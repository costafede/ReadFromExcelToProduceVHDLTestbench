-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            18, -8, -8, 4, 14, -9, -14, 20, -15, 16, 9, -2, -3, -12     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -4, -23, 70, 97, -125, -115, 123, -86, -83, -65, 28, 89, -22, 29, 65, -105, -18, -124, 98, 24, -37, 84, -37, -12, -125, 6, 16, 107, 117, -77, -22, -83, 30, 112, -96, -95, 52, 36, -53, -113, 31, -62, 67, 88, 78, 18, 25, 83, 50, 55, 24, 112, -75, -35, 72, 56, -120, -122, 2, -25, -3, -127, -114, -115, -123, 26, -11, 91, -7, 53, 94, 45, -118, -36, 17, 17, 81, -49, 26, -58, -3, -2, -69, -92, -40, -70, 67, -96, -6, -115, 116, -80, 111, 41, 42, -71, -114, -76, -124, -62, 27, 72, -98, -42, -33, -52, 42, -74, 36, -68, 112, 93, 110, -63, 110, -128, -121, 108, -32, -21, 95, 50, -21, -36, -16, -49, 93, 91, -9, -45, -48, 43, -88, 73, -105, -126, -62, 44, 41, -45, -6, 93, 40, 56, -42, 121, 109, -103, -103, 103, -48, 95, 83, -37, 31, -33, -20, 127, -112, 86, -122, -26, -71, 127, -4, -70, -115, 113, -69, 84, 23, 27, -1, 10, 103, 43, 91, 48, 46, 109, 94, -78, -102, 73, 15, -4, 84, 18, -13, -84, -126, 23, 4, -105, -101, -53, -46, 8, -91, 79, -90, -97, -49, 120, 8, 46, 120, 70, 8, 79, -101, -28, 14, -105, 31, 57, 45, 90, 68, -47, -20, 59, -55, 47, 18, -3, -123, 16, 42, 53, 116, -103, -18, 108, 107, -35, 47, -16, -68, 94, 112, -39, 85, -9, 74, 103, -19, -127, -20, 30, -3, -58, 117, 69, -92, 47, -25, 65, 49, 9, -39, -41, 78, 99, -62, 84, -86, 84, -34, 106, 40, -4, 30, -96, 87, 56, -4, -37, 8, -119, -113, 37, 53, -13, -88, 88, -58, -34, 113, -79, -100, -52, -82, -23, 97, 65, -30, 84, 7, -117, 60, 124, 122, 120, 105, 55, -105, -30, 72, -13, 41, -101, -96, 126, 104, -57, 108, -96, -97, -87, 22, 29, -21, 110, -32, -109, 1, -9, 31, -72, 21, 74, 74, 107, 26, -90, -50, -8, 118, -113, 98, 17, -60, 114, 60, 97, 100, -44, -17, -75, 122, -38, -6, 13, 77, 106, 8, -77, -94, -57, 2, 9, 16, -18, -63, -78, -3, 110, -4, -30, -75, 91, 54, -31, -57, 4, 117, -76, 86, -44, 80, 46, 79, -68, 68, 17, 64, -124, 85, -90, 60, 103, -117, -33, -17, 91, 85, -60, -19, -92, -68, 108, 13, -109, 97, -107, 72, 104, 51, -48, -4, -112, 36, 0, -77, -52, 118, -57, 90, -68, -44, -80, -114, -65, -61, -82, 95, 109, 85, 62, 65, 21, -18, -7, 60, -39, -54, -43, 74, 105, -36, -96, 39, -81, -63, 82, -85, -90, -43, 108, -31, 96, -80, 113, 96, 18, -76, -13, -90, -58, 20, 91, -6, -44, 82, -66, 114, 116, 118, 97, -108, 35, 45, -33, -58, 70, 6, -68, 7, -23, 121, 112, 11, -121, -125, 67, 26, -12, -59, 121, 91, 0, -38, 64, -94, -126, -39, -64, 104, 28, 109, 4, 68, -18, -99, 56, -26, 47, -45, 126, 119, 65, -25, 71, 32, -113, -32, 55, -103, 48, 14, 4, -66, -22, 103, 60, -46, 6, 52, 41, 82, -4, 88, 64, -53, 21, 111, 64, 118, -45, -70, 37, -112, -38, 102, 95, 82, -114, -42, 3, -38, 3, -123, -53, -58, 80, 39, -73, -30, 72, 65, -12, 32, 126, -3, 31, 76, -120, 85, -63, 104, 26, -18, -112, -38, 75, 84, -63, -125, -87, -78, 8, 94, 66, -27, 122, -84, 84, 25, -3, 36, -51, 26, 1, 53, 113, -2, 25, 121, -21, -88, -61, 51, 20, 63, 10, 97, -96, -23, 58, -30, -103, 2, 87, 85, -37, 125, 59, -12, 74, 76, 105, -80, 126, -124, -9, 66, 29, -5, -27, -60, 46, 2, 67, 27, 32, -33, -117, -101, 1, 82, 29, -78, -116, -54, 3, -124, -104, -89, 49, -98, 58, -38, -97, -67, 30, -67, -2, 45, 61, 82, -3, 67, -19, 74, -27, 94, 107, -15, -70, 71, -79, 48, 5, -128, 69, -22, 116, 88, -45, -80, -58, 123, 100, 28, -95, 46, -41, 3, 16, -124, -94, 35, 115, -122, 5, -127, -122, -13, -120, 97, -92, 93, -89, -120, 10, -102, -22, 85, -67, 61, -126, -70, -98, -49, 3, 72, 67, 111, -42, 72, -122, -124, 8, -107, -109, 99, 5, 53, 74, -85, 8, -94, -49, -120, 53, -16, 85, -96, -62, 88, 54, 72, -20, -127, 97, 28, 9, -16, 44, 32, -89, -24, -19, -61, 14, 61, 51, 52, -87, 62, -117, 2, 62, -105, 0, 64, -84, 55, 6, 120, 73, -6, -122, 124, -128, -7, -16, -9, -41, 1, -35, 84, 44, -126, -93, 77, 16, 29, 99, 16, -113, 52, 49, -62, 7, -14, 85, -15, 42, -79, -50, 87, 49, 96, 46, 89, -86, 87, -99, -126, 69, -1, 29, -7, 95, -2, 50, 82, -55, 24, 93, -77, -11, -21, -34, 98, -106, -53, 100, 121, 50, 33, 111, -110, -91, 101, 17, 64, 27, 25, -15, 41, -10, -47, -52, 83, -103, 84, 106, -61, 47, 111, 70, -31, -98, -50, -116, 29, 73, 43, -48, 92, 118, -42, -69, 86, 110, -88, -10, 7, -100, -95, 83, 71, -23, -78, -90, -72, 12, -14, -79, 121, 79, -90, 31, -18, -52, 61, -92, -106, 82, -84, -25, -44, -17, -21, -64, 108, 59, 65, -118, -97, 111, -59, 22, -18, -20, -13, -51, 113, -61, -24, -66, -94, -91, 33, -73, 5, -53, 5, 7, 20, -121, -81, 20, -128, -117, -99, 24, 112, -89, -100, -127, -89, 90, 14, -59, 74, -60, -77, -128, -88, -67, 68, 68, -44, -89, -20, 58, -40, -72, 127, -112, 35, -8, 15, 28, -119, -112, -102, 73, -96, -32, 79, 81, -61, -81, -52, 106, -104, -128, 11, 110, 88, 111, -22, 107, 121, 67, 5, -52, 32, -115, -2, -82, -118, 46, -123, 50, -88, 127, -42, 45, 68, -54, -104, -102, -5, 10, -62, 101, -79, 117, 67, 10, -5, -75, 76, 54, -55, -43, 113, -128, 33, 66, -102, -52, -30, 109, 82, -21, -55, -99, -37, -15, -110, -88, 77, -69, 87, -126, 51, 76, -104, 33, 91, -29, 78, -47, -42, 91, -109, -98, 72, -126, 37, -120, -110, 62, -61, 62, -1, -110, 78, -11, 82, 121, -27, 27, -21, 81, -78, 120, -37, 89, 22, -97, 92, 24, -110, 15, -41, -97, -9, -23, -78, 75, -128, 73, 81, -120, 104, 89, -40, 93, 116, -118, -11, -128, -38, 100, -126, -103, -10, -60, -42, -11, -28, -46, -104, -46, 74, 91, -92, 17, -111, -92, -71, 127, -109, 57, -35, -23, 67, 37, 126, -70, -84, 47, -95, -18, -53, -69, 105, 102, -73, -42, -91, 81, 97, -74, 17, -98, -53, 112, -90, 29, -126, -47, -28, 68, -73, 8, 43, -66, -116, -116, -110, -14, -114, 12, 9, 84, 7, -121, 62, -64, -23, 109, 25, 1, 99, 17, -35, -6, 12, -45, -82, -89, 55, -3, -32, 103, -72, -125, 55, -8, 94, 56, -122, -98, -118, -92, -112, -3, -47, 119, 34, 90, -123, -50, -5, 53, 97, 30, -66, -38, -44, 2, 88, 12, -97, -62, 4, 109, 53, 40, 127, 36, -2, -83, 115, -14, 42, 46, 106, 39, -120, -27, -74, 126, -82, -71, 124, -9, 98, -5, 85, 27, -69, -43, -57, 98, 89, 9, 87, 60, -79, 30, -48, 55, -66, -67, -77, 79, 70, 29, -22, 38, 23, -127, 23, 63, -28, 12, 51, -36, 23, -41, 123, 13, 116, -108, 109, 76, 15, -125, -94, 34, -12, -63, -48, -85, -77, 22, 27, 20, -90, 2, -108, 116, -106, -28, 66, 51, -55, -75, -101, -76, 73, -114, -56, -65, 38, 93, 58, -37, -103, -82, -72, 5, -18, -83, 127, 35, 6, 101, -36, -48, -44, 69, 90, -2, 52, 115, -2, 24, -112, -97, -74, 96, 116, -72, 82, 103, -32, 17, -64, 91, 120, 84, 66, -122, 8, -9, -96, -128, -109, 34, 69, -30, 50, -89, 43, -35, 45, -107, -120, 105, 87, -39, 75, 95, -122, -79, 43, -20, 112, -18, -124, 28, -100, -105, 88, 1, -26, 72, -17, -71, 45, 126, 40, 47, 97, -79, -8, -88, 12, 70, 20, 26, 88, -56, 118, -10, 68, -40, -63, -59, -49, -52, -75, -49, 64, -60, 77, 104, -49, -4, -118, 61, -120, 96, -51, -30, -7, 62, 30, 86, -66, 44, 70, 8, -51, 74, 9, 90, -107, -7, -115, 118, 27, -27, 79, 112, -38, 118, -73, 76, -28, -24, -63, -24, -70, 99, 102, -100, 114, 122, -90, -88, 127, -92, 17, 52, 62, 42, -7, 45, -41, -95, 118, -127, 94, -15, 73, 84, -118, -55, 78, 74, -76, -35, -17, -80, -4, -18, -22, 31, 41, 23, -48, -72, -110, 112, -32, -27, 36, 23, -25, 73, 117, -117, -55, 13, 0, 98, -40, 99, 120, -11, 36, 72, -17, -90, -86, -86, 99, -20, 36, -103, 65, 16, -28, -64, -85, 59, 6, -61, 84, 71, -107, 70, 57, 95, -126, 82, 68, 64, 50, 20, 124, 98, 63, -67, 75, -5, -23, -102, 18, -44, -60, 72, -78, 104, 107, -15, -82, 82, -126, -16, 93, 121, -63, -116, 4, -37, -83, 47, -44, 103, -67, -63, 3, -15, -59, 101, -91, -63, -79, -39, -3, -70, -116, 125, 107, 122, 99, 4, 107, -106, 0, 29, 25, -56, 21, 21, 77, -65, -90, 75, -123, -25, -59, 14, 5, 37, 24, -41, 19, 25, -89, -21, -41, 99, -60, -96, 66, 87, 1, 51, 9, -35, 1, -55, 55, 6, -15, 0, -81, 126, 109, -84, 115, 24, 62, 62, 1, -41, 106, 1, -85, 95, 64, -127, 31, 108, -70, 78, -36, -4, -51, -11, -39, -82, 51, -13, -125, -47, 124, 75, 4, 16, 21, 49, 72, 112, -101, 101, 33, -15, -96, -121, -109, -97, -123, -17, 102, 64, 19, 54, -22, -105, 37, 70, -62, 24, 30, 103, 32, -29, 59, 101, 12, 127, -54, -103, -123, -111, 91, 50, -100, -108, 34, 10, -44, -8, -61, -31, -80, -109, -59, -48, 84, -128, 70, -101, -61, -48, -86, 99, -23, -17, 20, 125, 113, 74, 18, -14, -100, -86, 72, 19, 99, 63, -33, -34, -6, 81, -31, 54, 105, -32, 97, 15, 102, 4, -95, -87, 2, 83, -9, 2, 35, 44, -128, 29, -42, 105, -61, -19, -17, -52, 95, -43, 27, 33, -16, 109, -87, -45, 42, 116, -37, 51, -36, -118, -70, 84, 40, -115, 87, 51, -27, -40, -92, 25, 77, -70, 67, 127, 10, -93, -83, 74, 46, -98, 53, 98, 54, 37, -101, 82, -49, 121, 101, -30, -14, 59, -105, -39, 63, 3, -87, -117, -14, 91, -37, 118, -51, 81, -110, 4, -102, -82, -102, 90, -4, -54, 86, -115, 74, -24, 116, -89, -104, 7, 12, 80, -22, 59, -33, 66, 10, 122, -29, 73, -124, -4, 33, -17, -17, -12, -69, -110, -19, 36, 20, 37, -103, -112, -25, 13, -30, 91, -78, 91, -7, -51, 15, -25, 31, -77, 84, -107, -119, -43, 17, -23, -25, -30, 118, -54, -82, -5, 59, 36, 91, 84, -31, 1, 98, -93, 74, 112, 86, -97, 84, -14, -127, -68, -19, -17, -20, 2, 5, -28, 127, 36, 79, 18, 110, -124, 51, 116, -10, 10, -99, -4, 6, -2, 46, 15, -76, -54, 37, -119, -28, 50, -59, -16, 121, 21, 11, -101, 89, -25, 56, -57, 48, 109, -117, -27, -121, -50, 16, -127, 100, 59, -78, 80, 96, 17, -88, 36, -92, 84, 17, 76, 47, 53, -1, 41, -38, 83, -29, 18, 80, 90, 48, -4, -64, -41, 48, -58, 15, -10, 21, 69, 41, -47, 66, 14, 16, 107, 57, 119, 93, 1, -23, 15, 115, -97, 22, -59, 65, -55, 13, -82, 56, -68, 99, 33, 82, -62, -90, 11, -97, -43, -73, 26, 53, -31, 72, -35, -1, 119, -85, 125, 16, 121, 116, -118, 52, -27, -108, 101, 7, -83, 40, -97, 58, 42, 53, 30, -104, 93, 63, 34, 17, 127, -49, 77, -126, -76, -27, -87, -38, 104, -51, -56, 19, 30, 115, -46, -57, -80, 3, 57, -33, 69, 89, -54, 66, -98, 76, -31, 102, -60, 79, 55, -72, 112, -82, 26, -30, 0, 103, 44, -16, -11, -77, 94, -120, 28, 3, -80, -77, -94, -68, -121, 117, -118, -31, -49, -9, 57, -127, 89, 70, 47, -89, -104, 85, -42, 28, 5, -28, 35, -76, 93, -7, -96, 25, -86, -37, 121, 78, -1, 19, -38, -40, -120, 77, 104, 124, 92, 22, -38, 118, -85, -16, 70, -43, -83, 112, 75, -8, 15, 19, -47, 46, 84, -114, -22, -34, -101, 19, -124, 76, 47, 102, -115, 65, -114, -110, -62, -82, -70, -112, -96, 100, 10, 88, 10, -108, -87, 96, 92, 0, -16, -28, -47, -122, 63, -67, 35, 77, 56, -44, 19, -61, -15, 78, -14, -103, 48, 37, -7, 105, -64, 27, 54, 47, 116, 109, -88, -10, 77, -125, -77, -19, -122, -14, 94, -60, -20, 120, 69, -64, -86, 23, -98, 108, -121, 100, 103, 46, 64, 18, 90, -30, -95, 51, 101, 98, 62, 54, -6, -14, 10, -31, -66, 65, 82, -79, -83, -68, -49, -119, 48, -17, -56, -19, 7, -123, -35, -35, 65, -39, 24, 21, 61, 125, -11, -3, 42, -127, -114, -44, 86, 37, 1, -119, 56, -53, 54, -24, 25, 17, -5, -127, 2, 79, -67, -103, 84, 26, -85, 74, 64, 110, -23, 51, 9, -12, -100, -70, -1, 94, -43, 74, 6, -128, 12, 14, 113, -19, -61, -116, 121, -53, 73, 74, -108, 99, 99, 36, 16, -2, -48, 80, -37, 124, 3, 33, -24, 35, 31, 62, -94, 5, -34, 86, -74, 1, -87, -116, 63, 68, 86, -126, 78, 115, 80, 68, 1, 58, 40, -73, -62, -96, 6, -27, -91, 124, -39, -126, -110, -23, -108, 50, -83, -91, 27, -75, 69, 13, -105, -49, 109, -79, 119, 117, -66, -65, -77, -68, 17, -82, 8, 118, 38, -12, -47, -120, 91, 47, 114, 111, 125, -21, 89, -24, 21, 80, 81, -102, -123, -78, 37, 82, -39, 79, -127, 105, -110, 30, 119, -10, 91, -45, 8, 104, -46, -107, -2, -82, -24, 119, -53, 94, 38, -2, -40, -23, 40, -107, 39, -113, 85, -99, 121, 16, 72, -69, 10, -36, -117, 0, -23, 69, 36, -51, -45, 61, -23, 43, -62, -1, -19, -7, 126, 29, 109, -45, 89, 60, -121, -1, 14, 95, -63, -67, -25, 41, 23, -40, -33, -22, -51, -16, -66, 64, 92, -106, -72, -50, -47, -107, -113, -97, -59, -38, -105, 47, 23, -14, 104, 31, -76, -8, 115, 5, -114, -14, -64, -13, -57, -101, -63, -116, -29, -17, -2, 112, -46, -15, 44, -19, -64, 77, -19, -32, -127, 102, 13, -105, -122, -92, 21, 107, 72, 21, 125, 10, -93, 82, 104, 13, -33, -25, 68, -121, 124, -21, -79, -116, 3, -15, 87, -87, -11, -6, 90, 80, -23, 119, -23, 70, -101, -31, -35, -103, -113, -7, -50, 13, -111, -89, 65, 83, 99, 56, -86, 39, -46, -20, 105, 113, 102, -9, 73, 88, 54, 62, 29, 63, -27, -9, -128, 90, -120, 97, 3, 57, 47, -9, 58, -79, 26, -20, 47, -99, -55, -55, -94, -123, 9, -11, -101, -100, 100, 120, -116, -59, -128, 50, 115, 114, -100, 37, 83, 6, 87, -8, -122, 70, 103, -120, -54, 24, -40, 80, -89, -65, -44, 54, 108, 29, 85, -45, 25, -4, 59, -56, -40, -59, 22, -102, -121, -21, -76, -115, -109, -11, -55, 11, -28, 40, 120, 2, 16, -5, 38, 63, -124, -114, -102, -99, 16, -3, 31, 77, 110, -31, -109, 97, -35, 48, -123, 62, 52, -35, -48, 33, -67, -113, -115, -50, -86, 111, 21, -4, -32, -53, -103, 68, 37, 11, 31, -57, -119, -77, 103, -111, 13, -106, -31, 32, -18, 49, -6, -125, -7, 60, 115, -27, 28, 42, 101, -18, -83, -70, -57, -68, 77, -25, -68, -112, 88, -86, -54, 127, -77, 72, -76, 89, -94, -111, -33, 35, 87, -30, -96, -44, 48, -35, -86, -115, -80, 14, 55, 12, -81, 80, 98, -91, -80, -47, -21, -118, -50, -117, -90, 107, -80, -24, -39, 11, -30, 109, 92, 95, 15, 112, -106, -40, 111, -40, -69, 104, 46, -60, -28, 105, 16, -110, 20, 11, -7, -30, -113, -120, 83, -102, -34, 67, -44, -91, 107, 92, -98, 46, 23, -22, 30, 36, -4, 82, -107, 78, -128, -98, -90, 70, 41, -28, -128, 104, 106, 40, 69, 46, 49, -122, 115, -94, 11, -86, -91, -13, 31, -116, 38, 47, -122, 11, -21, 74, -14, -89, -104, 108, 49, -79, -28, -58, -119, -38, 117, 53, -12, 25, 29, -122, -72, -69, -62, -69, -38, -125, 97, 54, -37, 36, 43, -53, -106, -102, -101, -51, -111, 26, -19, -31, 87, -126, -128, 18, 101, -2, -122, 118, 1, -25, 47, -108, -53, 118, 42, -8, 62, -34, -12, 40, 105, -93, 53, -117, 10, 47, -128, 120, 66, 36, 72, -112, 19, 94, 74, 121, -80, 38, 126, 120, -48, -126, -97, -32, 125, -124, 73, 121, 79, -109, -90, -111, 10, 78, -49, 24, -61, 12, -6, 82, -121, 127, -39, -80, -46, -127, 97, -12, -8, 51, -2, 36, -113, -115, 58, -104, -52, 2, -53, -67, 24, -18, -122, -105, -109, 111, 64, -45, 18, -72, -74, -68, -96, -1, 95, 43, 24, -68, -40, 24, 110, -32, -124, -49, -86, -8, 97, -124, -86, -45, -31, -125, -78, -95, -59, 61, -99, -86, -101, 89, 46, -50, 96, 45, 36, 62, 66, -101, -21, 3, 3, 92, 20, -64, -92, -32, -118, -55, -115, -56, 95, 49, -121, -58, 24, 16, 126, 122, -85, -46, -124, 21, 25, -56, 15, -126, 43, 113, 51, 69, 15, 75, -90, 24, -78, 121, 94, 97, 63, 98, 119, 42, 93, -61, -106, -80, 88, 83, 123, -57, -111, 53, -67, -87, -122, -117, 97, 118, 114, -2, -24, -114, 46, 126, -26, 8, -57, -112, -9, -114, -95, -48, 94, 38, 15, -2, 57, 66, -3, -16, -69, 42, -101, 82, -119, 71, -28, 34, -91, -109, 4, -111, -38, -64, -123, -108, 27, 71, -22, -57, -118, -11, -73, 127, -9, -87, -85, -54, 22, -20, 82, -94, -121, 5, -97, -46, 127, -59, -52, -4, -33, 85, -3, -106, -64, -105, -90, 0, -105, -58, -110, 124, -114, 102, 92, 59, -18, -121, -113, 12, 96, -47, -9, 28, -69, 88, 120, -109, 28, 83, 89, 31, -96, 116, -7, -107, 108, -37, -22, 74, -82, 9, 124, 52, -1, -26, -99, -118, 22, 108, 66, -61, -99, 47, -61, 104, -24, 53, -11, -63, -41, 90, 76, 22, -107, -12, -59, -61, -92, 117, 125, 48, 95, 9, -95, 123, -101, -28, -109, -31, 116, 11, -47, -108, -7, 50, -79, -69, -6, 57, 127, -11, 2, 62, 0, 73, 52, -86, 4, 108, -109, 25, -93, -5, 63, 49, -89, -47, -72, -127, -46, 56, -62, 76, 25, 92, -28, -118, -83, -27, 35, 20, 107, -47, -57, 94, -111, -100, 74, -68, 105, 33, 7, 17, -83, 75, -20, -77, 50, -6, -28, 77, 51, 97, -70, -119, 102, 73, 90, -46, 63, -114, -2, -17, -61, -29, -79, 81, 15, 10, -7, -59, -110, 0, -60, 49, -119, 74, -33, -94, 21, 106, 95, 118, -108, -101, 96, 75, -104, -52, -106, 108, -51, -118, 33, 2, 56, -27, -62, -67, -46, 87, 118, 115, 109, -74, -123, -100, 111, -109, -36, -98, -66, 54, -88, -108, 82, 120, 29, 46, -17, -32, -54, -94, -13, 43, -3, 38, 47, -74, -67, 96, 94, 22, -10, 124, 31, -99, -84, 35, -126, -14, -14, 97, 81, 109, 22, 12, -128, 126, -90, -7, -80, 79, 22, -112, -110, 19, 125, 29, 55, -75, -108, -88, -69, -12, -115, -59, -97, 126, 46, -17, 101, 109, -125, 123, -44, -116, -38, 41, -93, 4, 115, -64, 127, -60, 95, -125, 59, -53, 41, -115, 3, -15, 94, -53, -61, -91, 66, -13, 97, -79, -30, 62, 115, 72, -7, -50, -36, -93, 13, 47, 47, -109, -97, 11, -88, 73, -62, 0, -51, 16, -65, 121, -100, -106, -22, -115, -14, -18, 39, 110, -96, -15, -87, -105, 70, 100, 121, 3, 111, -105, 96, 51, -81, 27, -65, -105, 121, 57, 127, 51, -74, 14, 28, 74, -123, -67, -69, -126, -56, 30, -69, -45, -73, -33, 123, 89, -51, -47, 22, -62, 6, 94, -58, 51, -43, -72, -73, -108, 77, 54, -112, 76, 22, 125, 15, 94, -112, 45, 16, -100, 49, 101, -7, -15, 94, 124, -37, 79, -87, -72, -66, -10, -52, -92, -90, -20, 9, -124, 100, 100, -105, -13, 2, -49, 62, -100, 56, 127, -88, -92, 29, -86, 92, 10, 113, 127, -65, -95, 124, 103, -87, 62, 107, 50, -114, 3, -37, 80, -53, 30, -81, 123, 11, 78, 12, -101, -13, 90, 29, 56, -29, 94, 19, 61, 124, 4, 89, 42, 61, -51, 95, 37, -81, -22, 27, -68, -81, -125, 16, 37, 31, -49, 42, 110, -65, 54, 111, -62, -93, 2, 59, 11, -20, 78, 65, 126, -123, -15, -103, -65, -57, 71, 76, -48, -77, 126, 98, 2, -115, 1, 53, 84, 90, 121, -23, 74, 115, -78, -67, 21, 10, 115, 89, -20, -12, 51, 29, -6, 73, -1, -71, 88, -64, -125, 4, -92, -6, 55, 121, 115, 119, 102, 126, 30, 101, -113, -76, -85, 63, -96, -51, 110, -61, -108, -51, 97, -36, 88, 12, -103, 100, 9, -126, -67, 62, 42, 117, 47, -74, -110, 62, 98, -28, -111, -28, -102, -81, 84, -14, -87, 4, 47, -47, -71, -27, -115, -40, 68, 63, -114, 123, 33, 6, 83, -118, 81, -122, -105, 96, 60, 119, 19, 66, 90, 121, 102, 118, -65, -104, 80, 35, -68, -81, -31, -24, -81, 42, 83, -85, -115, -20, -60, 78, 80, 57, -67, -124, -107, 39, 27, -29, -85, 59, 65, 42, -23, -103, -4, 93, -128, 10, -4, -91, -77, -14, -109, -71, -49, -8, -107, 82, 95, 109, 4, -56, 74, 28, -93, -46, 12, -49, -39, -91, 48, -62, 77, -79, 46, 46, 101, -5, 84, -5, -108, -34, -98, -82, 19, 74, -102, 24, -77, -20, -47, 9, 96, -112, 113, -104, 121, 15, 26, 16, -113, -43, 106, -37, -103, -105, -33, -10, -124, 97, -108, -51, -81, 46, 37, -82, 13, 120, 99, 45, 86, 74, 36, 87, 103, 7, 40, 35, -8, -117, -25, 47, -116, -37, 60, -98, 93, -15, 63, 106, 83, -42, 50, -117, -117, 98, 70, -90, 62, -118, -17, 0, 106, 91, -6, -13, 24, 73, -41, -118, 29, 82, -43, 78, -10, 113, -116, 121, 88, -96, 23, 119, 7, -111, 21, 100, 121, 64, 107, -117, 17, -87, 5, -22, 102, 80, -121, -77, 39, -56, 43, -46, -124, 90, -2, -4, -73, 32, 23, -34, 11, -2, 71, -66, -1, -79, 11, 60, 77, -94, 122, 113, -44, 17, -95, -106, 2, -111, -12, 127, -18, -80, 18, -6, -109, -33, 20, 54, -22, 36, -3, 11, 74, 84, 81, 66, 81, -124, 61, -125, 97, 102, -97, -63, 11, 98, 127, -87, -14, -46, -43, 67, 78, -56, 38, -26, 9, -115, -1, -70, 89, 103, 74, -20, -67, -17, 5, -6, 87, 80, -24, 52, -51, -3, 36, 111, 76, -40, -47, -103, 43, -34, -117, -74, 46, -97, -22, 70, 81, 44, -77, 81, 94, -63, 43, 65, -63, -17, 92, -128, -25, -8, -21, 25, -74, 105, -102, -81, 22, -119, 107, -56, -5, -49, 79, -74, -99, 68, -119, -48, 81, -112, 119, 62, -124, 93, -19, 69, -26, -24, -128, 91, -57, 92, -63, 74, -116, -116, 15, 47, -77, 72, 48, 118, -68, -122, 68, -63, 57, 18, 74, 11, 58, -80, -47, -51, -50, -79, 46, 6, -24, 99, -56, -1, 102, 22, -107, 14, -80, -114, 18, -81, -4, 27, -46, -18, 31, -100, 60, -2, -85, 101, -97, 84, -74, -112, 42, 113, -25, -47, -22, 60, 26, -73, -29, 84, 61, 41, -80, 84, 22, 64, -32, -6, 74, -91, 121, -101, -91, -102, 64, -28, -43, 120, 20, -61, -20, -82, -19, 115, -122, 20, 90, 88, 125, 95, -90, -67, -29, -37, 80, 34, -28, -36, 113, -37, -57, 58, -75, -27, 38, -79, 52, 104, -4, -94, -22, 41, -8, -59, -22, -107, 0, 54, -42, -32, 59, 10, -6, -121, 15, -63, 81, 18, -19, -118, 121, -44, -93, -27, -124, 112, 69, 2, -27, -38, -15, -48, 56, -120, -53, 37, -59, 90, -38, 34, -19, 86, 75, -112, -43, -39, -125, 37, -86, -105, 53, 72, 118, 69, 14, -53, -115, 38, -79, -24, -85, -16, 99, 75, 36, -92, 40, -115, -114, 64, -55, 88, 9, 93, 101, -95, -98, -54, 122, 9, 95, 112, -80, 111, -128, -102, 62, 78, -2, -57, 85, -121, -7, -97, -58, 29, -5, -93, 122, -57, 16, -44, -87, 40, 103, -76, 9, 51, 95, 98, 98, 48, 83, 11, -124, 42, -52, -16, -77, 52, 20, -25, 10, -16, -6, -36, -74, -100, -91, -89, 22, -95, 70, 49, -79, 89, 111, -61, -23, -45, -73, 21, -70, -40, 28, 31, 118, 57, 96, 121, 15, -38, -56, -91, 73, 57, 4, 36, 78, -115, 46, 74, 44, -21, -19, 105, 50, -31, -107, -78, -106, 67, -32, 79, 15, 36, -114, -64, -109, 118, 107, 101, 126, 103, 86, -36, -71, -4, 105, -18, 95, 22, -6, -38, 122, 53, 5, -106, 120, -89, -97, -48, 89, 64, 123, -77, 102, -42, -113, 113, -77, 42, 125, -9, -30, -2, 3, 44, -14, 77, 30, -114, 103, -27, 80, 6, -72, -101, 117, 81, 22, -115, 76, 126, 102, -89, 2, -28, -77, 90, -107, -54, -44, 24, 0, 33, 110, 59, 89, 50, 25, 36, -127, 123, -117, 38, 83, 17, -110, -57, 57, 23, 20, -64, 56, -62, 40, -123, -83, -124, 6, -16, 46, -24, 15, -44, -70, 63, -5, 31, -40, -19, 109, -36, -90, -64, -44, -70, 107, -71, 105, -93, 119, -25, 122, -127, -37, 81, 17, 47, -81, 5, 114, 73, -50, -45, 10, 70, -114, -128, -83, -46, -46, -67, -55, 101, 46, 62, 127, 86, 11, -112, 49, 101, -125, 11, 99, 99, 19, -123, -9, 36, -78, 42, 15, 103, -111, -41, 42, 18, 125, 91, -128, 104, 31, -8, -56, -50, -40, 44, -21, 86, -27, 86, -99, 90, -93, 117, -60, -59, 25, 77, -6, 4, 45, 38, 105, 29, 15, 86, 57, -82, -94, 105, -51, 38, -27, 43, -13, 125, 55, 7, -97, -104, -32, 114, 23, 78, 88, 26, 21, -7, 81, -14, 93, -39, -93, 93, 112, 98, -85, 5, 40, 119, -32, -119, -82, -39, -118, -120, -100, -112, -89, 70, -97, 56, -28, -123, -9, -26, -39, 37, -114, 95, 116, -28, 111, -95, 28, -70, 93, -82, 101, -26, -76, 108, 125, -56, 67, -76, -23, -6, -43, 6, -19, -65, 109, -39, -56, -111, 33, 102, 15, -95, -73, -11, -105, 109, -66, 41, -90, 72, 88, -100, -42, -32, 89, -100, -59, -63, -77, 83, 67, 7, 115, 14, 30, 15, 36, 40, 80, -68, -4, 19, 56, -70, 79, 108, 64, 33, 123, -59, -58, -23, -94, 44, 127, 119, 117, -15, -6, 97, 93, 108, 101, 119, 81, -34, -21, -94, -22, 43, -123, -55, -67, -44, 41, 80, 57, 14, -109, -37, -96, 27, -67, -58, 123, 84, -92, 67, -66, -116, 68, -60, -32, 15, -30, -57, -20, -105, 39, -107, -73, -66, -16, -64, -120, 51, 10, 52, 28, 1, -101, 103, -88, -60, -98, -124, -73, 68, -15, 61, -124, -92, 108, 91, 26, -68, 84, 118, -90, -72, 34, 89, -21, 109, 78, 107, 112, 63, 28, 52, 108, 71, 10, -94, -68, -103, 116, -114, 82, 110, 36, 34, -27, 109, -121, -72, 94, -93, 110, 54, 82, -120, -77, 52, -83, -112, 36, -119, 51, 57, 123, 42, 36, -97, 124, 15, 54, -2, 93, 11, -111, 108, -71, 120, 64, 103, -95, -13, -42, 34, 89, -62, -20, 75, -107, -95, -68, 102, -37, 96, -70, -106, 28, -87, 18, 94, -39, -29, 32, -128, 23, 37, 27, -20, 16, 55, -126, -125, -48, -119, -118, -6, 114, 51, 61, 25, -121, -3, -55, 7, 100, -94, -12, 89, -14, -122, 28, 64, 105, 80, 23, -55, -102, 93, -2, 83, 17, -88, -48, -63, 3, -102, -127, -104, -68, -111, -18, -103, -30, 34, -73, -36, -97, -119, 7, 97, -52, -71, -36, 60, 55, 52, -83, -58, -62, -33, 127, -103, 11, 2, -15, 49, 29, 45, 70, 77, -121, 33, 67, 1, 115, -87, 19, 92, 41, -70, 109, -49, 80, 9, 38, 103, -92, 119, 85, -85, 74, 86, 10, 26, -35, -22, 118, 66, 19, -14, -37, 124, 24, -82, -30, 31, -15, 92, 123, 14, -117, -106, -65, -101, -78, -46, -37, -28, 38, 23, -128, 70, -87, -87, -24, 100, -41, 110, 17, 111, 100, 28, -4, -113, 49, 25, 27, 33, 10, -68, -91, 36, 61, -23, -9, 68, 110, -70, -103, 27, 105, 44, 2, -119, -127, -70, 124, 6, 0, 18, -27, 50, -99, -79, 19, 71, 73, 103, 37, -105, 8, 37, 116, -57, 16, -14, 65, 25, -37, 96, -81, 72, -61, -87, 69, 123, -110, 16, 125, -60, -66, 112, -115, -118, -71, -71, -13, -75, 33, 110, 42, -105, -73, 10, 49, 115, -11, -46, 88, -63, -18, 82, -42, 85, -25, -55, -32, 77, -106, 93, 57, -54, 71, 84, -19, 123, -37, -51, -126, 121, -125, -64, 98, -32, 44, -63, -122, -17, -15, 87, -89, 41, 94, 64, 46, 99, -75, 17, -85, -29, -36, -65, -92, 11, -20, -21, 52, 64, -96, -70, -22, -40, 101, -86, -57, 125, 61, -21, -123, -122, 22, -18, -69, -44, 43, -19, 42, -123, 14, 23, -66, -37, 24, -119, 4, -36, -53, 117, 103, -33, 18, -68, -57, 112, 9, 87, -40, 87, -2, -46, -42, 73, -73, 124, 92, -88, -116, 67, -58, 80, 103, -102, 75, -91, -49, -88, 11, -80, 83, 108, -86, 38, -43, -66, 34, -6, -102, -11, 75, 31, -103, -59, 126, 75, -51, -60, 74, -22, 26, 65, 5, 73, -58, 96, 102, -63, 119, -70, 84, 112, -112, 95, -45, -44, -64, -34, 41, 21, 97, 118, 72, -107, -23, -24, -8, -126, 21, 56, 48, 102, -125, -95, 111, -81, -2, -4, -37, 32, -68, 88, 52, 109, 93, -109, 69, 7, 95, 111, -48, 123, -71, 28, 29, -11, -118, 30, 56, -52, -83, -57, -16, -2, 105, -47, -49, 57, -119, 63, -104, -12, 47, -95, -80, -93, 35, -36, -120, -89, 18, -37, 57, 44, -3, -70, 39, -57, -69, -90, -70, -63, -108, -84, 33, 30, 37, -34, 55, -35, -95, 84, 13, 82, 71, 120, -34, -24, -66, 21, 44, -40, -103, 70, 124, -27, -92, -61, -48, -9, -63, 5, 31, -105, -126, -24, 80, 6, 74, 86, 120, -59, 18, -95, 96, 116, 92, -15, 24, -20, -22, -127, -103, 53, 115, -20, -34, -90, -39, -68, 44, 123, 60, -79, -87, 50, -66, -55, -10, 118, -75, 75, -48, 77, 3, 125, -65, -87, 76, 102, -25, 71, -115, -62, -39, -99, -2, 103, -42, 118, -27, -87, -4, -15, -118, 19, 68, 46, -30, -124, -106, 117, -31, 124, 79, -54, 79, 46, -60, -43, -29, -86, 16, -49, -119, -25, 84, -63, 31, 126, -119, -27, -10, -9, 124, 124, -48, -32, 116, 50, -43, 15, -110, -95, 77, -43, -44, -35, 52, 38, 11, -2, -18, 93, 11, -83, 0, -12, 26, 114, -68, -4, 27, -90, -11, 12, -34, -91, 32, 72, -110, 22, 43, 72, 55, 36, 127, 106, -67, 94, 94, -77, 91, -15, 73, 69, -65, -10, 89, 41, 67, 79, -86, -11, 61, 2, -23, 70, -4, 61, -13, -122, -16, 15, 45, 112, 44, -4, 122, 0, -9, 40, 126, 93, -44, 50, 2, -125, -114, -98, 30, -30, -86, 9, 67, 38, -52, -14, -103, 73, -10, -80, -84, -106, -57, 102, 76, 81, 59, 2, -53, -9, 116, 42, -8, 97, -5, -39, -6, 77, 118, -64, 4, 78, -81, -15, 6, -39, 103, -3, 5, 100, -31, 47, 17, 22, -62, 95, -65, -51, -105, -123, -81, -100, -55, 102, 93, -103, 119, -8, -117, -124, 111, -127, -34, -8, 55, -44, 110, -55, 81, 2, -69, -91, -3, -17, 56, 55, -65, -107, -60, -104, -2, -81, -67, 89, 97, 30, -121, -61, -127, 73, 61, -46, 16, 73, -113, -9, -116, -116, -77, -107, -122, 59, 73, 56, -83, 25, -21, -2, 73, -101, 40, -64, 112, -6, 35, 20, -22, 32, 29, 110, -107, -40, -25, 6, -123, -23, -8, 6, -71, 68, 74, 104, 113, 119, 15, -95, -125, -104, -26, -53, -122, 122, -45, 27, -3, 20, 18, -104, 34, -31, -50, -101, -33, 127, 84, -83, 101, -62, 97, 76, 54, 92, -27, 100, -4, 4, 122, -9, 94, 9, -105, -44, 61, 25, 61, 87, 9, -28, -32, -9, -14, -29, 73, 52, -90, -39, -52, 124, 97, -52, 2, -128, 111, 86, 107, 76, 18, 114, -109, 73, 22, 125, -59, 56, -50, 118, -32, -86, -97, -21, -117, 49, 7, -42, -98, 95, -20, 27, -67, -4, -72, -41, -104, -12, -59, 24, 110, -94, -54, -5, 83, -69, -85, -66, 86, 31, -59, 123, -93, 108, 57, 79, -44, 82, -8, 29, -25, -42, -76, -40, 10, -91, 83, 42, 11, 57, 100, 41, 111, -128, -91, 14, -8, 16, -35, -112, 36, 127, -35, 75, 55, 88, -11, 22, -78, -9, 43, -7, -47, -124, 26, 56, -6, -100, 58, 110, -91, 1, -99, -48, 111, -113, 121, -120, 35, 117, 115, 116, -18, -127, -43, -47, 11, -15, 30, -26, -108, -31, -101, -51, 74, 119, -12, -107, 52, -40, -121, 48, 97, -31, 16, 5, -85, -1, 33, 28, 117, -57, -57, 47, 51, -12, -121, -77, 10, -38, 18, -67, 86, 74, -8, -51, -67, 67, 74, 104, -104, -21, 59, -96, -15, 8, -54, -25, -127, -55, 101, 50, 15, 57, -116, 122, 83, -38, 11, -37, -29, -52, -100, 37, 118, 38, 100, -50, 18, -48, -92, -115, 9, 29, -19, -46, 37, 83, 46, 44, 38, 62, -102, 5, 121, 23, 68, -100, -28, -116, 101, -19, 72, 11, -77, 120, -41, -21, 110, 30, -56, 46, 96, -102, -71, -73, -88, 125, 37, 12, -7, 77, -35, 65, -128, -50, 17, 5, -62, -63, 19, -44, 10, -56, 83, 17, 86, -103, -93, 29, -127, -22, -13, -5, 72, 46, -102, 125, 75, -97, -77, -46, -127, -86, 17, 60, 52, -3, -76, 70, 11, -51, 23, -12, 116, 107, -91, -101, -60, -98, -87, -90, -78, -35, 85, 31, 67, -48, -28, -115, 37, -41, 60, 103, -96, 79, -119, 88, 107, 83, 9, 60, 21, -60, 121, -27, 39, 33, 57, 50, 87, -89, 23, 106, 82, 41, -89, 43, -36, -71, -120, -28, 14, 81, -33, -55, -50, 9, -38, -23, -117, 17, -76, 65, -10, 68, -25, 7, 86, -91, 115, 89, -68, -53, -55, -55, -32, 44, 94, 60, -102, -86, 97, -97, 42, -127, 80, 103, 11, -88, 50, -5, 81, -118, -86, 124, 67, 79, 22, 90, 82, -69, 15, -7, -79, 21, -15, -46, 24, -53, -121, -126, 92, 123, 72, 75, -82, 49, -51, 69, 68, -33, 118, 17, -70, -55, 70, 106, 15, -58, -116, 98, 100, -75, -37, -8, 21, -103, -84, 121, -48, -15, -46, -41, -16, -26, 80, -57, -25, -19, -56, 4, -18, 30, 90, 80, 8, -125, -52, -49, -15, -72, -57, 112, 88, -121, 124, 119, 12, -66, 99, -89, -48, -15, -110, 32, -70, -79, -57, -101, -119, -77, 17, -82, -63, -46, -110, -128, 59, 78, 59, -91, -98, -85, -63, 47, 26, -110, -34, -17, 118, -100, -88, -10, -77, 60, 72, -38, 109, -80, -89, 74, -35, -3, 84, 86, 73, -12, -18, -121, 48, 91, 15, 56, -66, -75, -47, 94, 66, -39, -55, -42, 0, 0, 5, 63, 9, 97, -5, -9, -48, 58, -114, -82, -83, 83, 18, 32, -83, 18, 19, -121, -126, -71, -3, 61, -99, 35, -109, -72, 123, -14, 118, -12, 53, 58, 51, -103, -68, -81, -21, -54, 60, 51, 78, -27, 62, 43, -32, -83, 21, -11, -67, -82, -86, 57, -13, -18, -94, -60, -26, 114, 59, 72, 6, -61, 33, 16, -116, -18, -69, -109, -19, -17, -116, 38, 110, -103, 70, -88, 71, 34, -24, 28, -33, 20, 58, 5, -9, -4, -15, -114, 96, 104, -67, 81, -97, -103, 89, 43, 42, 41, -88, -127, -92, 104, -5, 52, -24, -58, -75, 4, 100, -126, -25, 94, 91, 16, -99, 89, -109, 84, -82, -98, 51, 57, -43, -81, 15, 91, -12, 66, -77, 20, -113, 33, 3, -59, -84, -54, 108, 71, -113, -34, -30, -41, 96, -98, 35, 95, 114, 29, 91, -113, 48, 127, 72, 43, -1, 12, -118, -11, -58, 70, -78, -97, 122, -93, 21, -97, 98, 91, 16, -20, -10, 78, -32, -107, -99, -27, -62, 32, 115, 24, -92, 126, -52, -116, 57, -119, -33, -1, -44, -5, -40, -116, 33, -83, 71, -115, 43, 113, 36, -104, 12, -9, -19, 106, -112, 63, -41, -26, -74, -54, 83, -82, -50, -107, -118, 29, 123, 51, 95, -124, 42, 44, 46, -97, 94, -117, 87, 42, -5, -123, -8, -1, -85, 94, 118, -62, -16, -73, 8, 63, -20, -10, -96, -122, 95, -70, -22, -100, -44, 80, 84, -83, 61, 117, -83, -23, 119, -111, -42, 50, -118, -30, -22, 126, -109, 27, 3, 119, -120, 70, -6, -96, 10, 9, -54, 67, -27, 41, -105, -42, 82, 29, -111, 54, -44, -87, 20, -3, -112, -81, 127, -115, 96, 88, -1, 119, -26, -44, 71, -125, 126, -49, -31, -99, -34, 124, -99, -12, -115, -114, 70, -45, -27, 38, -64, 46, -108, -102, -122, -58, -59, 112, -47, -86, 87, 68, -51, 70, -122, -117, -47, -69, 30, 88, 96, -103, -126, -62, 2, -125, -118, -35, -45, 10, -3, 1, -8, -7, 7, -8, 2, 67, -114, 50, 15, 2, -100, -38, -121, -46, 43, -58, 63, 50, 111, -50, 11, -14, -105, -52, -89, 41, -87, -70, -93, -53, 11, 6, -95, -28, -92, -32, -51, 59, -117, 86, -3, -72, 49, -55, -80, 71, 82, -123, 78, -66, -123, 6, 48, -84, 113, -77, -84, 37, -126, 122, -5, 118, 78, 89, 25, -66, -55, -81, 95, 25, -110, -115, -22, 20, -77, -28, 24, 22, -27, 114, 101, 4, 99, 63, 68, -23, -102, 88, 97, 98, 88, 76, -114, -9, 98, 48, 14, -88, -51, 34, -98, -67, -112, -3, -12, 25, -112, 118, 96, -66, -44, -93, 45, 90, 40, -37, 18, 59, -39, 92, -50, 110, 3, 83, -47, 26, -52, 103, -101, -95, -95, -91, -43, -56, 60, 29, -7, -55, -126, -10, -68, 38, 99, 125, -1, 122, -27, 58, 8, -68, 75, -49, 98, 107, -126, 94, -46, 119, 109, -62, 89, -7, -67, 22, 100, 68, 18, -93, -110, 59, -12, 11, -5, 102, -52, 77, -8, -15, 80, 61, 96, 52, -44, 55, -110, 120, -36, -82, 51, 115, 26, 95, -54, 125, 94, 5, 28, -121, 4, -79, 83, 76, -80, -47, 20, -72, 25, 80, 44, -50, 95, 35, 40, -107, -38, -24, 56, 124, 80, 27, -82, 46, -64, -43, -71, 19, -13, 5, 61, -28, 24, 109, 10, 116, 98, -1, -65, -95, 87, 115, -32, 68, -47, -85, 89, -55, -100, 54, 65, 41, 27, -11, 42, -7, 47, -86, -1, -107, 47, 1, -98, 25, -64, -111, -121, -105, 3, 108, 5, 123, -35, 1, 125, 99, -13, -39, 11, 7, -67, -22, -123, 44, 27, 38, -19, 71, 90, -10, 124, 84, -40, 12, 35, 112, -41, 5, 89, 29, -22, 78, 19, 85, -125, -13, 53, 121, 115, 104, 126, 73, -22, -126, 109, 71, -47, 69, 118, -45, -48, 94, -48, 51, -75, -24, 64, 61, 14, -77, 5, -48, -31, 109, -22, -87, 122, 122, -33, 24, 0, 58, -87, 4, 8, -127, 111, 10, 27, -60, -82, 51, 22, -54, -46, -81, 1, 113, 88, 56, -115, -74, 1, -112, 26, 70, -34, 61, 46, -17, -21, -110, -82, -84, -125, -115, -39, 127, -27, 109, -57, 79, -47, 100, 79, -22, 98, 44, 69, 118, -96, -50, -11, 1, 30, 117, 23, 45, 110, 58, -90, 116, 104, 75, 8, -68, 102, -32, 125, 99, -43, 13, -6, 110, -62, -66, -10, -41, 20, -68, -73, 93, -57, 90, -79, 65, -61, -64, 110, 68, 97, 127, -9, -101, -21, -91, -2, -46, 77, 42, -64, 62, 5, -115, 60, -15, 93, 55, 117, 1, -110, 75, -77, -1, -36, -125, -92, -10, -12, -46, 121, 104, -22, 29, -3, -23, -39, 101, -86, -21, -39, 24, -111, 72, -102, 81, -89, -49, 74, -41, 35, -92, -53, 90, 7, -45, -41, -1, -9, 15, 30, 59, 31, -108, -102, -10, -52, 127, -37, 98, -23, 14, 96, 38, 28, -23, 37, -18, -86, -98, 94, -121, -119, -43, 96, 96, 59, 106, 122, 23, -120, -93, 30, 85, 54, -115, 67, 106, 10, 26, 2, 116, 123, 116, 50, 80, 65, -21, 95, -64, 63, 11, -122, -30, 79, -47, 97, 100, 113, 21, -86, 4, 27, 8, 48, 101, -62, -115, -7, 119, 34, -120, -23, 53, -2, -97, 24, -29, 76, 4, -93, -91, -46, -25, -112, 34, 33, 7, 48, 47, 124, 105, 60, -16, 71, 40, -99, 91, -117, -24, 119, -11, 104, 18, 63, -38, 89, -53, 115, 77, -25, 60, -87, 11, 107, -9, -27, -42, -36, -27, -79, 17, 99, -73, 7, 93, 1, 26, -21, -114, -60, 17, -86, 7, -27, -56, -48, -47, 98, 31, 92, -110, 98, 100, -82, 103, 42, -126, 102, 124, -55, -56, -126, -33, 56, -81, 49, -1, 51, -70, -120, -120, 49, 25, 31, 112, -80, -82, 90, -15, 8, -19, -8, -80, 107, -91, 85, 7, -14, 28, 106, 2, -54, -54, 50, -86, 12, 105, 117, 32, 67, 69, 6, -111, -4, -31, -8, 118, 58, 107, -71, 13, -82, -66, 6, -42, -97, 39, 48, 65, -107, 50, 92, -29, 27, 126, -46, 14, 2, 82, -20, 14, 72, 85, -112, -108, -96, -97, 115, -61, -9, 31, -26, -27, -62, 100, -109, 62, -95, 33, -127, 51, -32, 112, -105, -112, -14, -7, -112, 2, -34, 81, 36, -106, 8, -38, -52, -121, 46, -42, 50, 28, -72, 48, 34, -3, -118, 1, 55, -22, -58, 94, -69, 64, 68, -21, 121, 4, -3, -37, -55, 74, -14, 16, 114, 96, -117, 113, -114, -73, -6, -84, 68, -45, -20, 8, 124, -11, -88, 105, 20, -43, 31, -90, -18, 36, 84, 47, -26, -112, -44, 114, 13, 121, 48, 93, 68, -105, 110, 48, -97, 101, -16, 76, 46, 99, -81, -41, 29, -96, -25, 73, -104, 115, -18, -115, -7, 78, 4, -120, -33, 13, -16, -55, -72, -57, -16, 115, -2, 77, 3, -35, 54, 6, 10, -28, 20, -32, -7, -64, -46, 77, -110, -48, 127, -89, 3, -36, -30, 97, 55, -104, 43, -119, -30, -58, -51, -42, -62, -123, -32, 102, -80, 72, -37, -77, 28, 42, 108, 103, -40, 26, -26, 86, 20, 62, 79, -29, 6, -107, 97, -114, 82, -4, 116, 11, -87, -61, 44, -85, 25, 26, -10, 113, 27, -96, -54, -44, -109, -19, -98, 95, -98, -1, -55, 114, 113, 56, -27, -105, 25, -107, 126, 115, 74, 98, 72, 67, 56, 89, 20, 102, 22, 102, -23, 56, 56, -72, 121, -105, 47, -23, -19, -35, -75, -35, 64, -112, -74, -106, 61, -38, 89, 28, 3, -46, -12, 2, 5, -51, 70, -26, -58, 4, -27, 58, 77, -37, -32, -55, 20, -123, 70, 55, -36, 119, -11, -123, -42, 60, -84, 1, -74, -30, 44, -49, 118, 21, 93, 33, -58, 90, 49, 10, -68, 55, -11, 3, 16, 108, 75, 83, 81, 95, 114, 98, -49, -83, -44, 24, 72, 11, -38, 110, -106, 54, 50, -118, -74, 122, -24, 96, 122, 37, -45, -19, 30, -76, -73, 54, 121, -77, -90, -47, 28, 42, 28, 83, 107, 6, 76, -122, 106, -61, 53, 99, -123, 120, 48, -107, -84, 27, -38, -21, 55, -125, 120, 42, 122, -34, -90, 61, 109, 55, 38, -86, -46, -20, -57, 47, 54, 65, 112, -4, -6, -8, -105, -100, 124, -96, -74, 117, 52, -63, 48, 3, -36, 16, -97, -111, -32, 37, -63, -106, -40, 15, -83, -21, -19, 113, 86, -96, 45, 30, 104, 29, 69, -34, -15, 115, 64, -96, -76, -77, 23, 68, 90, 66, -106, -92, 83, -26, 72, -70, 119, -2, -97, 88, 69, -76, -109, 76, -84, 17, 9, 87, 24, 31, 95, -36, -42, -127, -73, -89, 122, 54, -58, 7, -59, 56, 61, -12, -71, -12, 24, -42, -30, 111, -95, 75, -113, -98, 96, -111, 117, 118, 121, 60, 87, 101, 19, -47, 41, 115, 70, 108, 3, -112, -84, 36, -120, 64, -75, -57, -89, 72, -4, -39, -46, -29, 70, 10, -48, -27, -21, -111, 77, 49, 16, -67, 36, -127, -126, -1, 73, 66, -92, 87, -8, -40, 80, 0, -97, -45, 89, 4, 24, 120, 94, -114, -82, 99, 46, -101, 121, 7, -72, 69, -16, -116, -79, 57, 59, 88, 91, -120, -14, -71, 15, 38, 124, -114, -37, 49, 125, 25, -56, -9, -7, 101, 117, -115, -85, -59, -24, 110, -113, 108, -11, -70, 13, 106, -128, 54, 51, -36, 97, -56, -8, -59, 64, 16, 86, -83, 31, 34, 44, 71, -62, 40, 86, -126, 27, 124, -86, 24, 0, 26, -50, 38, -111, 106, 12, -28, 94, -90, 27, -14, 126, 12, -82, -14, 16, 72, 1, 53, -122, -9, 115, -107, -40, -5, -16, -1, 47, 3, -121, -56, -27, -19, 23, -15, -27, -50, 37, -20, -46, -29, 55, 83, 74, 114, -59, -46, -96, -2, 114, 125, 51, 77, 41, 24, 54, 17, 42, 41, 72, 45, 44, 84, -45, 83, 49, 70, 127, 94, 115, 118, -53, -6, -58, -106, 33, 58, 62, -79, 53, 72, -29, -79, -95, -13, 107, -8, 63, 63, -7, 85, 44, 116, -83, -81, 110, -19, 113, 99, 105, -105, 74, -23, 74, 127, 66, 26, -83, 78, -62, -128, 49, 74, 66, 77, -27, -74, 5, -127, -65, 92, 113, -111, 110, -59, 103, 93, 108, -83, -10, -4, 27, 49, -38, -95, 43, -77, -50, -56, 16, 3, -60, -6, -63, 17, 64, 53, 39, 106, 104, 74, -98, -48, -118, -18, 74, -34, -26, -62, -47, -56, 3, 126, -87, -63, 100, -34, 61, -61, -123, 15, -47, -45, 63, 125, -120, 116, 33, -116, -75, -20, -79, 105, 6, -44, -31, 88, -10, -58, -56, -41, 73, 113, 18, -81, 54, 17, -123, -95, -11, -114, -102, -55, 0, -40, 22, -118, -49, -55, -121, 121, -64, 32, -21, 109, 102, 86, 24, 113, 72, 32, 95, -126, 28, -50, 61, -66, -3, -28, 79, 127, -103, 23, -46, 110, -71, 53, 65, -119, -37, -92, -103, 0, 18, -92, 111, 6, -75, -112, -92, 51, -103, -49, -52, -123, -63, -49, 82, 48, -6, -127, -22, -109, 46, 83, -89, -104, -12, -37, -42, 7, 32, 123, 84, -55, 42, 13, -82, -26, -91, -90, -114, -36, -115, -81, 118, -71, 79, 70, -77, -9, 56, 100, 75, -73, 89, 88, -74, 86, 57, -78, 55, 22, -52, 18, -118, -116, -91, 97, 98, -73, 57, 89, 13, 125, -127, -69, -26, -52, -64, -105, -115, -104, -4, 90, 91, 74, 111, 16, -51, -29, 66, -41, 112, -51, 43, -48, 83, 33, -15, -76, 7, -13, 16, 14, 58, -9, 78, -36, 47, 106, -15, -88, -40, -26, -101, 40, -41, 92, -50, -127, 35, -40, 103, 98, 113, -41, -38, 34, 24, 109, 29, -81, -36, -9, 17, 47, -45, 87, 66, 13, -7, 108, 2, -47, -69, -47, 24, 52, 6, -52, 63, 29, -106, 76, -40, 19, 27, 119, 115, -127, 110, 25, -40, 9, -68, 20, -70, 92, 123, 115, -23, 80, -11, 97, 24, -83, 88, 46, -118, -19, 112, -69, -62, 55, -66, -103, -36, 92, -88, -127, 63, -58, -128, -85, 84, -4, 92, -85, -30, -52, 58, 52, 32, 75, -16, 32, 92, 16, 13, -125, 80, 42, -26, -100, 21, -45, -3, -27, -85, 48, -61, -111, -43, -83, 91, 89, 107, 78, -90, 113, 83, -114, 31, 80, -24, 70, 44, 111, 17, -122, 70, -86, -62, -54, -47, -2, 116, -98, 23, -6, -1, 124, -88, 105, 92, 0, -8, 25, -62, 48, 19, -18, 35, -40, -32, 57, -92, -81, 53, 92, -36, -85, -23, 32, 36, -74, 94, -124, 117, -31, 20, 29, 112, 62, 38, 84, -21, 120, -76, -111, -16, 52, -42, 46, 13, 88, 102, -8, 5, -35, 122, -36, -128, -98, -2, -16, 114, 23, 35, 0, 120, 5, 23, 105, -107, -90, -107, 56, 36, 82, -15, -98, -128, -16, 58, -65, 35, -118, -6, -58, 56, 37, 20, -19, -51, 83, 6, 119, -89, 63, -7, -55, 89, -8, 105, 20, 118, 57, 105, -47, 26, -100, -92, -110, 124, -94, -68, -110, -110, 19, 61, -122, -22, 125, -7, 107, 123, -74, 73, 34, -12, -7, 83, -71, -60, -6, -32, -99, 117, 34, 44, 62, 119, -128, 109, -30, -71, 14, 44, -42, 17, -25, -64, -78, -66, -90, 10, -44, 63, -43, 29, -16, -69, -51, -41, -37, -121, -32, 5, -17, 81, 38, -87, 70, -68, -57, -105, 57, -125, 32, -94, 56, 62, 39, 78, 49, 43, -61, -71, -89, -75, -102, -108, 120, 78, 109, -68, -19, 106, 76, 26, 107, -23, -33, -117, 68, 59, -52, 12, 67, -70, -63, 61, 72, 120, -110, 115, -30, -121, 102, -47, -116, 14, -44, 119, 8, 2, 32, 16, -59, -59, -33, -24, 64, 95, 89, -78, 54, -64, -45, -100, -106, 20, -61, -97, -96, -54, 74, 75, 111, 91, -2, -88, -4, 18, -45, 17, -55, 103, -34, -88, 109, 70, -87, 69, 78, 126, -124, 75, -60, 73, 89, -10, 30, -57, 24, -25, -23, 72, -112, 82, -44, -71, 54, 27, -88, -12, 107, -46, 103, -119, -69, -121, -89, 104, 126, 62, 85, 89, -78, 76, 88, -95, 26, 65, -4, 108, 77, -25, -8, 89, 9, -122, 91, -77, -28, 43, -16, 125, 126, -73, 17, -85, 30, 9, 13, -14, 67, 18, 21, -42, -91, -20, 93, -89, -76, -44, -112, 123, 21, 1, -100, 6, 56, 24, 111, 20, -116, 29, -65, 16, -75, -58, 99, -99, 4, -54, -116, 35, -121, -53, -71, 96, 79, 3, 21, 112, 102, -70, -83, -32, -36, -98, -81, 81, 112, -24, 91, 19, 48, 76, -88, 71, -43, 113, 13, 72, -13, 11, -88, -83, 49, -76, -47, -62, 112, 9, -26, 72, -3, -103, 64, -49, -55, -82, -127, -72, -46, -18, -23, -24, -38, 108, 27, -87, 78, -10, 52, 19, -15, -102, 41, -124, 99, 33, 49, 47, -59, -17, -46, -47, 54, -17, 114, -94, -55, 79, 118, 106, 94, 78, -10, 94, 37, 18, -70, 0, -34, 41, -56, -32, -86, -42, 58, -26, 75, -38, -76, -68, -111, -122, -34, 109, -22, -25, -73, -101, 116, 62, 103, 67, -33, -1, -49, -100, 11, -2, -103, 84, -26, 83, -91, 99, 2, 70, 86, 67, 121, 118, 64, 25, -115, 120, 86, 40, -69, -125, -121, 30, 9, 7, -42, -32, 10, -57, -78, -123, 56, 7, 40, 123, 109, 68, 100, 66, 56, 110, -125, -112, -78, -19, -20, 71, -21, 22, 63, -50, 57, 0, -68, -1, 127, -12, -4, -107, 75, -44, 35, -104, 26, -60, 63, -111, 88, -77, -19, 72, 74, -125, 24, 78, 59, 94, 73, 13, -38, -18, -64, -26, 89, 54, 110, -66, -59, -55, 99, -96, 110, -19, 37, -117, -88, 80, 13, 90, 116, -65, 123, 81, -83, 56, -77, 59, 54, 75, 89, -67, 79, -117, -81, -43, 35, -112, 123, -97, 89, 115, 3, 115, 99, 87, -97, -87, 8, -75, -116, -64, 29, -76, 87, 76, 119, -44, -91, 100, 107, 12, -47, 100, 51, 43, 78, 75, 25, -113, -118, -8, 123, 11, -36, -57, 118, 1, 32, -66, 107, 13, 93, 33, -92, -44, -73, 61, 26, 104, 91, 8, -119, 124, -125, 48, 112, 123, -18, 97, -41, 32, 17, 42, 35, 125, -124, 127, -111, 120, 100, -94, 117, 59, -112, -99, -25, -34, -58, -89, -30, -69, -116, 33, 115, 78, 2, -101, -4, 83, -33, 11, 20, 16, -112, -84, -90, -121, 119, -69, -70, 97, 31, 6, 11, 46, -112, -16, -53, 109, -94, 61, 51, 14, 112, -124, -89, -72, -66, -63, -41, 122, -19, -64, -100, 53, 125, 38, -85, 44, 126, 98, 107, 76, 32, -35, -79, 73, -58, -33, 51, -79, -81, 79, 29, 122, 55, -88, -17, -98, 88, -91, 62, 5, 23, 100, 114, -39, -115, 31, -71, -60, -30, 108, 115, 122, 58, -77, -99, 5, 115, -53, -18, 43, -51, -49, 3, 15, -93, -24, -49, 111, 43, 122, -102, -10, -16, -123, 36, 29, 42, -41, -8, -47, -20, 72, -68, 39, -24, 59, -121, -52, 123, 114, -126, 11, -20, -87, -71, -127, 42, -90, 83, 84, -115, -41, 95, 104, -9, 92, -79, -48, 6, -15, -37, -49, 50, -61, 120, 26, -120, 105, -73, -104, -88, -85, -1, 99, -75, -57, -114, 45, 81, 111, 39, -90, 86, -103, -82, -16, -42, 85, 105, 17, 39, 126, 88, -19, 99, 42, 46, -42, 68, -126, -121, 46, -73, -52, -47, -20, -13, -117, 112, 60, -74, 52, 116, -28, 124, -60, -55, 36, 46, -123, -118, 18, -16, -36, -105, -6, 22, 89, -70, 108, -100, 96, 86, 91, 16, 6, 100, -55, -31, -13, -69, -13, -4, 43, -9, -72, 16, 84, -56, 98, -37, 8, -20, -83, -49, -15, -8, 74, 8, -81, 1, -22, -118, 97, -56, -92, -12, 20, 33, 28, -88, 28, 57, 9, 117, 118, 52, -48, 36, 112, 110, -35, 32, -60, 89, -43, -121, 47, 27, 102, -74, 92, 53, 12, 64, -26, 52, -25, -5, 121, 79, 123, 52, 117, 33, -39, 4, 76, 20, -36, -104, -13, -6, 23, 124, -106, -31, -71, -37, -65, 89, 101, 69, 31, 89, -105, 61, 105, -42, -126, -40, -28, 55, -52, -40, 88, -1, -22, -6, 46, -28, -72, 126, -55, 109, 72, -4, -23, 7, -52, 99, 1, 13, -49, 104, 45, -48, -82, 59, -42, -37, 0, -1, 32, 25, -42, -86, -48, -4, 20, -84, -13, -30, 49, 66, -69, 95, -127, -5, 79, 72, -79, 52, 32, 46, -24, -100, 48, -125, -36, 22, -6, -26, -10, 90, -31, -37, 107, 20, 66, -60, 1, -14, 47, -124, -6, -4, -59, -70, -105, 7, -119, 69, -127, 40, 67, -49, -16, 28, -18, -21, 31, 65, 23, 21, -21, 87, 77, -30, -75, 108, -115, 52, 59, -25, -7, -73, 60, -87, 61, -125, 65, 19, -122, -7, -73, -57, -3, 42, 122, 106, -115, 111, 5, 40, -90, 125, 112, 14, -116, 74, -1, 21, -43, 36, -41, 102, -68, 49, 50, 55, -128, 50, 68, -108, -117, -87, 29, 11, -59, 96, -10, 105, -5, -69, -47, -76, 37, 109, 89, -38, 92, -46, 115, -115, -1, 3, -53, 2, 1, -61, -114, 23, 29, 121, 42, 56, -128, -46, 100, -99, -81, -46, 14, -41, 98, -118, 110, -124, -32, 4, 62, -96, 75, -44, 99, 111, -67, 69, 27, -86, 115, 115, -14, -66, -18, -4, 100, 71, 17, -82, 11, 97, 70, -91, 113, 9, -66, 75, 72, -2, 84, 79, -6, 95, 3, 62, -63, 107, 6, -52, -99, 70, 98, 39, 111, -50, -121, 91, -39, -38, -116, -68, -29, -55, -24, -127, 61, -83, 88, -28, 88, 111, 34, -7, -26, -97, -60, 32, 85, -42, 78, -16, 44, -50, 73, 114, -32, -76, 37, 79, -33, -101, 71, -91, -85, -38, -126, -102, -44, 16, -40, 112, 89, -91, -107, 96, -53, 57, 24, -46, 81, -95, -38, 62, 53, -4, 95, 108, -70, -13, 12, 125, -86, 33, 103, -90, -15, -97, -15, -64, 78, -36, -111, 1, 52, 115, -35, 35, -68, -82, 51, 51, 22, 10, -61, -118, 29, -57, -11, 72, -88, 119, 103, -9, -28, 31, -125, -54, 98, -102, -14, -42, 56, -42, 81, 96, 39, 33, -73, 59, 16, 107, -41, -109, 51, 10, 48, 36, 6, 81, -56, -12, -5, -107, -71, -116, 105, 94, 75, 110, 26, 123, -123, -12, 100, -66, -74, 71, 10, -101, -31, 65, -106, -94, -27, -98, -25, 7, -76, 58, -55, 119, -103, -25, -52, -52, 70, 51, -70, -5, -43, 64, -3, -77, -77, 107, -9, 91, 116, -52, -48, 43, 103, -41, -98, 106, 104, -105, 19, 108, -84, -116, 108, 61, -12, 124, 18, -94, 10, -33, 113, 93, -82, 92, -100, -54, 123, 104, 8, -82, 62, 123, -76, -40, 56, -92, 104, 90, -118, 92, 102, -80, 89, -44, -127, 19, 10, 56, -50, 68, 16, -13, 66, -54, -79, 109, -106, -76, -114, 59, 51, 97, 99, -101, -5, 35, 79, 107, 50, 10, 90, -95, 95, -40, 103, 58, -44, 107, 64, -9, -43, 106, 67, -90, -127, 14, 87, -57, -21, -56, -90, 51, -65, -44, -116, -125, 124, 41, 83, -6, -30, 110, -105, 39, 105, 102, 125, -98, 2, 75, -86, -32, -87, 39, -56, 81, -84, -97, 75, -89, 39, 58, -14, -120, -77, -11, -10, -36, -24, -12, 121, 54, -87, 2, 8, 52, 96, -32, -91, -92, -127, 118, -117, 127, -38, -102, -95, 108, 88, 17, -44, -5, -30, -33, -100, -126, -57, -74, 101, -9, 85, -65, -69, 49, 21, 89, 28, -62, 36, 36, 3, -61, -56, 26, 80, 22, -99, 41, 70, 102, 16, -114, -108, -116, -92, -32, -55, -104, 87, -43, -50, -32, -19, 26, -50, -110, -63, -33, -70, 76, 47, -76, -125, -24, 86, -15, 74, 9, -105, 9, 24, -50, -104, -17, -21, -101, -18, -33, -79, -69, 13, 76, 120, -8, 81, 74, 8, 33, -49, 36, -73, 61, -102, 81, 97, 103, -30, -123, -29, -32, 72, 112, -45, -68, 116, 48, 64, -97, 2, -118, 54, -25, 81, 22, 9, 101, 4, 13, 66, -27, -58, 34, -40, -38, -104, 37, -5, -124, 77, 44, -57, -34, 9, -87, -59, 29, -121, -5, -81, -102, -123, -121, -113, -126, 60, 115, -108, 44, 127, -58, -61, 87, 87, -113, -7, -99, -77, -12, -58, 77, -29, 113, -72, -98, -27, -52, -88, -11, 55, 61, -26, -11, -12, -6, 72, 56, 125, -3, -37, 47, -19, -52, 59, -20, -107, -83, -34, 107, -90, -61, -29, -8, 20, -92, -70, -109, 96, -109, -4, 21, -125, 45, -17, -103, -125, 16, 62, 14, 28, -99, -117, -5, -74, 117, 0, -15, -51, -69, 69, -57, 79, 50, -13, -128, 85, -32, 54, 39, -91, 41, 90, 52, 123, 5, 40, -107, 20, -103, -79, 96, 17, -50, -18, -25, -32, 25, 17, 44, 99, -101, -15, -93, 32, 54, 9, 23, -83, 2, -12, -44, -32, 79, 116, -118, -116, -53, 31, 113, 55, 109, -54, -23, 0, 115, 67, -100, -43, 20, 9, 3, -47, 102, -38, -95, 92, -97, -14, -50, -113, -8, -95, -91, 127, -93, -49, 69, 112, -119, 28, -66, 97, 71, -88, 80, 126, -68, 98, 37, 106, 18, -12, 22, -30, -62, 40, -87, -99, -7, 50, -33, 37, 88, -26, 9, 99, -100, -122, -58, 24, -94, 74, 2, 127, 71, 94, 52, 39, 69, -10, 34, 10, -98, 97, 7, 21, -32, -74, 58, 69, 39, 84, -68, -22, 24, -59, 1, -124, -127, -68, -88, -40, 68, -39, 24, -87, 70, -53, -96, -79, -67, -3, -58, 88, -48, 126, -5, 71, -41, -43, 96, 53, -86, 8, -11, 104, -111, 49, -38, -1, -79, 124, -19, 110, -112, 12, -120, 72, 30, 77, -70, 49, 110, -15, -23, 120, -79, 122, 50, -9, 48, 95, 123, -31, -62, -126, -116, 20, -17, -57, 78, -125, -12, 106, -37, 23, 39, -10, 34, -20, 127, 118, -111, -89, 127, -25, 28, 102, -77, -74, -106, 75, 34, -72, -116, 89, -31, 112, -103, 124, 20, -90, -124, -119, -57, -33, -45, -115, -87, 68, -100, -29, 31, 29, -51, 29, 80, -35, 119, -113, 35, -116, -10, 14, 87, -20, 67, 55, 23, -120, -8, -66, 115, 34, -12, -127, 66, 60, 0, 94, 39, -75, -51, -8, 50, -45, 56, -77, -111, 77, 9, -18, -23, 41, -56, 22, -111, -79, -2, 98, 33, 21, 105, 19, -50, 77, 72, -2, 82, 19, 4, 82, 36, 47, -109, 88, 121, 42, -109, -53, -85, -34, 41, 99, 25, -28, 31, 98, 104, -69, -73, -47, -22, 72, 60, 90, -14, 65, 121, 11, 80, -68, 21, -124, 77, 66, 109, -44, -39, 76, 118, -115, -12, 125, -4, -30, 108, -126, 97, 99, -118, 60, 13, 27, 109, 65, 117, -88, -45, 11, 126, -41, 34, -28, 50, 62, 93, 83, -72, -36, 94, 81, 37, 34, -58, -7, 116, 22, 9, -33, -22, 110, -40, -98, 121, -55, 5, 54, -6, 104, 17, -118, -1, -62, 0, 41, -12, 52, -107, -118, 30, 114, 6, 21, 112, -32, 102, -96, -70, 104, -78, 18, -10, -56, -25, 18, -76, 89, -32, -79, 49, -84, 93, -7, -96, -7, -57, 78, 114, -112, -13, -12, -42, 46, -122, 115, -33, -76, 12, -71, 39, 97, 116, 72, -125, 15, -35, 51, -62, 49, 37, 34, 70, 6, 9, -5, 76, -19, -126, 102, -93, 92, -86, 111, 52, -21, 24, -45, -50, -122, -109, -80, -29, 39, -30, -5, -74, -53, 12, 80, 16, -57, -46, 122, -128, 10, 26, -28, 3, 77, -38, -50, -112, -10, -1, -97, 125, 81, -18, 124, -27, -67, 2, -18, 89, -56, -115, 52, -80, 55, -21, -55, 97, 15, 25, -102, 117, 15, 9, -30, 35, -116, -56, 121, -4, -23, 8, -119, 78, -92, 7, -7, -121, -119, -86, 111, -6, -121, -61, 26, -122, -91, -81, -44, -17, 25, 46, -82, -65, 97, 46, 46, 84, 27, 38, 70, -26, 101, -71, 122, -34, 12, 10, -20, 70, -59, -48, -4, 101, 59, 2, 16, -104, 118, 116, -73, -100, -90, 127, -52, -105, 68, -40, -41, -74, 57, 95, 101, 15, 116, 51, -116, 31, -110, 59, -59, 26, -78, 106, -103, 28, 98, 90, 58, 36, -35, -97, 38, 75, 68, -65, 106, -42, -121, 74, -63, 118, -24, -55, -99, 24, -91, 84, -11, 26, -37, 89, -69, -35, -47, -61, -77, -121, -47, -14, 117, -30, 120, 43, 105, 70, 89, 42, 126, -101, -4, 8, -54, -107, 30, -127, 25, -125, 81, 24, -54, 46, 87, -126, -115, 12, -45, 27, -126, 76, -81, -55, 60, -65, -70, -33, 87, -128, 48, 102, 25, 58, -42, 90, -76, 94, -55, -29, 21, 30, -61, -18, 56, 97, 85, 1, -38, 93, -31, -25, -33, 4, 24, 41, -109, 4, -46, 37, 7, -13, 86, 39, 67, 31, -100, 89, 117, 123, 57, 124, -1, -104, 123, -53, 103, -119, 82, 35, -123, -20, 89, 34, -95, 56, 48, 19, -90, -33, 22, 78, -55, -44, 65, -78, 106, 117, 21, 10, -90, -128, 126, -80, -87, 115, -84, -45, 94, 5, -112, 10, 4, 9, -84, 118, 60, 3, 33, -60, -68, 82, -62, -118, -50, 48, 41, -55, 73, -85, 83, 38, 115, 120, 86, -101, -38, -104, 52, 21, -69, -31, -68, 67, -106, -65, -63, -69, -50, 53, -68, -26, -119, 86, 76, -124, 107, -87, -62, -56, -48, 14, -109, -74, 100, 53, -128, -114, -35, 11, -8, -77, 43, -82, -97, 52, 62, 98, -116, -40, 41, 64, 59, -121, -81, -10, 97, 96, -120, -87, -84, -74, 33, -88, -41, 61, -1, 40, 82, -77, -55, 21, 120, -92, 96, -33, -83, -11, 83, -98, -9, -102, 110, -115, 126, -17, 113, 73, 29, -30, 48, -109, 36, -117, -85, -41, 74, 126, -34, 54, -100, -88, -97, -120, -111, 85, -109, -39, 0, 106, -100, 102, 54, -66, 29, -101, -96, -61, -87, -65, -95, -117, -94, -39, 62, 50, 21, -39, -31, 41, -124, 20, -87, 8, -4, 26, 75, 15, 81, 113, -103, -25, -41, 88, 73, -111, 1, 108, -69, 91, 31, -114, -123, 113, 48, 96, -83, 69, 11, 12, -16, 109, -13, 12, -34, -21, 110, 112, -23, -80, -88, 2, 38, 84, 92, 19, 70, -110, 98, -9, -89, 95, 33, -57, -38, -77, -88, -79, -127, -121, -116, -63, -114, 34, -23, -100, -64, -2, 14, 92, 88, -101, 75, -91, -46, -12, 104, 39, -114, 62, 83, 45, -46, 15, -26, 17, -52, 77, -49, 93, 23, -46, -42, 1, -27, -82, -125, 119, 127, 99, 85, 101, -11, -50, 62, -89, -98, -15, -23, 66, 69, -24, -98, 122, 1, -56, -88, -83, -105, 62, -85, 117, 67, -47, -125, 83, -50, -128, -23, 19, 28, 107, 73, 73, 121, 116, -109, 11, -3, -84, -9, -47, 101, 110, -23, 68, -15, -14, 54, 24, -37, -30, -26, -4, -102, 105, 49, 108, 46, 57, 75, -91, 40, 86, 9, -1, 8, 18, 34, -72, 102, 96, 97, 68, 77, -32, -61, 90, 122, 122, -67, -87, 61, 78, 81, 122, 63, -28, -113, -14, 30, -8, 79, 3, 92, 76, 12, -47, -98, -112, -25, 83, 64, 127, 91, 28, 35, 127, 23, -51, 78, -118, -52, 91, -127, 80, 65, 85, -62, -25, -108, 16, 9, 65, 65, 10, 68, -107, 41, 85, 16, 24, -68, -86, -71, 120, 81, -73, 32, 90, 67, 125, -120, -9, 105, 27, 2, 104, -41, 109, 9, 83, 126, -57, 89, -108, 61, -56, 67, 125, 73, 96, 114, -79, 104, -51, 33, -85, 82, -64, 105, 62, -104, 9, 97, -77, -110, -80, -107, 31, 3, 13, -25, 62, -56, 110, -35, 19, 84, -81, -5, 80, 8, -20, 94, 59, -117, 43, -67, 110, 43, 112, -108, 109, 90, -109, -114, -48, -60, 64, 4, -92, 8, -53, -114, -24, 14, 31, -37, -117, 112, 99, 81, 22, 98, -82, -13, 115, -122, 18, 99, -85, -31, 19, 39, 90, -29, -66, -34, 50, -103, 125, 34, -87, -80, -81, 67, -41, -25, 19, 1, 123, 102, 50, 53, 66, -111, 78, 8, 110, 67, 39, 98, -118, 114, -62, 48, 19, -55, 4, 41, -94, 62, 64, -56, -32, 95, 53, -111, -87, -8, 3, -54, 10, 13, 103, 63, 40, 109, 31, 30, -96, 64, -21, 16, -23, 0, -65, 19, -114, -115, 112, 57, -128, -63, 74, -87, -125, -117, -94, -8, 95, 46, 37, 12, 81, -109, -9, -102, -58, -87, 8, -83, -11, -74, 11, -66, -26, 57, 64, -66, 82, 91, 40, -18, 83, -57, -9, 44, -92, -75, 85, 36, 84, 36, 44, 78, -46, -89, -2, 87, 18, 89, -101, -111, -93, 117, -103, 105, -20, -23, -8, 54, -57, 79, 97, -112, -29, 27, -53, 12, -105, -82, -100, 72, 46, 10, 92, -91, 48, -47, -52, 81, -33, 8, 76, -45, 111, -29, 48, -36, -8, 105, 51, -15, 105, -113, 71, -25, 51, -68, -91, -52, 53, 50, -72, -115, -4, -109, -32, -99, -112, 77, 102, 107, -75, -83, -28, 16, 39, -92, -25, -48, -104, 88, -83, -65, 22, -98, 31, 122, -116, 103, -63, 13, -29, -55, -46, 105, -15, 73, 101, 59, 114, -49, -50, 95, 122, -63, -116, -76, 90, 62, 6, -45, 9, 102, 65, 46, 26, 29, 124, 87, -75, 85, 69, 94, 83, -106, -5, -27, 29, -114, 118, -88, 17, -109, 99, 76, 41, 30, 91, -59, -122, -90, -99, 58, 121, 10, -86, -106, 24, 119, 48, 92, 116, -93, 49, -64, -100, -68, 31, -18, -22, -20, -57, 74, 32, 115, -62, -111, -11, -110, -49, -81, -120, 56, -50, 92, -60, 21, -127, 7, -87, 93, -31, -54, 4, 50, -96, -44, 79, -85, 1, 79, 107, -125, 44, -113, 26, -33, 23, -125, 91, 117, 15, 74, 102, -90, -97, -86, -7, 0, -114, -1, 64, -106, -44, -13, 48, -33, 90, 68, -80, -120, 32, -63, -93, 107, -12, 110, -100, -32, 47, 21, -115, -81, 97, -104, -118, 55, 51, 10, 111, 95, -69, -108, -69, 47, -47, -28, -23, -49, 50, 116, -47, 94, -78, -110, -56, 57, -36, -83, -54, 106, -79, -71, 74, -100, -92, -5, 110, 0, 0, 68, 4, 73, -3, 55, -15, 0, -78, -37, 119, 125, 77, -124, -11, 89, -80, -67, -93, -35, -54, -81, 92, 4, 32, -75, -99, -111, 102, -43, -59, 47, -84, -80, 61, 98, -69, 50, 11, -19, -127, 118, 81, 41, -34, -52, 31, -69, -30, 97, 86, -90, 57, -44, 36, -81, -126, -124, 123, 4, -110, 6, -83, -106, -121, 95, -82, 96, -69, -54, 11, 25, 125, -67, 82, -109, -6, 53, -1, 100, -78, -80, 98, -66, 6, -18, -68, 25, -19, -68, -51, 127, 89, -41, 69, 68, -88, 103, 27, 17, -93, -54, -97, -29, 56, 16, 45, 74, -112, -21, 79, -9, -109, -19, 122, 89, 115, -98, -127, 24, -49, 24, -84, -86, -70, -13, -107, 42, 91, -46, -41, -117, 111, 1, -68, 50, 105, 21, 71, 59, -115, -62, 101, 63, 29, -33, -71, -63, -102, -92, 18, -10, -88, 23, 20, -105, -32, -74, -75, -65, 55, -67, -18, -18, 70, 116, -95, 89, -105, 44, 59, 92, -24, 46, 104, 19, 60, 88, 49, 19, -39, 46, -72, 111, -94, 104, -108, 26, 99, 41, 98, -85, -64, -120, -78, -99, -71, -17, 25, 94, -38, 39, 25, -49, 59, -25, 39, -77, -29, 96, -35, -38, -92, -123, 1, -113, 121, 64, 118, -1, -128, 94, 7, 69, -92, 25, 94, 127, -29, 111, -33, -78, -95, -96, 61, 107, 118, 90, 91, 116, 120, -15, -121, -31, 62, -37, -64, -45, 61, 73, 83, 88, 0, -66, -43, -109, 35, 63, -57, 121, -63, -103, -72, -5, 110, 12, -50, 70, 41, -92, -21, -22, -60, -47, -108, 44, -8, -31, 123, 1, 66, -35, -73, -101, -3, -58, -58, 45, 72, -55, 119, 48, -81, -113, -115, -23, -22, 127, -65, 53, 70, -125, 47, 17, 94, -47, 12, -125, 43, 66, -4, -33, -26, -123, 9, 49, -117, -107, -123, 18, -97, 78, 46, -111, -36, -2, -116, -63, -91, -44, -54, 5, 26, -70, 75, -46, -59, 87, -66, -5, 107, -82, 126, -78, 21, -19, -29, 14, -8, -107, 117, 70, 97, -12, -16, -4, -25, -97, 94, 25, 45, -63, 108, 14, 20, -21, -54, 25, -45, 2, 5, -41, 28, 49, 71, -68, -40, -14, -8, 74, 67, 43, -63, -86, -22, -61, -93, 39, 46, -29, -75, -77, -79, 25, -65, -86, 107, 86, -28, -9, 55, 27, 3, -90, 37, 7, 120, -109, -110, 22, -1, 50, -30, -12, -89, -29, 18, -71, 71, 41, -126, 110, -12, 58, 12, 74, -77, -100, 111, -128, 105, -24, -93, 49, 123, -70, -104, 15, -59, -113, 116, -106, 87, -76, -10, 68, 56, -125, 99, 43, 67, 120, -24, -49, 23, 52, 113, 99, 21, -31, 54, -113, -54, 67, -92, -45, -54, 112, 88, -84, -48, -56, -98, -106, 46, -97, 29, -25, -20, -96, 67, 121, -80, 83, -81, -128, 112, -35, 5, -112, 86, 81, 5, -59, -18, 111, 53, -91, -116, -100, -70, 17, -59, 105, 94, 14, 33, -14, -105, -27, 22, -120, 108, -110, -128, 52, 86, -21, 56, 125, -14, 43, -117, -67, -13, -31, -2, -68, -112, 76, -54, -118, 114, -44, 82, -118, 91, 38, 117, -4, -86, 75, -49, 86, -107, 82, 113, -74, 97, 97, 19, -120, -46, 61, 91, 102, 94, -127, 0, 38, 45, -115, 110, 114, 80, 96, -52, 28, 3, -17, -52, 6, 10, 22, 19, -119, -128, 50, -125, 91, 10, 4, -50, -32, 64, 86, -60, 84, -1, 103, 111, -62, 61, 14, -125, -116, -103, 2, 38, 22, -106, -120, -128, -126, 67, -44, -98, -126, -106, -9, 40, -18, 70, 49, -94, -78, -85, 118, -120, -11, 30, 52, 60, 59, -81, 3, 103, 114, -31, -50, -82, 118, -82, 25, 84, 124, -41, -20, -107, 80, -125, 5, 90, -103, 98, -44, -26, -104, -113, 91, 34, 79, 100, 50, 27, -65, 86, 124, 91, 36, -43, -63, 66, -83, -1, 18, 45, -114, -86, 35, -116, -101, 20, 86, -115, 9, -84, -96, -81, 28, 83, 2, -14, -64, -15, 69, -22, -98, -55, -1, -26, -128, 81, 37, 20, -30, 103, 85, -69, -29, -30, 16, 23, -92, -53, 73, 91, 99, -75, -94, -53, -15, -73, -127, 83, 123, -110, -5, -45, -9, 15, -65, -88, -115, 61, -83, -96, 22, 39, -31, -126, -73, -83, 77, 38, 91, -124, -65, 41, 94, -78, -87, -7, -121, 60, 41, -14, 29, -123, -52, -84, -18, 6, 20, -97, -101, 116, -75, 26, -88, 49, 40, -26, 26, 49, -17, 38, 125, 62, 11, -10, -38, 76, -52, 72, 65, -83, -3, 62, 27, -21, 18, -48, 5, -32, -121, -20, -49, 48, 93, 22, 95, 95, 79, -29, -81, 87, 114, -5, 83, 35, -53, 64, -36, -117, -105, -52, -27, -109, -106, -82, 69, 69, 83, 34, 126, 10, 118, -53, -90, 55, -56, 95, -2, 59, -117, -112, -21, 5, 19, 0, 78, 38, 22, -58, 82, -117, -22, 40, 109, 18, 38, 30, -128, 17, 73, -93, 74, -78, -16, -72, -48, -12, -67, 107, -79, 47, 127, 84, -109, 67, 83, 108, 30, -81, -62, -2, -98, 97, -13, 14, 46, 9, -34, 68, -84, -81, 92, 31, -105, 125, 107, 94, 54, -62, -90, 7, 126, -48, -112, -28, 51, 41, -120, -18, -6, -102, 96, -102, 36, 5, 56, 28, 101, -122, 0, 11, -63, -114, -54, 69, -88, 62, -100, 113, -6, 40, 32, -120, 121, -86, 78, 41, -59, -103, -38, -65, 99, 25, 47, 105, -16, -98, 62, 53, 45, 42, -15, 39, -47, 77, -30, -19, -124, -82, 45, 99, 64, 1, -110, 55, 70, -60, 87, 23, 32, -35, -93, -51, -47, 84, -65, -45, -57, -88, -12, 77, -46, -112, -111, -84, -38, 36, -87, 90, -114, -70, -42, -37, -97, -78, -49, 19, 117, 107, 26, 118, 52, 38, 72, 110, 44, 100, -51, 110, 127, 83, -109, -26, 35, -8, 67, 8, -14, 41, 34, 15, -30, -60, 103, -89, 34, -81, 31, -95, 25, -105, 50, -112, -89, -53, 40, 68, 91, 4, 78, 30, -123, -111, 112, -74, -67, 75, -9, 24, -27, -9, 86, -122, 63, 88, 116, 85, 68, 75, -18, -21, 12, 13, 68, 21, -89, 105, 44, 11, 3, -17, -110, 88, 118, -54, 10, -76, 92, 36, -121, 65, -5, 15, 127, -88, 92, 22, 52, 13, -53, -60, -112, 107, 60, 13, -22, -27, 6, 11, 100, -58, 36, -112, -85, 72, -45, -52, 17, -2, -45, 89, -40, -5, -22, 43, -23, -97, -26, -49, 11, 10, -119, 45, -76, -85, -28, 119, -77, -90, -2, 80, 58, 78, 122, 29, 42, 16, -72, -104, -3, -63, -74, 38, -19, -81, 61, -18, 117, -71, 36, 10, -111, 35, 115, -86, -74, 57, -123, 81, 59, 16, 78, 67, 62, -80, 123, 12, -27, -20, 33, 100, 2, 60, 98, -9, 53, 121, 103, 28, 62, -83, -87, -91, -80, -16, -128, -104, 4, 26, 49, 19, -114, 109, -106, -69, -10, -100, 64, -8, -121, -123, 106, 90, 47, -104, 95, 52, 12, -68, -75, 126, -128, -48, -86, 63, -39, 70, -92, -27, -87, -119, 86, 116, -37, -25, 53, 10, -14, 106, -24, 8, -4, 45, -49, -36, 113, 125, -48, -12, -56, 8, -123, -71, 65, -8, 56, 127, 66, -18, 123, 64, 115, 107, 67, 1, 79, 65, -21, -54, 80, -124, -118, -107, -4, -124, -72, -10, 31, 2, -99, 54, -121, 10, 79, 75, 67, 95, -20, 121, -103, -41, -17, -15, -15, -44, 109, -60, 47, -68, -84, -7, -115, 54, 6, -91, -115, -60, 73, -111, -116, 19, -74, 73, 47, 14, -66, 40, -67, 90, 116, 50, -28, 78, 63, -13, -106, -54, -48, 0, 23, -110, 53, -63, -122, 89, -55, 92, -33, -7, 28, -2, -49, 58, 120, 69, -75, 109, 105, 76, 92, 7, -33, 26, -8, 95, 0, 21, -13, -118, -98, 7, 45, 101, 99, 61, -123, -70, -98, -53, 106, 5, 67, 16, -97, 52, -114, -94, 54, -6, 12, -127, -75, 123, 31, -22, 55, -41, 68, 57, 32, -104, -119, 104, -103, -118, -35, 12, -51, 38, -116, -57, 38, -24, 70, 19, -63, 87, -48, -106, 112, -112, -31, -40, 66, 26, -51, 52, -118, -51, -125, 75, -46, -114, -66, 38, -10, -8, 110, -123, -99, 9, 56, 0, -29, -48, 10, -32, -89, 79, -41, -58, -83, 33, 38, -111, 69, 51, -25, -10, -79, 62, 104, 36, -89, -102, -52, 73, 87, -29, -23, 45, 96, -16, 59, -87, -56, -100, 20, 48, 70, 44, -14, 25, 114, -123, 102, 49, 120, 11, -37, -45, 56, -109, -81, -12, -18, -19, 122, 111, 76, -49, 93, -95, -25, 52, -95, 40, -8, -117, -78, -110, 96, -91, 114, -59, 38, -113, -128, -55, -3, -10, -8, 11, -120, -123, 40, -77, -114, -101, -67, -100, -8, -102, 5, -64, -51, -57, 52, -42, -104, 25, -108, 126, 52, 36, 3, -126, -65, 97, 120, 94, 43, 109, 69, -111, -82, -30, 118, 36, -101, -48, 119, 110, 8, -1, -79, -35, -53, -105, -1, -85, 64, 1, -108, -68, -60, -86, -23, -6, -86, -80, -62, -121, 115, -18, 65, 107, -35, -55, -22, 61, -97, -111, -115, 18, -74, -49, 78, -47, 91, 92, 48, -47, -105, -48, 117, 16, -91, 123, 110, 108, -95, 52, 10, -96, -94, 86, 56, 66, 48, -35, 107, -6, -65, 90, -90, -45, -9, 100, 32, 124, 61, -8, -53, -5, 21, 14, -74, -107, 68, 113, -67, 36, -79, 20, -80, -67, -92, 37, 19, 5, -118, -95, 11, 74, 73, -122, 24, -114, -62, -2, -39, 36, 126, -14, 37, -12, 54, 21, -46, -37, 35, 88, 101, 28, 66, 35, 52, -116, -14, 23, 102, -21, -108, 16, -84, 14, 15, 65, -102, 125, 106, -48, 11, 34, -6, 81, -74, -128, 72, -66, 68, -43, -38, -18, -100, 26, 84, -29, -15, -10, 51, 51, 115, 54, 120, 17, 8, -115, -73, 30, 20, -90, -10, 103, -32, -74, 58, -5, -50, 14, 30, 77, -102, -61, -26, 82, -84, 101, -82, 108, 38, 127, -125, 22, -94, 56, -94, -115, -115, 36, 70, 59, -108, 46, -63, 71, -70, 71, -92, 115, -105, -94, 95, 71, -36, -67, 22, 54, -86, 127, -105, 28, -90, 18, -53, 56, 10, -10, 78, 99, 78, 0, -106, 22, 42, -92, -47, 24, 76, -67, -41, -3, -35, 60, 52, -35, -96, 41, -38, 106, -83, -14, 46, 121, 94, -26, 36, -57, 81, 98, -15, 107, 49, 12, -64, 60, 32, -10, 38, 73, -45, -64, -123, 38, -18, 87, 17, 112, 35, -14, 104, -126, -64, 85, 68, 56, -7, 103, -34, 46, 50, 122, -22, -27, -78, -55, -93, 114, 25, 87, -48, 6, -97, -92, -108, 9, 53, 36, 75, 107, -97, 32, 6, 122, -99, 114, -6, -37, -125, 50, 29, -50, 95, 111, 26, 13, -123, 51, 117, 14, 98, -70, -25, 112, -32, 117, -55, 124, 121, -112, 26, -37, -89, -81, -32, 40, -52, 100, -22, -36, 57, 33, 89, -104, 122, -46, -26, -91, 34, -110, 0, -100, 13, 67, 47, 73, -70, -78, -18, -61, -102, 77, -112, -39, 3, 90, -87, -109, -88, -87, -5, -4, -49, 55, 122, -86, -43, 17, -13, 11, -19, -65, -96, -60, 28, 120, 115, -47, 4, 18, -47, 70, -21, -73, -81, -100, -110, 41, -51, 77, 113, -118, -125, 102, -92, -87, 66, -47, 12, -112, 126, 105, -27, -38, -2, 46, 88, 43, -122, -126, 0, -125, -82, -128, -86, 83, -83, -62, -79, 34, 45, -40, 121, 65, -33, -4, 13, -90, 118, -55, -44, 13, 87, 102, -118, 50, -33, -6, -125, 72, 66, 67, -18, 35, 16, 116, -88, -87, -15, -87, -9, 101, -71, 56, 76, 99, 52, -117, 68, -23, -19, -26, -76, -96, 50, 72, 114, 57, -126, -72, 103, 104, -15, -50, -60, 0, 84, 15, -94, 34, -128, 120, -98, -22, -15, -22, -74, 93, -62, 85, 0, -107, 13, 79, 28, -70, -58, 105, -47, -65, 38, 20, -40, 124, 71, -19, -56, -83, 18, 90, 76, -41, 37, 25, -2, -58, -96, 8, 64, -98, 73, 13, 50, 97, 50, -118, -19, 46, -63, 12, -127, -23, 91, 50, 24, -16, 109, -102, 74, 30, 46, -19, -126, 78, 3, -10, 112, -107, -25, 122, 35, 32, 27, 84, 80, 1, -103, -33, -77, 20, 85, -97, -109, 44, 66, -118, -88, -123, 89, 72, -107, -76, -121, 67, 58, 22, -104, 70, -76, 87, -102, -7, -47, 39, 10, 123, 80, -119, 69, -28, 87, 57, -25, 28, 19, 80, -33, -112, 9, -30, -1, -49, 118, -19, -98, 112, 54, -82, 31, -93, 93, 53, 16, 38, 86, 14, 21, 13, 59, -109, -61, 58, -88, -89, -25, -84, 49, -117, -71, -127, -27, -90, 42, -8, 98, 85, -49, 70, -97, -98, -29, -55, 30, -105, -17, -15, 73, 115, -8, -97, -10, -8, 61, -51, 97, 88, 44, -17, -106, -23, 22, 102, -7, -71, 35, 86, -96, -81, 93, -112, -8, 79, 8, 48, 112, -60, 20, -18, -72, 124, 115, -40, 69, -90, 44, 98, -105, 96, 96, 98, -88, -100, 59, -36, 83, -2, -14, 123, 102, 33, -88, 2, -85, 39, -40, 74, 86, -75, -33, 60, -95, 84, -45, -105, -126, 29, 15, -105, 85, 75, 83, -61, 33, 76, 43, 121, 65, 66, 113, -67, 67, -26, -70, -65, 47, -83, 52, -32, -30, -26, 110, 68, 87, -44, 59, 68, 47, -25, 123, 65, -72, -90, 91, 89, -106, -33, 70, -78, -78, -117, -108, -26, 77, -21, -15, -31, -127, -18, 93, -39, 39, -30, -98, -91, 55, 116, 96, 52, 46, 120, -51, -128, 3, -16, -21, 36, -32, -44, -87, 69, 96, -16, -41, 93, -71, -88, 68, -23, -22, -88, 18, 43, -97, -73, -12, 8, -45, -37, -114, -28, 21, -93, -53, 22, 30, 72, 71, -41, 8, 115, 45, 113, 89, -34, -18, 102, -58, 51, 23, -59, -78, -117, -11, 109, 12, -102, 68, 120, -53, 2, -47, 93, -84, -56, 100, 117, -19, -37, -93, 110, -72, -18, -59, 27, 77, 115, 105, 79, -49, -4, -60, 89, -71, -116, -115, 7, 45, 9, 45, 4, -77, 38, -60, 26, -87, -116, 124, 67, 45, 52, 69, 36, 4, 64, 4, -70, 81, -94, 107, -51, 96, 17, -76, -44, 69, -34, 79, -11, 49, 109, -111, 75, -55, 57, -59, 25, 26, -47, 102, -111, -27, 47, -125, -66, 119, 96, -126, 44, 59, 119, 15, 124, -127, 32, -114, 0, 99, -122, 81, 11, -65, 62, -122, 19, 18, -53, 67, 43, 48, 99, 53, 59, 105, 108, -3, -84, 112, 50, -89, -108, -80, -47, -50, 53, 12, 13, -68, 64, 60, -75, -11, 38, 32, -90, 51, 29, 63, -122, 83, -22, -86, -11, -48, -67, 109, -113, -52, 8, 21, -71, 118, -83, 17, 49, 59, -108, 47, 49, -12, -80, 106, -64, -93, -61, -62, 78, 57, -114, 87, -47, 20, -113, 84, -91, -39, -69, 16, 0, -78, -89, 53, -81, 88, 100, -63, 56, 66, -94, 118, -65, 7, -102, 53, -8, 114, -54, 91, -25, 41, -23, -7, -111, -102, 68, 20, -119, -68, 1, -15, 44, -109, -28, -52, 113, -103, 5, 86, -121, -70, 25, 86, -51, 27, 25, -37, 106, -69, -17, -125, 3, 89, -126, -30, 20, 28, 33, 71, 25, -110, 109, -121, -108, 95, -62, -109, 22, 19, 98, 79, -51, -19, 105, 113, -43, -75, 59, -102, -74, 14, 124, -60, -88, 39, 105, 8, 90, -84, 67, -117, -68, -100, 12, -98, -23, -17, -49, 90, -77, 76, 76, 25, -19, -43, 121, 43, -40, -19, -123, 109, -24, 118, -112, 14, -115, 18, 70, 93, -6, 18, 6, -82, -49, 78, 65, 82, 127, 93, 105, -15, -94, -121, 82, -30, 84, -78, -52, -95, 78, 70, -59, -42, 117, -26, 35, -1, -28, -100, 86, -89, 67, -50, -48, 10, -9, -42, 6, -9, -107, -117, 111, 43, 32, 18, -14, -6, -11, -71, -92, -10, -49, 74, 51, 125, 42, 123, 37, -41, -63, -66, 4, 30, -90, -101, 119, -86, -123, 28, 78, -114, 118, 90, 8, 43, -1, -84, 18, 79, 7, -43, -11, 36, -21, -6, 28, -35, -97, -95, 18, 13, 71, -17, 53, 9, 34, 13, 73, 7, -11, -27, -68, -24, -28, -12, 2, 127, 47, 49, -46, -105, 19, -89, 41, -29, -106, 39, 40, -126, -111, 121, -115, -36, -124, 13, -64, 34, -109, -29, -86, 103, -98, -117, -7, -55, -89, 40, 67, -24, -122, -106, 38, -73, -95, -10, 108, 6, -97, -61, 97, 73, 63, 91, 102, -93, -84, -51, 58, 1, -110, -100, -29, -88, 66, -77, -25, 77, 65, 69, 31, 67, -47, 120, 85, -127, 119, -31, 64, -35, -111, -53, 119, 104, 118, -77, -2, 126, -8, 60, -85, 0, 100, -3, 115, -2, 78, -91, 100, 82, -75, -12, 11, -122, 123, 70, -57, -35, 80, 65, 0, -3, 26, -97, 111, -7, -43, 71, -92, -53, -108, 46, 98, 73, 112, 2, -38, 95, -127, 65, -31, -84, -109, -118, 31, 5, 70, 96, 25, 91, 88, 3, -41, -16, 109, -85, 96, 8, -124, -112, -27, 9, 36, -61, 90, 29, 8, 105, -115, -26, 76, -13, -114, 4, -11, -98, -31, 30, 40, -120, -82, -126, 61, 73, 126, 98, -62, -55, -17, -17, -71, -51, 105, 123, -76, -92, 109, 23, -89, -100, 90, 11, 64, 40, -103, -26, -14, 28, -59, -113, 54, -59, 103, 1, -121, 18, -18, -104, -43, 19, 60, -99, 28, 109, -73, 92, 115, 52, -5, -72, 118, 119, -19, 50, -106, 50, 75, 67, 117, 10, 99, -114, -42, 94, -114, 4, 18, -22, 14, -122, -111, 87, 118, 62, -69, -124, -84, -51, -88, 89, 87, 111, -53, -83, 105, -53, 82, -21, 49, 88, -96, 21, -87, 60, -29, -25, 59, -24, 6, -94, 24, 41, -84, -11, -7, -91, -8, -4, -56, 5, 65, -66, -29, 5, 18, -22, 43, 86, -53, 33, 84, -103, -40, -44, 92, -64, -41, -67, -44, 79, 54, 3, -64, 49, 15, -88, 74, -61, -97, 76, -74, -90, -65, -110, -64, -33, 120, 64, 87, -77, -125, -72, 17, -96, -72, 67, 103, 27, 72, 51, 65, -72, -30, 4, -19, -57, 32, -9, 114, -72, 26, 101, 2, 123, -91, -75, -8, 12, 36, 112, -57, -102, -16, 127, -94, 51, 16, 117, -58, 21, 79, 86, -60, 63, -86, -40, 104, 79, 71, 126, 57, -118, 36, 101, 62, -120, 28, 96, -42, 114, 20, 111, -112, -125, 23, -85, 29, -54, -99, -97, 89, -85, 25, -82, 124, -37, -56, -12, 115, -22, -107, -71, -113, 41, -126, -86, 100, 28, 12, -43, 104, -51, 113, -76, -24, 26, -95, -124, 69, 18, -20, -5, 36, 33, 11, 26, 102, 67, -113, 88, -34, 86, 48, 1, -95, -120, -21, 56, -79, 25, 24, 70, -14, 54, 62, 43, -50, -44, 89, -103, 20, -108, -90, 2, 8, -80, 84, -34, 92, -80, 115, -93, 30, 58, 53, -68, 56, -47, -65, 64, 36, 20, 59, -87, 68, -10, 47, 7, 109, 63, 122, 38, -39, 16, -117, 78, 39, 91, -73, -86, -42, 119, 73, 86, -111, 11, -117, 127, -53, -8, 44, -72, -101, -38, -9, -15, -84, 23, 55, -107, 39, 32, 37, 66, -35, -32, -100, 94, -15, 110, -100, -61, 23, 66, 45, 120, -101, 91, -75, 113, -103, -36, 101, -106, -125, 45, 121, -72, -30, -17, 31, -101, -66, 86, 113, -1, -23, 53, -89, -21, -93, 57, -20, -31, 51, 32, 5, 22, 86, -29, -107, 7, -8, 120, -38, 49, 21, 28, -98, -74, -34, -47, 54, -35, -83, 82, -97, 123, 62, 110, -6, -73, -52, 17, 52, -60, -120, -46, -90, -121, 58, 64, 103, -42, -48, 94, -57, -79, -25, -46, -6, 100, 4, -61, -96, -1, -71, 62, 1, 105, 77, -121, 61, 42, 89, -38, 66, -111, 37, 29, 20, 29, -109, -64, 16, -113, 36, 14, 79, -108, -82, -9, 3, 99, 109, -17, 62, -119, 81, -29, -32, -81, 121, 18, -41, -43, -74, 83, -49, -6, 80, 18, 69, -76, 83, 76, 3, -65, -3, 81, -42, -61, 14, 92, 58, -7, 37, 7, -99, 96, -122, 85, -74, -10, 32, -55, 40, -1, -40, -94, 114, 14, -66, -105, -74, -42, 43, 80, -88, -118, -43, -89, 7, 77, 127, 87, 73, -112, 110, 101, 67, 27, 40, 69, -4, -78, -67, -104, 104, 43, -34, 84, -23, 106, 46, -122, 97, -12, -51, -116, -82, 71, -52, -19, 22, -51, 56, -42, 85, -26, -82, 41, 17, -19, -33, -105, 108, -16, 15, -49, -64, -102, 100, 116, 40, 122, 124, 55, 67, -99, 80, -31, -90, 1, 27, 80, -105, 96, 103, -77, -84, 61, 43, 37, 80, -118, 110, 8, -106, 88, 59, -69, 46, 79, -114, -123, 56, 99, 67, -111, -45, 17, 67, 118, -61, 72, -89, -31, 64, -30, -65, 62, 57, 49, 73, -12, 35, 81, 12, -43, -89, -58, -105, 74, -45, -120, -89, 10, 107, 80, -32, -4, -3, 18, -26, -80, -46, 102, -116, 113, -36, -105, -92, 112, -48, 104, 17, 49, 116, 31, 101, 47, 20, 108, -35, 100, -86, -124, 48, 78, -118, -117, -18, -12, -41, 27, -92, 112, 124, -1, 56, -91, 21, -80, -27, -115, 40, 8, -71, -102, 50, 78, 99, -64, 72, 111, -46, 65, -75, 32, 52, 61, -6, -60, 109, 93, -99, -52, 69, 60, 39, -77, 120, 82, -81, 45, 1, -121, 31, 47, 113, 14, 126, -118, -72, -92, 11, -61, -6, 113, 18, 10, 33, -96, 13, 28, -74, -17, -74, 82, 39, 71, -116, -34, -24, -17, -51, -100, -99, -95, -111, 101, 9, -122, 64, -72, 127, 29, 105, 123, 20, 3, 20, 104, -120, 4, 108, -79, -110, 125, 90, -38, 82, 48, 4, 32, 116, 100, 50, 125, 98, -96, -84, -50, -107, 71, -46, 40, 85, 74, -45, -105, 91, -107, 40, 28, 70, 34, 73, 96, 68, 123, -112, 82, 87, 65, 115, 108, -111, -47, 67, 74, -23, 123, -13, -85, 66, -77, -13, -117, -69, 64, 39, 90, -118, -96, -95, 16, 24, 120, -101, -12, 44, 113, 91, -21, 126, 29, -60, 73, -73, -39, -110, 53, 40, 116, 49, 56, -35, 49, 102, -16, -99, 10, -3, 64, 24, 45, -103, 33, 83, -72, 23, -8, -96, -35, 115, -92, 21, 44, -22, -126, -47, 73, -37, -25, 75, -72, -95, -31, 65, -45, 109, 54, -118, -42, -107, -37, 90, 112, 82, -59, -96, -125, 72, -123, -74, 57, -112, -26, -25, -121, 31, 111, -79, -98, -111, 15, -92, 26, 0, 49, -36, -22, -116, 83, -1, -64, 110, 75, 126, 86, -91, 48, 48, 42, -35, -52, -75, 109, 22, 46, 16, 11, 50, -105, 4, 75, -95, -118, 37, 51, 108, 60, -77, 104, 12, 41, 32, -2, -64, -43, -13, 85, 62, -1, 109, -60, 92, 45, -32, -126, 7, 74, -77, 17, 68, -58, -117, -73, -57, 21, 70, -84, 65, 4, -76, -101, -7, -82, -85, 92, 40, 8, 13, -46, -12, 99, -60, 107, -45, -94, 64, -17, -110, -36, -10, 47, -57, 90, 98, -40, -79, -52, -57, 62, 4, -54, 62, -45, -17, -106, -91, -84, -50, 107, 100, -91, -46, -2, 14, 90, 79, 23, 76, -58, 107, -122, -114, 98, -79, 64, -123, -108, -6, 36, -43, -53, -116, -5, 126, 41, 47, -18, -70, 39, -118, 86, 111, 89, 75, 109, 99, -104, 71, 121, 87, 79, -88, -13, -92, 84, -75, -6, -52, 1, -72, 52, 10, 62, 68, -118, 76, -8, -30, -45, -49, -62, -53, -104, 12, -116, 39, 120, 42, -94, 0, -99, 32, -110, -10, -126, -113, 119, -33, -16, 20, -110, 57, -64, 53, -113, 64, 104, 88, 63, 36, -46, 44, 60, 43, 119, 37, 108, -37, -67, -38, -7, -31, 67, -9, -53, -24, -50, 121, 69, -71, 43, -66, -74, -51, -27, 95, 57, 31, -119, -99, 126, 103, 47, -10, 26, -125, -4, -46, 71, 69, 85, -118, -65, -18, -68, -117, 90, -26, 28, -36, 90, 111, 56, -68, 97, 51, -34, -103, 85, -65, -42, 116, 7, 30, -84, 12, -18, 21, 72, 43, 119, 26, 104, -24, -92, -98, 120, 99, -93, 30, -65, -18, 46, 70, -30, 48, -114, 124, 12, -4, 65, -115, -49, -124, 49, 25, -43, -9, 93, -6, -78, 24, -53, 71, 78, 81, -37, 32, 29, -11, 18, 21, -35, 72, -14, 26, 121, 18, -69, -97, 27, -56, -73, -88, 38, 85, -86, -38, 25, 91, -25, 99, -48, 5, -100, 51, -29, -126, 80, 68, -46, -89, 36, -20, -44, 95, -7, -118, 32, -65, -112, -62, -80, -14, -124, 47, 90, -115, -94, 53, -116, -49, -3, 70, 84, 89, 57, 0, 71, 73, 41, 20, 98, -115, -2, -118, 6, -58, 36, -104, -60, -37, 94, 15, -85, -37, -38, 73, 75, 97, -105, 97, -33, -115, 110, 81, 92, -59, -95, -56, 58, -126, 109, -85, -66, 55, 8, -101, 109, -126, 42, -95, -46, 90, -96, 69, 75, 81, 81, 14, -48, 65, 60, -98, 95, -34, 50, 15, -87, 78, 110, 125, 52, 117, 71, -121, 46, -72, -78, -66, -57, -109, 36, -68, 76, 122, 92, -30, -5, 90, 60, -39, -96, -127, -104, -61, -117, -30, -106, -117, 57, -100, 43, -113, -29, 127, -87, -117, -36, 50, -3, 58, 45, 5, 56, 37, 10, 13, 3, -93, 68, -19, -23, 94, 87, 55, -124, -36, 49, -120, 48, -56, -28, 75, 38, 118, -94, -17, 109, 103, -45, -82, 69, -103, 127, -12, -16, -47, -31, -2, -86, -21, 93, 24, 54, -64, -90, -74, -105, -91, -70, -14, -93, -2, 56, 11, 105, 111, 48, 61, 121, 90, 48, 13, 9, -89, -11, 66, -127, -30, 11, 44, -24, 7, -4, 121, 101, 21, 114, 75, 94, 72, -82, 35, 93, -2, -27, -36, -103, -113, 55, -27, -120, 68, 104, 20, 3, 63, 36, -86, 82, -42, -58, 42, -17, 47, -111, 22, 37, -93, -61, -22, 77, -80, -16, 15, -57, -54, -37, 71, -83, -99, -66, 4, 43, 27, -128, 57, 14, 68, 14, -19, 80, -5, -9, 8, 65, -100, -85, -128, -33, -81, -79, 50, -91, -107, 89, 31, -90, 35, -7, -56, -21, -37, 60, 40, 119, 86, -79, -65, -87, 46, -8, -69, 23, 42, -123, -6, -45, 19, 28, 74, 117, 45, -24, -54, -127, -51, 12, 94, 92, 79, -95, -96, 49, 36, -12, -88, -57, -38, -5, 112, 26, -48, 9, 16, 40, -24, 83, -115, -55, -86, -12, -38, -44, 16, -90, -114, -90, -25, -109, -76, -83, -50, 42, 122, -116, 17, 17, 81, 77, 111, -54, 100, 67, -7, 121, -32, 49, 56, 59, 98, -49, 58, -85, -29, -29, 13, 58, 70, -63, -54, -96, 82, 19, 76, -60, -99, 28, -101, -28, 67, 111, -40, -62, 45, -102, -123, 33, -78, 47, 16, 13, 45, 78, 15, 10, -24, -125, -108, -2, 95, 7, -103, 13, -32, 37, -35, -48, -126, -126, -97, 30, -40, -51, 24, 48, 96, -112, 101, -127, -116, -47, 1, -5, -41, -18, 26, -110, 56, 21, -111, -91, 73, 57, -113, -21, -102, 75, -76, 55, -52, -71, 74, 104, 76, 14, -41, -24, -17, 103, -86, 46, -39, 114, 5, 104, 95, 27, 108, 52, 44, 108, 35, -48, 75, 13, 68, 42, 106, -41, 58, 56, -30, -21, 103, 122, 36, -13, -76, 79, 12, -107, -9, 7, -4, 105, -71, 72, 70, 83, -116, -42, -54, -79, 88, 43, 79, -112, -4, 36, -124, 19, 113, 4, 69, -42, 102, 31, -19, -48, -29, 29, 31, -22, 115, -10, 44, -20, -54, 2, 89, -29, 75, 59, 33, 93, -117, -13, 47, -109, -61, 11, -49, -98, -107, 80, 5, 57, -12, 34, 114, -81, 127, 68, 54, 30, 78, 91, -121, 8, -93, -62, -43, -89, 1, 70, -23, -16, -98, 60, -12, -109, 4, -11, -109, 114, 84, 110, 84, -119, 64, -83, -14, 119, 34, 109, 63, -55, -122, 62, -23, 96, 61, -72, 35, 4, -89, -36, 20, -72, -62, -17, -31, -119, 8, -17, -82, 55, -7, -30, 17, 83, -98, 28, 5, -120, 81, -37, -103, -81, -96, 26, 76, -103, 74, 37, -18, -125, 120, -71, -2, -22, 2, -74, -88, 88, -1, 118, 76, 50, 14, 58, 9, 19, -12, -119, 39, 38, -120, -5, -36, -117, 110, 28, -121, -25, -23, 87, 42, 58, 83, 76, 37, 100, -23, 32, -33, -118, -103, 97, 96, 70, 10, 36, 65, 23, 5, -70, 11, -60, 93, 9, -13, 26, 71, 80, -43, 82, -48, -63, 50, 44, 47, -119, -123, -105, -52, 34, -71, 49, -17, 112, -71, 56, 106, -75, 119, -85, -127, -42, 6, -124, 4, -111, -104, -1, 124, -41, -85, 21, -6, 101, -98, 109, -119, -58, -122, 86, -16, -75, -35, 127, 79, -7, -128, 22, -83, -23, -100, -26, -50, -111, -16, -85, -22, 86, -38, 43, -10, -75, -44, -3, 109, 58, 14, -18, 23, 106, 73, -105, -14, -100, -66, 124, 67, 29, -15, 105, -11, 60, -4, -46, 86, 41, -126, -122, 34, -34, -43, 27, 93, 14, -67, 49, -89, -24, 22, -71, 124, -31, 83, 117, 32, -104, -95, -35, -57, -83, -49, -127, 30, 85, -97, -100, 120, 62, -127, -37, -112, 89, -34, -9, -71, 10, -37, -17, 115, 102, -96, 99, -27, 110, 107, -78, -3, -121, -91, -42, 75, -72, 49, 6, -122, 6, -25, -29, 51, 0, 118, -90, -41, 101, -34, -16, 73, 28, -13, -116, 118, 73, 122, -5, -21, 48, -82, 98, 77, 41, 102, 26, -98, 122, -125, -76, -6, -94, 120, -64, -85, 0, 22, -22, 73, -62, -34, -94, -39, 36, -40, 20, 90, 121, -1, -29, -72, -16, 32, 27, 48, -19, 14, -110, 32, -55, 50, 18, -57, -109, -15, -13, -69, -79, 39, -87, 0, -128, -114, -53, -77, 104, -89, 102, 47, 4, -54, -126, -120, -122, 21, -91, 80, -106, -3, 70, 94, -23, 62, -92, -69, -31, -111, -92, -99, 42, 47, -6, -81, -50, -128, 86, -127, 100, 113, -3, 29, -39, 9, -116, 110, -92, 125, -64, -35, 114, 125, 94, -106, 7, -55, -21, -7, -58, 95, 78, -122, 44, 42, 25, 79, 35, -30, -11, 127, 115, -100, 106, 45, -84, -74, -47, -118, 23, -99, 0, -108, 46, 12, -109, -122, 29, -78, 66, 84, -69, 85, 22, 48, 27, 101, -117, 1, 14, 106, 35, 125, 86, -119, -5, 64, -44, -72, 5, 127, -65, 49, 89, -14, 22, 119, -120, -47, -128, -102, 122, 73, 93, 36, 37, 107, 92, 119, 37, -44, 96, -10, -70, 53, 94, -113, 121, 66, -89, -9, -64, -20, 6, 58, -127, -26, 84, -31, -23, 38, -90, -6, -60, -127, 47, 39, 96, 58, 4, -44, 68, -31, -96, 83, 14, 127, -60, 64, -74, -40, 42, 117, -65, -117, -63, 69, 93, -74, -28, -94, 56, -12, 107, 84, 56, -6, -9, -14, 55, 123, -17, -64, 121, -56, 48, 87, -117, -73, -45, -73, 48, -70, -6, -76, -45, -15, 79, -77, -47, -88, 112, 51, -47, -99, -95, -74, -11, 72, -29, -109, -77, 70, 30, -96, -97, 53, 115, 104, -80, -67, -3, 109, 88, 8, -106, 23, 27, -49, 77, -17, -82, -86, 19, -43, -125, 53, -23, 79, 88, -75, -49, -46, 100, -102, 104, -108, 28, -18, 121, -4, 57, -45, 38, -102, -18, -102, -46, 51, -109, -91, 37, 86, -128, -74, -11, 22, 79, -72, -27, -9, -72, 41, -34, 53, -31, -53, -123, -33, -58, 8, -13, 4, -66, 32, 7, -125, 15, -93, -93, -46, 22, 14, 43, 125, 120, 75, -123, 3, -92, 96, 68, 36, -32, -114, -7, -49, 117, -28, -3, 99, -37, 67, -72, -53, 33, -77, -94, -55, -33, -17, -77, 17, 11, -57, -56, 90, -41, -110, 75, -25, 65, -10, -90, 12, 63, -19, -51, -122, -54, -71, -127, -91, -51, 72, 116, 84, -98, 8, 24, 40, -85, 57, 1, -39, 18, 18, -26, 99, -15, -96, 103, -22, -78, -12, -14, -45, -61, 83, -121, -40, -24, -83, 79, 64, -48, -44, 48, -3, -11, -82, 115, -93, -127, -13, 17, -96, 126, -39, 37, 4, -84, -19, -66, -9, 81, -77, 19, 91, -53, -3, -62, 33, -47, -123, -41, -105, -81, 65, -93, 57, 23, 20, -33, 10, -104, -122, 29, 60, 9, -1, 54, 93, 34, -19, -75, -100, -120, -32, -47, 67, 98, 62, -127, -96, -84, 33, 32, 79, -4, -24, 49, 71, 124, -11, 60, 78, 48, -8, 60, -110, -123, -126, -78, 80, 46, 25, -30, 14, -94, 91, 103, 27, -106, -110, 71, 70, -55, 116, -25, 43, 5, -88, -98, 69, 104, 124, 64, -91, -119, -44, -107, 47, -67, 73, -8, 114, -106, 113, 75, -12, 27, 33, -84, 50, 97, -128, -5, -33, 11, -33, -23, 83, -29, 90, 99, -124, -70, -89, 8, -125, 60, -55, -99, -63, 65, 109, 33, 45, -118, -41, -58, 43, -65, -47, 72, 75, -2, 123, -54, 94, 99, -65, -48, -2, -72, 107, 50, 107, -68, 103, -88, 106, -62, -56, -51, -123, -105, 101, 81, 118, -2, -49, -5, -63, -49, 71, 80, -107, -24, -11, -34, -16, -25, 107, 122, 111, 66, -86, 71, 51, 82, 101, 18, -62, -63, -38, -110, 45, 3, -30, 18, 99, -123, 83, -78, 25, -52, -19, -90, -97, 84, -15, 96, -97, 119, 69, 15, 52, -38, 38, 71, -84, 47, -31, 29, 93, -67, -123, 75, 105, -2, 76, -19, 65, -8, -39, -5, -115, 14, -116, 24, 45, 25, -113, 96, -101, -47, -7, -85, 99, 110, -31, -112, -75, 111, -75, 70, -108, 94, 20, -53, 10, 16, 67, 4, -93, 68, -99, -120, -12, 119, -122, 120, -37, -35, -2, 115, -113, 63, 47, -111, -55, 90, -118, -60, 36, 19, 6, 77, 120, 62, 3, -53, -3, 78, -68, 42, 113, -28, -119, 4, 76, -99, -71, -19, 99, -76, -33, 38, -33, -20, -85, 124, 125, 16, 61, 81, -125, -2, 50, -24, -87, 93, 66, 91, 49, -61, 57, 74, 43, 85, -29, -105, -79, -10, 124, -26, -89, -45, 84, -59, 24, -40, -110, 111, 101, 24, -91, 91, 82, -9, 72, -79, 49, 75, 5, 105, 17, 19, -105, 117, -101, -114, 25, 72, 102, 114, -21, -72, -17, 59, 97, -62, -45, 8, 37, -65, -19, -13, -35, -124, -70, -44, -26, 113, 88, -105, -64, 94, 36, -42, -17, -63, -42, 117, 30, -58, 6, 90, 28, 84, -58, 46, 54, 98, 89, 46, 66, -91, -29, -111, 8, -61, 7, -80, -14, -1, -15, 111, -115, 59, 117, 83, -127, 113, -82, -23, -23, 18, 18, 107, 51, -78, 126, 41, 126, -118, -70, -22, -41, -2, 28, -46, 16, -48, 40, 93, 97, -48, 29, 83, -38, -35, 5, 37, -97, 64, 27, -60, 79, -8, -113, 71, 103, 36, -124, 113, -70, 59, -49, 80, -97, -113, -18, -88, 3, 110, 41, 13, -11, -4, 121, -50, -9, 47, 105, -10, -15, -86, -23, 87, -52, 57, 30, 113, -111, -99, -121, -101, 105, 63, 107, 126, -40, -92, 28, 5, 0, -52, -41, -90, -56, -34, -127, 85, 121, 64, -128, 41, 28, 75, 43, -28, 48, 38, -31, 27, 81, -71, 69, -59, -97, 113, 120, -105, -107, -60, -22, 85, -66, 118, -68, -11, -99, -128, -54, 72, -20, 110, 53, -93, -16, 53, 108, 9, 99, -83, 14, -39, 99, 113, 97, -97, -10, 119, 61, 13, 106, -52, 124, 123, -57, 9, -19, -54, 74, -61, -21, -113, -44, 13, 82, -1, 32, 93, 124, 60, -94, -115, 123, 77, -119, 81, 6, -32, 70, 114, 29, 53, 76, 109, 72, 36, -9, -48, 113, 9, 66, 2, -36, 71, 88, 0, -74, 14, -55, 95, 115, 42, 76, -118, 16, 32, 56, -11, 110, 19, 44, 45, 79, -53, 119, -68, -86, -97, -84, -114, -108, -45, 11, -99, 126, 83, -1, 37, 118, 47, 123, -128, 33, -13, -7, -75, -101, -8, 108, 39, 123, -118, 114, 46, -8, 74, -55, 51, 116, 70, 73, 112, 52, -95, -41, -99, -101, -53, -106, 96, -28, -70, 81, 100, 72, 58, 51, -73, 53, -94, -13, -116, 94, -125, 99, 7, 98, -41, -78, 3, -71, -98, 112, 12, -122, 64, 40, 19, 120, 56, 76, 22, -4, 80, -19, -10, 29, 118, 49, 59, -50, 67, 52, -72, 7, 76, -92, 77, 115, 76, -22, -34, 81, -115, -29, -113, 84, 96, -57, 9, 18, 123, -127, 86, -40, 14, -53, 91, -82, 19, -122, 15, 43, 24, -72, -13, -10, -16, -26, 21, 81, -13, -118, 76, 47, 123, -79, -44, 76, -67, 106, 29, -96, -97, -62, 29, -13, 49, -21, 104, 78, -77, -94, 14, -55, -69, -105, 81, 85, 8, 114, -27, 19, 110, -76, 72, -47, -105, -103, 47, 12, -59, -92, 72, -9, -112, 58, 6, 118, -106, -85, -37, -123, 66, -47, 15, -127, 68, 80, -115, 109, 11, -34, -78, -116, -44, -19, -50, 46, -56, 18, -25, -36, 7, -62, -25, 101, -79, 5, 118, 10, -46, 84, -87, 3, 10, 42, -32, -51, -51, -55, 108, -95, -20, 124, -58, -45, 43, -124, -68, -33, -5, -100, -124, -29, 2, -3, 124, -62, 11, -18, -70, -97, -111, -80, 72, -1, 0, 93, -6, 15, 91, -47, -80, -54, -34, 92, 116, 48, -108, -87, 10, -43, 127, 48, -21, -113, 30, 70, -3, 20, -101, 120, 73, -115, 11, 125, 113, -5, 26, -69, 109, -53, 50, -58, -41, -5, 76, 49, -114, 44, -99, -108, -16, 109, 92, 109, -33, 76, 22, 96, 9, -66, 30, 90, 19, 118, -66, 126, -39, 16, -10, 103, 91, 31, 127, -7, -127, -96, 118, -113, -103, 127, -70, 44, -74, -112, -42, 94, 38, -27, -108, -104, -114, 79, -106, -41, 7, 35, 124, -86, 78, -62, -117, 0, 113, -10, -71, -5, 95, -25, -18, -120, 55, 125, 28, -104, 60, -54, -89, -88, 55, 121, 54, 16, 64, -64, -11, -80, -33, -58, -58, -60, 100, -119, -77, -50, 10, -23, 41, 0, -111, 9, 19, -101, -93, 30, 1, -39, 65, 67, 93, 88, -3, -83, -81, -79, -102, 7, -62, -37, 122, 25, -7, -34, -66, 88, -47, 93, -58, -41, 98, 72, 118, 117, 115, -31, -115, -121, -64, -106, -70, 17, -65, -80, -29, -27, -54, 23, -110, 89, 39, 77, 73, -48, 40, -123, -81, 104, 111, 56, -99, 98, -107, 93, 68, -68, 44, -25, 56, -95, 4, 79, -53, -3, -106, -42, 42, 116, 56, -81, 125, 118, -40, 41, -68, 43, -30, 111, 43, 43, 120, 120, -85, 117, -48, -53, 93, -97, 103, -49, 92, -74, 68, -27, -68, 18, -75, -7, 109, -27, -35, 41, 45, 7, -21, -78, 30, -41, -16, -14, 115, 32, 112, -30, 58, 17, -3, 111, 47, 124, -9, -24, 116, -14, -120, -103, -28, -86, 25, 29, 127, -19, 57, -65, -127, 101, -67, -110, -125, 83, 52, 127, 103, -80, 76, -101, -122, 32, 32, -86, -109, 81, -72, 4, -46, 104, 76, 0, -48, 45, -43, 99, -118, -67, 110, -18, 59, 51, 47, -63, -108, -65, -58, 121, -123, 58, -7, 99, -112, -49, 55, 81, -77, -27, 106, -52, 88, 94, -84, 109, -9, 58, -91, -127, -22, 12, -6, 84, 11, -69, 55, -77, -113, 95, 110, 5, -119, 55, -4, 28, 117, 101, 3, -59, 99, 112, -53, -33, 22, 74, 41, -97, 35, -30, 122, -118, -48, 123, 18, 122, -109, -8, 94, -117, -109, -51, -32, 110, -118, 102, 13, -39, 59, 3, 30, -51, -88, -111, -118, 34, -86, 51, 108, -74, -97, -67, -121, 60, 81, -71, -12, -121, -30, 18, -105, 49, -128, -4, 25, -83, -42, 26, -68, 108, -71, -2, -62, 55, -90, 2, 15, -105, -112, -86, 77, -112, 48, 98, -33, -4, 101, 12, -52, 66, -6, 108, 102, -53, 36, 4, 40, 36, 111, -25, -10, 42, 68, 26, 7, 91, 56, -104, -6, -29, 47, -114, -107, 100, 23, 46, -22, -71, 0, -75, -67, -22, 7, -10, -7, -63, 12, 100, -38, 30, -88, 5, 25, 30, 7, 115, 32, -24, 25, 90, 121, 19, -26, -112, -16, 62, -112, 98, -101, -121, 123, 85, -100, -27, -115, -95, -128, 35, -116, 50, 63, 66, -39, 15, 33, -7, -2, 84, 94, -23, 23, 71, -80, -27, 93, 6, -10, -2, -7, 27, 51, -114, 96, 79, -30, 70, -81, -25, 71, -119, 45, -78, -42, -73, -100, 35, 54, -19, -54, 33, -119, -109, -127, -51, 115, -20, 38, 94, 32, -120, -90, 73, -17, 11, -85, 121, 14, -93, -55, 68, 126, -90, -99, 47, 20, -93, -39, -73, 70, -21, -18, -90, 18, 43, 87, -60, -56, -5, 40, -16, 103, 8, -13, -6, 116, 69, -45, 127, -52, 6, 87, 113, 4, 43, 125, 63, -101, -36, -99, -6, 16, 0, 59, 94, 106, 41, 121, 117, 73, 70, 24, 115, -99, 65, 89, 25, 49, -28, 65, 12, 33, -125, 13, 85, -113, -48, 82, 46, -13, 51, -88, -85, -40, -40, -3, -121, -65, 75, 39, -58, 42, -127, -16, -13, -24, 21, 81, 78, 60, 83, -64, -35, 96, -71, -119, 27, 126, -15, -102, -55, -16, 95, 51, -40, -49, -114, -2, 18, -11, -104, 115, -123, 58, -53, 73, -30, 4, 94, 5, 65, -77, 104, 103, 10, -103, 35, -28, 90, 47, 19, 7, -70, -98, -63, -107, 27, -79, 80, -87, 23, -125, -19, -80, -57, -114, -101, 97, -41, 83, 12, -33, 27, 55, 45, -115, 65, -78, -108, -34, -29, 17, -28, -36, -55, 54, -36, -6, -57, 16, 65, 36, 32, 123, 15, 104, -115, 111, 78, 101, -95, -45, 126, -63, 56, -4, -20, 1, 25, 53, 38, 89, 48, 107, -44, 44, -93, 55, 124, 1, -10, -52, 116, 41, -78, -115, -60, 10, -96, 19, 12, 93, -40, -115, -77, -20, 105, 46, 108, 50, -124, 124, 81, 114, 127, -11, 52, 118, -112, -32, -39, 83, -107, -29, 83, -25, 99, -13, 47, 94, 68, 21, -25, 86, 78, -93, 91, -47, -106, -80, 119, -6, -51, 104, -12, 18, -71, 5, -23, -70, 12, -88, -115, 101, -127, -33, 125, -112, -13, 125, -1, -120, -105, 66, -92, -57, -71, -26, -109, 95, 72, 123, 12, 15, 58, 51, -103, 45, 122, 87, 51, -116, 1, -59, 58, -6, -51, 80, 36, -65, 15, -2, 122, 107, 47, 59, 71, -67, 28, 74, 15, -93, 11, -4, 13, 43, 60, 2, 52, -90, 100, -29, 26, -36, -76, -48, 89, -90, -86, -20, -69, 52, -3, 9, -53, -103, 107, -28, 80, 61, 74, 20, 23, -70, -20, -28, -8, -119, 40, -47, -79, -112, -32, -53, -73, -31, 72, -113, 23, 81, -53, -62, 62, 42, 1, -35, 21, 83, 88, -87, -49, 55, 40, 102, 120, 14, -50, 3, -119, -121, -120, 16, 82, -66, -8, -27, 99, 28, 7, -20, 76, 53, 120, 19, 67, -4, 6, 5, -19, 27, 96, -33, 54, 108, 50, -62, -113, 94, -41, 115, 119, -82, 62, 32, 118, 38, -8, 88, -120, 50, -65, 11, 58, -64, -73, -31, 36, -67, 77, -121, -93, -25, -28, 66, -71, -90, -51, -118, -36, 16, 66, -121, 54, 97, -119, 124, -2, -124, 16, 91, 2, 104, -22, 32, -16, -51, -71, -89, 123, 61, -112, 107, 107, -78, 18, -76, 65, 123, 121, -44, -91, -43, -107, -94, 102, 91, 71, -46, -63, 87, -84, -20, 112, -43, -37, -41, -67, -4, -104, 121, 4, -47, 95, -6, -4, 66, 114, 84, -68, 77, -94, -68, -37, 47, -112, -86, 102, -24, -51, -127, -34, -42, -57, 80, 31, 41, 62, 27, -22, 95, -81, -78, 9, -94, -26, -14, -13, -112, -7, -81, -33, -59, 16, 112, -18, -101, -67, 11, -33, -66, -83, -120, -60, -4, 79, -65, 37, -29, 11, -74, -59, -121, 124, -64, -68, 105, -96, -16, -70, -108, 79, -16, -24, 62, 16, -115, -83, 14, -20, 92, -37, 91, 13, 14, 20, -113, 89, -6, -90, -26, -89, -48, 79, -11, 61, 27, 81, -58, -106, -88, 114, 48, -82, -68, 74, -24, -112, 20, 104, 66, 51, 120, -119, 10, -42, 1, -93, -22, -94, 54, -65, 45, 11, -5, -93, 104, -16, 49, -125, 76, -80, 80, -109, -80, 40, 87, -64, 127, -108, 31, 56, 54, 24, -64, -72, -86, 81, -51, 99, 97, 101, 47, -98, 103, -46, -52, -6, 54, -99, -52, -86, -13, 33, -34, -82, 22, 78, 56, -58, 70, -40, -19, -116, -118, 82, 14, 16, 91, 1, 5, 22, 0, -107, -109, 54, 58, -78, 72, 23, 87, 29, -119, 122, -102, 111, 119, 90, -106, -125, -40, -80, 95, 9, -32, 80, 52, -79, 46, 109, 101, -13, 65, 87, 54, 53, 98, 100, 75, -57, -39, -5, -92, 30, 73, -63, -69, 127, 30, 104, -45, 11, 106, -45, 52, -34, 27, -31, -103, -56, 53, 92, -20, -11, 37, 15, 25, 116, 78, -1, 88, 76, -25, -108, -93, 36, 40, 35, -101, -6, 83, 92, 56, -119, 0, 19, 9, -33, -10, 63, -56, -79, 1, 60, -64, 105, -48, 113, -37, 0, 76, -89, 24, 112, 25, -125, -76, 49, 120, -52, -50, 20, 51, 21, 98, -24, 73, 119, -73, 20, -76, -41, -109, 115, 103, 34, -60, 5, 84, 36, -21, 6, -109, -82, -91, -78, -27, 123, -25, 94, -116, -67, 121, -72, 100, 122, -94, 83, -67, 7, 67, 97, -20, 42, 124, -8, 13, 69, -77, -119, -84, 41, 53, 61, 5, -101, -21, 43, -62, -93, 66, -108, -63, -110, 77, -12, 0, -27, -54, 86, 18, 112, -41, 95, 72, 38, 86, 52, -75, -97, 3, 54, 121, 32, -43, -70, -124, 90, 30, 80, 91, -12, 112, 74, 22, 122, -89, 61, -57, 31, -86, -123, -110, 79, 15, 92, -110, -96, -82, 15, -122, -67, -62, -54, -36, 25, 66, 105, 13, 91, -21, 69, 11, -69, -11, 35, 10, 72, -13, 91, -51, -37, 48, 113, -4, -49, -39, -44, -114, 92, 50, -74, -73, 21, -72, 6, 73, 117, -121, -40, -35, -42, -70, -51, 91, -106, -121, -42, -29, -114, -93, -9, 51, -95, -22, -117, 81, -35, -15, 118, -41, -39, 93, 117, -17, -80, 115, 66, -68, 100, 50, -25, -81, 119, -50, -93, 3, -53, 12, 113, -37, 16, -91, 59, 31, -32, 54, 57, -3, 2, -73, -16, -118, 73, -118, -14, 66, 2, -75, -56, 49, -70, -78, -23, 8, 31, 57, 53, 30, 28, 80, 47, -8, -31, -66, -26, 102, -52, 24, 4, -49, -52, -102, -111, -77, -116, -81, 112, 0, -88, -63, 103, -47, -22, 55, -70, -7, 117, 23, 21, 14, -47, 51, 4, -52, -11, -58, 5, 33, 59, -51, 55, 16, 2, -15, 75, -17, -85, -112, -125, 60, -97, 79, -37, 90, -79, 101, 73, -28, -51, 120, -12, 49, 54, -60, -29, -39, 65, -128, 19, -97, -3, -71, -39, -99, -21, -41, -3, 77, 108, 53, 53, -86, 84, -44, 55, -26, 33, -51, -54, -77, 24, -59, 34, -125, -68, -86, -83, 10, 73, -64, 111, 106, 45, 105, -126, -18, -10, -103, 87, -103, -106, -76, -104, -31, 63, 94, -98, 28, 36, 54, 85, -40, 125, 51, -78, 8, 74, 79, -16, 37, -6, 66, 76, -51, -31, -99, -11, 110, 82, 53, -55, -122, -100, -107, -52, 96, -16, 113, -74, -87, 96, 38, 123, -9, 28, 28, 6, 38, -99, -80, 72, -81, 18, 47, 116, -123, 92, 90, -15, 100, 10, 36, 59, 19, -97, 50, -106, 31, 50, 12, 79, 15, 57, 41, -79, 37, -74, -10, 13, -71, -27, -74, -82, 117, -53, -64, 59, -107, -67, -122, -36, -77, -72, 44, 13, 125, -23, 38, 14, 46, 51, 86, -33, -127, 27, 96, -123, 57, -43, -112, -53, 42, -102, 93, 116, 54, -69, -70, -85, -8, -88, 10, -43, 51, 1, 11, -112, -83, 30, -79, 32, 76, 119, -41, -41, -85, -95, 120, -119, 123, -115, -68, -21, 39, 45, 65, -58, -116, 100, 44, -1, 97, 102, -34, 54, -33, -29, 66, -48, -76, -16, -90, -26, 41, -68, 119, 14, -63, -53, 77, -23, -120, 63, -28, -67, 79, -109, 1, 123, -34, 50, 52, 21, 23, 122, -126, 33, -40, -79, -5, -96, 6, -95, 30, -127, -36, 82, -26, 41, 32, -81, -11, 37, 69, 95, 38, 120, 5, -81, 99, -120, 45, 123, 90, -54, 41, -16, -6, -22, 122, 23, -77, -27, -68, -82, 99, 17, -10, 32, -84, 73, -10, 114, 90, 112, -121, -65, -14, 103, 65, 29, -101, -83, 35, -128, 68, -57, 107, 111, -79, 51, -104, -99, 62, -27, -46, 7, -25, -49, -65, 110, 106, 91, 80, -119, 105, -86, 84, 113, -99, -9, 71, -114, -34, 125, 101, 65, 37, 26, -84, -25, 89, -76, -27, 43, 33, 38, -114, -106, -42, -29, 110, 77, 63, -97, 121, -101, -79, 49, -72, -74, 82, 47, 24, -23, -58, -86, 114, -46, -65, 44, 89, -77, 96, -40, 49, -108, 112, 104, 113, -78, 67, -98, -25, 67, -105, -95, 29, 65, -68, -42, -24, -81, -60, -101, 71, 50, 100, 90, 63, 39, -100, -118, 19, 9, -62, -128, -6, -51, -84, -76, 115, 53, -39, -63, -17, 86, 100, 85, 86, -69, -64, -74, -99, 120, -2, -107, 10, 115, 39, -51, 50, 124, -67, -126, -106, 62, -39, -71, 48, -92, -50, 56, -94, 14, -45, 103, 18, 102, -16, -123, -78, -58, -109, 108, -69, -110, 2, 82, -72, -100, 120, -73, 79, -3, -2, 12, 114, -85, 72, 52, -98, -82, -87, 95, 28, -37, -100, -27, 91, -57, -118, -110, -111, -125, -14, -33, -96, 79, -89, 21, -13, 99, 115, -7, 108, 29, -112, -109, 14, 104, 37, -37, -51, 60, 68, -55, -62, -127, -118, 46, 16, -57, 12, 68, -66, 7, -114, -46, 119, -49, -40, 69, 88, 111, -116, 66, 100, -43, 59, -126, -125, 96, -68, 102, 117, -105, 88, 103, -45, -120, -109, -7, 38, -118, 81, 56, -102, -64, -34, 122, 9, -39, -8, 108, -109, -114, 67, 69, -51, 116, 42, -25, 101, 21, 24, -116, 63, -112, -65, -5, 47, 96, -71, -78, 88, -79, 123, 55, 94, -108, -122, 26, 20, -11, 69, 49, 67, 46, -122, -110, 104, -107, -89, 60, -92, 3, -112, -114, 26, -65, -20, 75, 20, -40, -75, -57, -57, -114, -53, -12, 16, 116, 44, -50, 99, 66, 1, 8, -125, -104, -20, -81, 95, 106, 61, -104, -37, -95, 114, -63, -109, -46, -18, -112, 33, 125, -12, 113, -48, -12, -81, 59, 22, -98, -13, -34, 117, -117, -50, 22, 20, -91, -70, -52, 22, -55, -107, -71, 66, 82, -59, -85, -40, 95, 76, 119, 70, 24, -115, 70, -57, -84, -103, 24, 95, -121, -36, 5, 70, -119, -63, 59, -61, -13, -47, -43, 17, -128, 96, -27, 59, -44, -99, 12, -43, -51, 91, 86, -6, -93, 116, 75, 77, 95, 87, 92, 40, 117, 58, 81, 68, -91, -57, 54, -18, -72, 76, 109, 108, 42, -51, 80, 40, -74, -24, -101, -6, 30, 25, -37, -71, -44, 60, 20, 19, -78, -59, 94, -128, 24, -32, -9, 118, 27, -58, 91, 91, 9, -37, 113, -128, -107, 20, -81, 98, -100, -63, -113, 113, -53, 35, -12, 16, 87, 68, -7, -81, -75, -85, -25, 63, -95, 47, -68, -29, -68, -113, 64, 70, -67, 51, 17, -35, -6, 77, 19, -40, -12, -6, -32, 72, -1, -122, 15, 110, 77, -42, 57, -2, -99, 99, -35, -23, -93, 26, 85, -49, 62, -117, -69, 107, -66, -103, 65, 110, -19, -53, 10, 97, 39, -91, 94, 47, -116, 76, 54, 115, 31, -122, -77, 30, 38, 22, -39, -33, -118, 51, 16, -19, -126, -3, -124, 120, 76, 124, -92, 47, 5, 102, -20, -124, -33, 21, -61, -30, -7, 47, 83, 53, 61, -48, 10, -67, 122, 0, -118, 14, -85, 2, -65, -47, 46, 113, 17, -89, -53, -65, 45, 74, 123, 92, -80, -116, -101, 33, 89, 68, 105, 78, 11, 93, -82, 102, -58, -19, -75, 13, 73, 6, 8, 102, -23, 67, -78, -48, -85, 63, 124, 78, 56, 41, 69, -101, 68, -98, -41, 17, 54, -18, -99, 121, 80, -7, -51, -116, 8, -91, -73, -33, -35, -10, -46, 81, 61, -75, -103, -9, 19, 1, -95, -122, 35, 60, -98, 13, -45, -86, -95, -109, 59, 9, 107, -66, -88, 14, 49, 106, 101, 48, 104, -118, 8, -68, -9, -91, -79, -107, -128, -40, -93, 66, 115, -4, -86, 13, -114, -103, -9, -108, 50, 11, 21, 52, -46, 45, 27, 12, 125, 25, 36, 123, -12, 63, 65, 10, -6, 108, -31, 71, -25, 12, 10, -64, -56, 110, 10, -14, 57, -100, -83, 26, 16, 115, -14, -23, -12, 28, -100, -103, -88, 106, 95, -107, -126, 103, -44, 110, -51, 69, 98, -113, -83, 33, -27, 81, 125, 23, -33, -13, -95, -55, -54, 60, -111, -87, 127, -17, -33, 114, -26, -25, -59, 14, 109, 72, -74, -31, 67, -85, 125, -75, 15, -24, -56, -109, -45, 104, -71, -92, 85, 62, 12, -105, 102, 70, -103, 93, 25, 125, 44, -62, -115, 118, 11, 60, 59, -66, -85, 64, -123, 26, 0, -36, -59, -117, 123, 59, 124, 115, -71, 119, -112, -94, 72, -101, -31, -122, -8, -20, 47, 106, 115, -34, 53, -61, 69, -95, 104, -4, 101, 24, 38, 116, -73, -112, -120, -104, -62, -10, 78, -77, -42, 87, 123, -88, -26, 62, -30, 54, 25, -86, -24, -95, -92, 46, -53, -18, -34, -9, 83, 69, -97, -104, -70, -77, 44, 34, 118, -107, -67, -37, -101, -78, -18, -81, 88, 115, 12, -61, -13, -12, -89, -116, -73, 52, -97, -114, 66, 25, -11, -71, -12, -87, -115, 27, -90, -54, -123, 24, 49, -15, -37, 66, -36, 71, 1, -57, 13, 6, -92, -23, -92, 98, -35, -115, 77, 40, 39, 81, -36, -109, 108, 110, -7, -2, -4, -27, 11, 48, -108, -64, 126, -35, -67, -87, 4, -121, 98, 116, -126, 105, 18, 106, -8, 79, 44, 88, -72, 30, 9, 80, 46, -23, -74, -88, -126, 50, 23, 1, -77, -101, -79, -91, 61, -76, 66, 84, -43, -18, 6, 63, 64, 34, 117, 79, 96, -11, 24, -82, -127, -2, -106, -42, 44, -24, 56, 126, -114, 44, 78, -53, 121, -55, 10, 121, -105, 84, 25, -75, 72, -33, -122, 41, -68, 12, -35, -99, 122, 61, -24, 3, 64, -54, -75, 59, -94, -33, 59, 118, -30, -90, 55, -28, -110, -112, -62, 103, 108, -104, 89, -45, 122, 70, 54, 79, 103, -25, -20, -101, -71, -67, 91, -5, -48, -11, 104, -112, -111, 15, 38, 38, 60, -26, 89, -78, -109, 48, 80, 55, -21, -35, -57, -50, -88, 19, 70, -56, 24, 70, 29, -69, -85, -25, 100, -22, 122, 94, -6, 127, 50, -18, 64, -75, -48, -77, 105, 8, -38, 88, -84, -51, 4, -35, 85, 84, 73, 96, 3, -55, 45, -119, 111, -58, 6, -24, -53, -49, -39, -83, 105, -109, -3, -44, 79, 86, -68, 62, -110, -22, 37, -25, -101, 11, 5, 67, 25, 40, -52, -7, 10, -73, 126, 61, -103, 67, -125, -43, 109, -53, -38, 8, -59, -4, -20, -65, 11, 16, -102, 70, 43, 83, 56, 117, 31, 127, -103, -80, 121, 28, -63, 65, 0, 75, 80, -31, -98, -31, 112, 108, 90, -30, -51, -72, 15, -35, -108, 71, 79, 19, 18, -85, -42, -7, 1, 108, -16, 7, -63, 13, 67, -69, 12, 68, 112, -56, 68, -125, 78, 125, -21, -31, 45, 103, 114, -84, 74, 40, -111, -63, 0, 39, -46, -41, 117, 90, 43, 120, -17, -75, 68, 113, 97, -42, 75, -77, -45, -114, 65, -6, 110, 28, -55, 21, -75, -113, -40, 38, 35, -67, -3, -14, 50, -125, 79, -55, 65, 110, -29, 25, -9, -8, 109, 106, 105, 119, -103, 13, -35, 16, 56, -29, -57, 119, -73, 103, 123, -65, -118, -126, 12, -42, -50, -126, -122, -28, 54, 91, -109, -32, 34, -50, -40, 19, 3, -87, -44, -7, 119, -16, 48, 98, 33, 33, 1, -68, 101, 87, -39, 83, -122, -78, 8, 66, 54, 54, 99, -92, 89, -18, 113, -3, -58, -61, 33, -70, -128, 99, 27, 5, 39, -65, 53, 71, 43, 21, -4, 30, -109, 37, 84, -49, 39, 36, -99, -92, 73, 19, -13, 34, 71, 119, -66, 92, -89, -111, -68, -68, -7, 55, 58, 124, -6, -20, 41, 38, 49, -74, -90, -1, -127, 5, 89, -60, 38, 44, -17, -117, -38, 15, -112, -11, 106, 39, 14, -108, -86, -106, 75, -23, 13, 109, 76, 66, 120, -89, -40, 105, 9, 88, -18, 13, 119, -83, -70, -39, 38, -97, 41, 36, 48, -24, 104, -124, -34, -69, -53, -4, -24, 37, 45, -51, 7, 38, 48, -25, -87, 71, 73, 62, 105, -37, 27, -6, 20, 15, -7, -22, 109, -35, -11, 51, 22, -83, -92, 61, -75, 103, 53, 96, -61, 50, -84, -85, -101, -74, -92, 22, 2, -85, -23, 93, 90, -102, 8, 32, 115, -105, 124, 7, 3, -105, 123, -84, 30, 96, 50, 28, -27, -94, 75, 118, -31, -68, 53, 55, -109, -17, -124, 46, 117, 95, -95, 41, 20, 10, -58, 39, 110, -22, 21, -96, 79, 89, -19, 84, 118, -28, 63, -12, 16, 14, -84, -7, -107, 101, 117, -35, 32, -52, -38, -102, 113, 98, -22, 120, 19, -7, -116, 5, 86, -116, 116, -90, -128, -86, 9, 83, -72, -120, -119, 19, -72, 24, 58, 14, -109, -15, -122, 13, -46, 22, -60, 67, 81, -115, 106, -53, 92, -9, 120, 60, -73, -3, -63, -70, 122, 33, 61, -115, -127, 34, 60, -5, -105, -5, 67, 37, 0, -19, -5, -78, -105, 81, 17, -32, -33, -48, 60, -16, -15, -81, 90, 0, -74, 127, 68, -103, -95, -4, 23, 86, 93, -103, 33, -39, -82, -41, -98, 45, 88, -40, -12, 5, -123, -34, 23, 5, 20, 8, -53, 0, 10, -38, 65, 64, -118, -8, -37, -107, 9, 34, -127, 77, 51, -72, 17, 1, -7, 76, -63, -62, 65, 69, -49, 116, -112, 92, -16, 64, -123, -96, -103, 55, -41, 25, 56, -3, -42, 126, -104, -13, -7, 88, 112, -126, 102, -62, 96, 47, 125, 50, -124, -28, -56, -124, -77, 0, 55, -116, -86, 110, 100, -72, -114, 87, -59, 109, 31, -94, -40, -94, 54, -82, -110, 110, -61, 54, 28, -75, 77, 57, 16, -100, 24, -85, 33, -8, -98, -85, -66, -29, -128, -45, -77, 119, 15, 107, 20, -2, -28, -81, -108, 122, -13, -16, -12, -42, -37, 26, -53, 91, -120, 29, -22, 15, -70, -39, -88, -77, -50, 52, 50, 92, 92, -65, 67, 99, 119, 32, -118, -44, 5, 24, 108, -89, 95, 108, 87, 76, 112, 87, 50, -102, -108, -126, 51, -27, 114, 82, 17, 63, 44, 61, 13, -123, 15, 60, 3, -54, 49, 35, -60, -32, 13, 43, 11, -3, 12, 13, -5, 96, 102, 88, -81, -51, 117, 20, 7, -69, 102, 15, -119, 116, 109, -57, 17, 52, 12, -73, 100, -65, 100, -18, 40, 98, -48, -80, 89, 47, 93, -26, -52, -121, 44, 105, -94, -76, 49, -36, 113, -26, 78, -13, -64, -40, -40, -20, 84, -122, -56, 9, -116, 73, 29, -34, 27, 116, 47, 108, -51, -108, -33, -24, -68, -16, -29, -12, 45, 31, -68, 35, -31, 118, 41, 45, -101, -42, -91, -74, 38, -116, 6, -47, -51, -95, -85, 100, 7, -10, 79, 108, -48, 88, -114, 57, 59, 89, -43, 80, -98, 6, 78, 88, -122, -35, 14, 89, -75, 116, 104, 88, 124, -105, -82, 80, -45, -1, -44, -39, -43, -74, 86, -108, 115, -64, -85, -5, -100, 22, -121, 92, 62, -101, -98, 6, 34, -66, 90, 51, 88, -88, -85, 6, -67, -112, -19, 19, -24, -70, -24, 65, 81, 43, 31, -40, -27, -79, -68, -103, -17, -39, -92, 122, -115, 81, 98, 103, -15, -72, -112, 0, -24, 44, 74, 37, -53, 19, 121, -49, -79, 72, -122, 46, -57, -43, 98, -117, -73, 117, -95, -104, 48, -76, -100, 111, 18, 29, -82, -97, 17, 99, 53, 27, -13, 125, -76, -50, 110, -48, -51, 41, -115, -97, -38, -35, -124, -128, -12, 60, -95, 92, -35, -50, 14, 65, 72, -7, 110, 6, 104, 115, -39, -19, 16, 114, -73, 106, -77, -34, 27, 108, -101, -22, -11, 97, -26, -35, -9, -62, 26, 122, -28, 111, -114, -46, 111, 84, 121, -125, -68, -41, 0, -51, 117, -82, 39, 119, 118, 59, -50, -31, 72, -127, -22, -122, -115, -106, 11, 115, 44, 92, -83, 60, 63, -60, 91, -41, -91, -20, 56, 56, -71, -16, -54, -54, 101, -34, -70, 75, -29, 89, -11, -46, 77, 120, -110, -122, -88, 125, -25, -123, 69, 33, 124, -55, -5, 29, -123, -122, -84, -20, -87, -82, -128, 111, -94, -61, -88, -41, 123, -113, -47, 5, 67, -95, 24, -47, 30, 88, 96, 121, -109, 0, -39, -118, 106, -120, 118, -128, -77, 18, 62, -87, 103, 16, -87, -70, -103, 73, 41, -116, 30, -61, -23, 123, 44, 58, 40, 27, 50, -31, 104, -50, -116, -126, -74, -107, 55, 52, 90, 37, 69, 16, -61, -121, 93, 86, 53, 103, 54, 32, -124, -21, -19, 49, -113, -61, 71, -89, 2, -55, 114, -57, 10, -104, 69, 6, 2, -41, -106, -89, -50, 35, -45, 55, 14, 7, -117, 105, 71, 3, -50, -57, 28, -120, 90, -55, 35, 82, 20, 89, -48, 84, -16, 85, 30, -18, 127, 54, -18, 83, -63, -95, 97, -60, 27, 2, -59, -52, 7, -83, -2, -33, -103, -42, 29, -34, -10, 97, -81, 124, -39, 13, 39, -27, -82, 26, -66, 65, -1, -96, 86, -105, -45, -64, 55, 33, 64, -15, -123, 6, 105, -10, -7, 59, -55, 82, -99, -63, 19, -11, 28, 51, -72, -38, -84, 119, 0, 90, 93, 60, 39, 70, 11, -58, -10, -79, 14, -38, -14, -126, 113, 33, 35, 81, -48, 117, -56, -81, -32, -11, -66, 84, 99, 85, 14, 86, -107, -34, 57, -100, -89, -92, 5, -36, -26, 96, -14, -124, 11, -95, -37, -62, -23, -68, 73, 41, 20, 126, 101, -21, -44, 63, 12, 61, -48, -10, 20, -34, -24, -102, -89, 41, -68, -57, -59, -2, -29, 97, 84, -89, -9, -58, -121, 85, 85, 82, 2, -5, 29, 34, 90, -74, -2, 112, 42, 74, 69, 39, 24, -15, -124, 18, -97, 48, 68, 75, -76, -74, -94, 0, 1, 66, 34, -44, -89, 75, -114, 18, -105, -14, 92, -28, -99, -24, -20, -65, 56, 3, 104, 52, -58, -4, 17, -112, 127, 61, -16, -41, 104, 18, -127, 6, 67, 71, 63, 4, -119, -19, 69, -93, 1, 8, -16, -32, 77, 110, 63, 8, -12, -89, -35, 28, 12, 79, 45, 81, -69, -106, -120, 38, -118, -25, 82, 100, -103, -128, 54, 76, -115, -9, 42, -50, -70, 114, -105, -4, 28, 116, 50, 123, 126, 55, 105, -79, -105, -64, -9, 76, 5, -35, 46, -2, 119, -50, -13, -53, 101, -17, 102, 55, -120, 87, -1, -116, -70, 26, 11, -74, 17, -86, -57, -54, 9, -8, -95, 57, 31, -77, -23, 73, -28, 31, 75, 10, 50, -54, -64, -81, 104, -2, 56, 14, 95, 37, -1, 125, -27, -13, 3, -11, 50, -71, 125, 8, -93, 66, 102, -83, -11, 103, -33, 67, -12, 34, -113, -101, -108, 98, 123, -80, 9, 116, 29, 4, -33, 19, -40, 90, -53, -125, 123, 2, 111, 69, 70, 83, -13, 49, 64, 68, -114, -80, -51, -98, 73, 52, -4, 103, 56, -16, -124, -64, -39, 35, -5, -62, 126, -12, 53, -128, 118, 57, -41, -18, 4, 49, 120, 92, -6, -71, -102, 10, 88, 34, 99, 101, -110, -40, -18, -26, -124, 58, -108, -85, -106, 78, -42, 61, -63, 102, -128, -93, -97, 77, -123, 105, -95, 103, 115, 74, 87, 67, -19, -102, -123, 64, 21, -31, 126, -18, -42, -80, 60, 109, 59, -50, -90, -104, 69, 45, -123, -122, -24, -104, 34, -89, 46, -90, -86, 2, 67, 4, -77, 111, 10, -115, -70, 116, 101, 114, 19, 114, 104, -26, -14, 40, -26, 25, 27, 3, -29, -21, 110, -122, -53, 21, -85, 32, 82, -68, -112, 87, 110, 33, -52, -6, -2, 107, 54, -74, -93, 110, -39, -17, -21, 55, 116, -1, 28, 50, 113, -49 );
    signal scenario_output : scenario_type :=( -78, 2, 127, -55, -128, 127, 127, -79, -128, 54, 127, 6, -98, 117, -90, -24, -128, 127, 127, -78, 31, 1, 34, -128, -12, 29, 119, 127, -114, -128, -128, -8, 127, 29, -128, -7, 127, 60, -128, 54, -1, 44, 86, 101, -73, -128, 2, 15, -7, -123, 122, -74, -128, 5, 127, -52, -128, 22, 127, 127, -47, -68, 6, -38, 127, 85, 127, -26, -63, 36, 127, -128, -128, 42, 65, 127, -70, -6, -75, -5, 68, 27, -95, 21, -36, 127, -10, 47, -128, 127, -54, 69, 28, 93, -81, -128, -12, 0, -6, 88, 127, -33, -121, 2, -8, 127, -39, 73, -128, 60, 81, 127, -128, 66, -50, -128, 119, 127, -96, 13, 127, -28, -128, -11, -92, 55, 127, 23, -128, -128, 127, -78, 127, 24, -123, -123, 127, 127, -21, -128, 76, 68, 50, -128, -16, 127, -57, -128, 116, 43, 31, 117, -68, -68, -42, -123, 127, -116, 80, -102, 0, -128, 127, 127, -32, -128, 127, 16, 57, 3, 28, -69, -97, 71, 8, 7, -44, -100, -18, 127, -85, -128, 27, 127, -42, 23, 49, 0, -73, -128, 44, 127, 22, -128, 5, 58, 127, -95, 127, 48, -96, -128, 127, 111, -78, 16, 76, -128, 42, -119, -128, 98, -53, -31, 101, 52, 8, 74, -106, -128, 88, -33, -2, 34, 98, -128, -60, 96, 58, 127, -128, -128, 29, 127, -98, -87, 0, -128, -16, 127, -87, -43, -85, -23, 107, 63, -128, -128, 124, 127, -128, 45, 127, -128, -78, -45, 58, 55, 28, -86, -128, 22, 127, -124, 22, -128, 78, -88, 80, 49, -59, 7, -128, 8, 127, 45, -128, 49, -23, -128, 37, 127, 117, -128, 88, 52, -128, 127, 79, -128, -53, 22, -24, 127, 127, -123, -23, 98, -128, -119, 127, 127, -18, -42, 15, -128, -128, 114, 66, 90, -69, -128, 74, 127, -128, 24, -32, -112, -128, 101, 127, -52, 109, 73, -128, -78, 58, 127, -81, -68, 63, 63, 65, 33, -128, -128, -69, 127, -124, -8, 92, -128, -7, 60, 21, 64, -108, -108, -128, 127, 59, -58, -98, 43, 127, 39, -128, -128, -50, 88, 97, 69, 23, -36, -107, -55, 127, 107, -49, -128, 60, 127, 12, -128, -116, 127, -76, 26, -108, 36, -6, 127, -128, -37, -11, 127, -128, 69, -79, -10, 127, -55, -128, -88, 127, 127, -74, -88, -76, -128, 127, 127, -128, 74, -79, -21, 112, 127, -128, -37, -128, 37, 127, 0, -128, 127, -7, 91, -54, -33, -34, -34, 12, 96, -65, 85, 127, 78, -81, -47, -36, -92, -114, 93, 29, -76, -128, 53, 127, 43, -128, 27, 52, -121, 127, 90, -112, -128, 127, 15, 116, -128, -8, 123, 87, -128, -47, -26, -50, 3, 127, 79, -128, 71, -100, 0, 71, 69, 78, -128, -128, 95, 66, -128, 48, 127, -88, -45, -71, 88, 127, 73, -128, -128, 88, 127, 75, -128, 42, 127, 16, -128, 69, 29, -128, -17, -17, 127, 52, 106, -96, 2, 0, -128, 16, 29, 107, -128, 27, 127, 78, -128, -70, 117, -124, -128, 127, -38, -3, 59, 93, -98, -128, 107, 127, -91, -128, 21, 28, 71, -102, -27, 90, -111, -128, 78, 43, 102, -74, -128, 53, -11, -128, 81, 127, 127, -128, -128, 37, 55, 107, -76, -33, -63, 127, 127, -63, -128, 45, 127, -43, -128, 122, 1, -124, 106, -128, 33, -92, 102, 60, 43, -128, -128, 96, 127, 22, -128, -96, 0, 52, 127, 127, -128, 88, -128, -11, 32, -21, 5, -79, -8, -17, -5, 127, -17, -128, 90, 64, -128, -128, 95, 91, 76, -86, 127, -109, -128, 79, 127, -128, -113, 124, 127, -128, -24, 86, -107, -95, 2, 127, -128, 91, -111, -128, 49, 127, -12, -49, -128, 52, 24, 65, -1, 23, -2, -109, -128, 5, 127, 127, -48, -128, -69, 127, 45, -59, -92, 127, -11, 88, 78, -47, -128, 127, 42, -32, 29, 69, 88, -95, -2, -106, 55, -107, -15, 127, 24, -128, 55, -45, 23, 121, -128, 17, -6, 100, 127, -24, -128, -128, 127, 127, 92, -128, -31, 8, 8, 108, -42, -128, -3, 127, -66, -37, -48, -95, 113, -49, 127, -54, 127, 12, -128, 44, 38, -48, 127, -11, 100, -85, -44, -55, 36, 43, 127, 48, 127, -128, 42, -69, -128, 79, 121, -128, 127, 127, 13, 96, -117, -31, -60, 50, -128, 127, 45, 127, -59, -128, 47, 127, 97, 0, -128, 13, 127, 49, -128, -1, 121, -92, -92, 52, -11, -18, 90, 70, 91, -128, 59, -92, -64, 127, -23, -123, 127, -45, -10, -49, 103, 87, 23, -128, 127, -16, -38, -10, 102, -34, 28, -68, 78, 127, -93, -128, 100, 127, -23, 49, 103, -128, -88, 127, -18, -66, -66, 127, -13, 53, -86, -128, 70, 98, 66, -69, 86, -128, 54, 5, -128, 45, 127, 74, -113, 90, -22, -59, 90, -86, -128, 127, -28, -98, -11, -59, 127, -12, -128, 12, 127, 39, -128, 107, -75, -128, 71, 127, 52, -43, -3, -98, 13, 28, -34, -128, 127, -88, -34, 127, -55, -128, 60, 127, -43, -128, -28, -86, 37, 127, 127, -128, -71, 127, 11, -128, -53, 127, -68, -128, 63, 21, -128, 71, 127, 60, -128, -107, -53, 111, 127, -128, 54, 127, -128, -112, 33, -70, 112, 37, -128, 127, 78, -7, -44, 52, 60, -119, 85, 111, 127, -128, -128, 127, 93, 8, -31, 3, 12, -121, 127, 26, -38, -47, -6, -100, 127, 44, 57, -34, 27, 26, 127, -79, -128, 127, 76, -63, -98, 71, 127, 55, -128, -128, -86, 127, 127, -118, 39, 39, -22, -116, -2, -21, 127, 127, 36, -128, -111, 127, 97, -128, 127, -37, -26, -17, 43, 107, -48, -119, -128, 127, 76, -107, 34, 127, -13, -128, -128, 127, 97, -128, -112, 127, 127, 93, -128, -103, 65, 55, -81, -128, 55, -88, 32, 45, -119, 127, -31, 127, -128, 127, -13, -36, 75, 33, -128, -128, 55, 127, -71, 127, -109, 32, 93, 11, -66, -128, 17, 127, -12, -128, 127, -69, -98, 127, 5, -128, -108, 127, 127, -7, -122, -128, -12, 127, 22, -128, 127, 10, 127, -128, -49, 127, -69, -128, 127, -12, 32, -36, -128, 127, 34, -128, 127, -11, 107, -7, -128, 127, 54, 81, 100, -128, 21, 24, 21, 127, -57, -95, -128, 127, -128, 100, -69, 45, 70, -128, -15, 127, -127, -64, 86, -54, -7, 118, -81, 127, -109, -15, 127, -128, -87, 127, -74, -118, 127, -123, -93, -121, -73, 127, 71, -128, 15, 109, 12, 38, 64, 48, -74, -92, 101, 127, -107, -36, -52, -38, -128, 127, -17, 17, -15, -52, 27, 8, 127, -44, -128, 58, 18, 10, 13, -100, 68, 127, -42, -128, -128, 66, 127, -58, -48, -81, -128, 127, 10, 57, -114, -33, -32, 127, -16, -71, 103, 65, -102, -74, -33, 127, 3, 49, 34, 127, 111, -128, 17, 37, -88, 100, 121, -119, 12, 59, -95, -102, 55, 38, -45, -128, 119, 127, -91, 127, 65, -128, 6, 68, 109, 127, -106, -128, -54, 81, -13, 127, -7, 127, 43, 127, -128, -128, -38, 101, 127, 81, -128, -116, -39, -7, 127, 127, -119, -128, -38, 127, 106, -103, 24, 22, -37, -128, 92, 45, -10, -76, 90, 111, -128, -111, -128, 127, 65, -128, 96, 57, 76, -112, 16, 48, -91, -102, -123, 101, 127, -50, -63, 91, -128, -50, -71, 127, 2, -45, -128, 101, 127, 70, -128, -44, 127, -128, -101, 127, 47, -90, 65, -29, 2, -128, 127, -17, 127, -128, -49, 107, 127, -128, -128, 90, 127, -1, -26, -6, -58, 66, 127, 127, -128, 21, -128, 127, 6, -121, 22, 127, -15, -107, -80, -88, 127, 49, -50, -93, 64, 127, 127, -32, -128, -88, -21, 117, 127, -128, 101, 127, -85, 37, 0, -103, -128, 52, 127, -26, -128, 92, -13, 0, -122, -108, -128, 127, 127, -119, -128, 127, -21, -64, -128, 3, 127, 68, 53, -128, -122, 100, 54, -97, -122, 98, 127, 0, 44, -128, 32, -32, 127, -23, -128, 55, 127, -60, -122, 127, -73, -128, 54, 38, 127, 92, -128, 2, 64, -128, 113, 127, -70, 27, 71, -128, -100, 127, 69, -116, 75, -109, -64, -123, -8, 127, 75, -80, 92, -128, 48, -43, 63, -47, -78, -69, 29, 58, 2, -60, 127, -22, -16, 127, -29, -50, -128, 127, -108, 127, 32, -29, -92, 100, 13, 121, -128, -98, 74, 85, -128, 8, -2, 127, -128, -22, -128, 127, 127, -80, -96, 127, -128, 50, -128, 31, -17, 6, -93, 36, -103, 71, 127, -128, -123, 127, -6, -128, 127, 38, -73, -2, 107, 27, -101, 10, 13, -128, 127, -87, 60, -33, 37, 127, -106, -128, 37, 127, -50, -128, 28, -21, 15, 57, 0, 11, 65, 68, -39, -58, -128, 127, 127, -68, -36, 95, -79, -48, 127, -87, -128, -2, 44, 127, -95, -50, 127, -37, -128, 34, 53, -116, -100, -128, 127, 96, 101, -128, 17, 103, 44, -71, -128, 96, 127, -113, -17, 127, -128, -98, 39, 127, -128, -96, 76, 87, -33, -128, 1, 59, 58, -128, -36, 37, 42, -128, 37, 80, -79, 127, -73, 6, 127, 59, -128, 100, -42, -128, 39, 127, 1, -128, -43, 127, -68, 79, -31, 127, 1, -128, -28, 112, -108, 127, 23, -70, -88, 31, 127, 80, -128, 73, 127, 96, -1, -128, 55, -128, -128, 12, 127, -91, -44, -5, 127, -8, -128, 127, 2, -13, -53, 90, 37, 54, 55, -79, -49, 112, -63, -50, -85, 127, 74, -128, -44, 127, 10, -47, -3, -70, -7, -86, 63, 70, -13, 13, -128, 47, 127, -128, -66, 2, 11, 0, -3, -128, 65, 124, -128, -34, 127, -128, -128, 127, -38, 1, -36, 15, -78, 24, 47, -103, 73, 127, -92, -128, 127, 127, -32, -127, -57, -2, -7, 127, -128, -60, 74, 64, -113, -101, -18, 86, -8, 0, 127, 127, -52, -23, 13, -128, -64, 127, -21, -85, -37, 127, 55, -128, -103, 123, -65, 85, -17, -128, -128, -128, 127, 127, -5, -128, 28, 127, 6, -6, -26, 36, 23, -47, 3, -11, 127, -100, 90, -17, -28, 7, -79, 127, 107, -49, -124, 92, 114, 12, -100, -57, -116, -128, 114, 93, 80, 68, -68, -128, -97, 127, -22, -74, 127, -88, -13, -73, 75, 33, -119, -128, -27, 127, 70, -80, -38, 127, -128, -28, -59, 127, -11, -69, -15, -81, 127, 6, -34, 23, -76, 127, -42, -128, -65, 127, -38, -29, 10, -103, -128, 127, 127, -128, -55, 127, 32, -75, -128, -12, 127, -59, -107, 127, 123, -128, -128, 76, 127, -128, -122, 123, 96, 34, -128, 36, -75, 59, 127, -37, -128, 93, -43, -128, 87, 127, -27, -128, -65, 127, -12, 111, -114, 103, -128, 23, -34, 16, -128, 127, 127, -118, 109, -119, 43, -69, 127, -18, -128, -52, 81, 127, -53, 23, -106, 32, -73, 127, -96, 78, -128, -98, 80, 87, -33, 21, 18, -116, -29, 127, 92, 113, -58, -128, -31, 127, -6, 127, -116, 43, 49, -79, -34, -7, 108, -128, 127, 22, -128, -86, 127, 103, 2, -124, 127, 71, -128, -118, 127, 49, 17, 87, -92, -128, 127, -109, -92, 86, 127, -128, -53, 112, -91, -128, 59, 117, 26, 13, 50, -112, 106, 38, 23, -128, 127, -128, -128, 127, 66, -27, -128, -39, 64, 32, 38, 86, -70, -128, 127, -17, -96, 127, 55, -128, 123, 103, 24, -128, 65, 16, 106, -123, -64, 127, -71, -81, -106, -12, 127, -101, 50, 127, -111, -108, 127, 114, -128, 5, -109, 87, 27, 63, -26, 15, -95, 8, -124, 76, -21, -75, -3, 101, 22, -52, -128, -128, 127, 6, 0, -13, -1, 52, 97, -128, -21, 28, -68, 32, -6, 5, 36, -65, -128, -128, 127, -85, -47, -119, 127, -26, 52, -128, 114, -87, 85, 16, 127, -64, -128, 39, 23, 23, -59, 57, 127, -38, 45, -29, -128, 127, -127, 26, -50, 31, 127, -128, -114, 66, -128, 57, 127, -117, 17, -91, 31, 64, 76, 63, -128, -27, 127, 53, -128, 123, -103, 70, -114, -127, 38, 50, -79, 127, 98, -128, -52, 24, 127, -3, -116, -128, 2, 127, -17, -34, 127, -106, 26, -128, 69, -64, 127, -122, -15, 114, -128, 76, -64, 0, -44, -48, 88, 116, -63, -55, -128, 127, -69, -18, 88, 26, -64, -31, 81, -128, 127, 48, -34, -58, 28, 127, -128, -22, 121, 127, -114, -128, 122, 86, 26, 6, -45, 64, -128, 80, 119, -128, 3, 3, -113, 109, 127, -44, -79, -57, 17, -128, 22, 127, 127, 10, -65, -128, 111, -34, -128, 85, 101, -128, 27, 127, -13, -122, 16, -86, -45, 127, -86, -122, 47, -50, 117, -102, 65, 71, 127, -128, 22, -18, -85, -13, 85, 88, 12, -121, 127, 116, 93, 47, -121, -128, 76, 127, 34, -121, -63, 36, -128, 127, 27, 0, 59, 127, -119, -33, -59, -76, 122, 127, -128, -47, 127, -36, 109, -76, -93, 8, 8, 13, 127, -128, -128, 127, 2, -128, 73, -2, -60, 127, 65, -128, 57, 127, -52, -128, 66, -86, 127, -128, -6, 124, 52, -57, -122, 58, 10, -128, -86, 127, 127, -34, -43, -81, -101, -1, 28, -128, 5, 127, -1, -128, -70, 116, -88, 106, 127, -8, -65, 127, -63, -45, -22, 127, 3, -18, -28, -5, 127, -22, -128, 65, -37, -128, -95, 127, 127, 73, -128, 38, -3, 103, -29, 6, 10, 92, -128, -106, 127, 107, -128, 34, 127, -128, -60, 54, 127, -118, -69, -21, 44, -107, -111, -18, 127, -26, 5, 92, -128, -91, 15, 127, 42, -73, -128, 127, 39, 7, 127, -128, -91, 127, 66, -97, -49, -128, 93, -74, 107, -7, 0, -124, -12, -3, 127, -128, -59, -78, 127, -37, 6, -21, -128, 38, 127, 127, -128, -128, 124, 111, -22, -128, -58, 73, -63, -88, -113, 81, 127, -128, 127, 127, -97, -128, 124, -12, 127, 73, -113, 76, -12, 87, 127, -75, -128, 127, -39, -13, 127, -13, -128, -92, -28, 127, 0, -70, 127, 127, -48, -70, -128, 68, 109, 81, -16, 90, -128, -39, -80, -87, -2, 127, -65, -128, -128, 103, 127, -48, 93, -128, 127, -80, -74, 127, 11, 34, -98, -128, 124, 85, -128, -13, 22, -69, 127, -21, 0, 31, 11, -116, -92, 127, -97, 80, -128, 127, -127, 113, 12, 123, -128, -42, 45, -107, -3, 22, 121, 116, -43, -128, 80, 23, 75, -79, -18, -3, -65, 127, 10, 90, -128, -47, 127, -128, -128, -12, 127, 0, -128, -101, 107, 127, -23, -75, 11, -5, 48, -79, 27, 127, -36, -128, -36, 124, 24, -28, -2, 71, 127, -64, 65, 127, -45, 45, 119, -128, -128, 127, 127, -128, -85, 2, 90, 54, -36, 24, -27, 48, 90, 3, 127, 6, -128, 15, 78, -128, 64, 80, 42, -128, 98, 127, -8, -128, -100, 63, 127, 127, -128, 24, 58, -128, -101, 127, 79, -128, -128, 127, -128, 90, 109, -12, -128, 42, 47, 127, -54, -81, -75, 107, 127, -128, 33, -75, 85, -128, -73, 45, 38, -114, 80, 71, 127, -18, -128, 47, 127, 114, 63, -128, -49, -5, -85, 33, 127, 106, -128, -124, 23, 2, -37, -86, 24, -63, 13, -128, 127, -90, 95, 11, 45, 12, -75, 52, -116, -12, -33, 127, -59, -71, 22, 65, -107, 74, 127, 28, -128, 66, 127, -49, -128, -128, 44, 127, 127, -128, -128, 93, 10, 28, 49, -128, -87, 127, -28, -128, 49, 16, 127, -16, -97, -106, 68, 127, 0, 32, -128, -57, -65, 121, -28, -55, -98, 127, 43, -128, 44, 127, 15, -91, 117, 70, 93, -13, -22, 127, 21, -80, -108, -15, 127, -58, -128, -39, -2, 127, 111, 31, 7, 127, 8, -128, 48, 47, 127, -128, -15, 127, 50, -128, 59, 70, -55, -109, 86, -47, 127, 127, 8, -86, -5, -128, 71, 127, 23, 11, 0, -127, -128, 127, 24, 38, -90, -28, 100, 43, 53, 92, -128, -121, 66, 127, -48, -122, -74, 127, 27, -128, -119, 27, -52, 127, 127, -8, -128, 127, 88, -128, 127, -7, 65, -128, 127, 5, -128, -96, 98, 127, 63, -128, -128, 127, 127, -27, -109, -59, 79, 127, 127, -128, -49, 127, -11, -128, -68, 127, -21, 33, 6, -111, 127, 96, -34, -76, 90, -69, 65, 81, 75, -128, 88, -128, -128, 127, 127, -128, 15, 127, -54, -128, 108, 127, -128, -100, 86, 75, 26, -52, -128, 127, 88, -97, 111, 127, -128, 8, 127, -127, -127, 60, -5, -43, 52, -57, 127, -128, 97, -31, -68, -128, 127, 127, 88, -128, -8, 127, 44, -78, -55, 90, -128, 98, -29, 49, -39, -68, -17, 127, -81, -39, 127, -80, -66, -24, 127, 79, -64, -128, 121, 127, -55, -118, 31, -55, -112, 127, 127, -65, -108, 103, -86, -107, 3, 85, 21, 112, -128, 100, 127, -32, -101, 88, 31, -116, -69, -6, 127, -28, 107, 116, -49, 127, 10, -128, -69, 127, 127, -128, 28, 127, -59, 47, -52, -128, 127, 127, -81, -10, -31, -90, -53, 127, -128, 21, -128, -33, 127, -128, 8, 127, 13, 54, -128, -128, 86, 87, 127, -128, -128, 39, 127, -29, -128, -128, -45, 127, -69, -107, 103, 127, -128, -128, -128, 47, 127, 16, 0, -90, 13, -37, 127, -128, 85, 80, -73, -42, -128, 127, 127, -29, 1, 0, 96, -64, -128, 127, 87, -57, 53, 91, -78, 50, 127, -38, -85, -128, 127, 127, -44, -54, -33, -38, 3, -34, -8, 127, 127, 29, -128, -128, -36, 127, 101, -128, -85, -5, 3, 127, 13, -128, -37, 127, -8, -10, 10, -10, 127, 70, -57, -128, 127, 127, -106, -27, 58, -18, -57, 117, -128, -128, 16, 15, 103, 96, -59, -128, 48, -2, 64, -8, -57, 127, 127, -106, -128, 43, 49, 80, 127, -116, -128, -128, 49, 127, 0, 60, -128, -47, 127, 98, -16, -122, 78, -128, -2, -128, 87, 111, 66, -109, -78, 32, -87, 22, -65, -128, -128, 122, 127, 127, -54, -128, 29, 114, 5, -71, -128, 122, 127, 127, -88, -96, -128, -59, 127, 49, -69, -44, -128, 68, 45, -31, -74, 127, 127, 0, -127, -17, 88, -5, -48, -128, 112, -107, 127, -123, 74, -8, 127, -39, -128, 88, 32, 34, 74, 13, -117, 65, 127, 93, -48, -128, 53, -65, 127, 127, -74, -128, -42, 127, 13, 127, 6, -128, 44, 64, -101, 127, 106, -128, -39, -28, 124, 127, -109, -85, -2, -24, 127, 49, 37, -128, 127, -54, 2, 88, 118, -37, -128, -128, -2, 127, 49, -117, 47, -97, -22, 127, -118, -128, 31, 127, 60, -128, 27, 127, -128, 44, 85, -92, 91, -36, -128, 112, 127, -50, -71, -68, -128, -10, 127, 127, -59, -128, 63, -26, 127, -22, 32, 0, -64, -128, 80, 127, 96, -128, -69, 28, 55, -128, 91, 127, 8, -38, -1, -128, 116, 1, -2, -124, -71, 127, 127, -26, -128, -55, 127, 50, -128, -52, 65, 127, -5, -128, -3, -27, 2, 107, -128, -128, 127, -53, -11, -93, -27, 78, 127, -90, -102, 21, -45, -55, 127, 3, 39, -8, 124, 17, -128, -128, 10, 127, 27, 127, -11, -128, 127, 44, -128, 113, 6, 91, 63, -16, -6, -128, 57, 101, -127, 0, 93, -71, 11, 33, 127, -44, -128, 5, 127, 127, -128, 33, -128, -37, 57, 21, 16, -108, 114, 107, 18, -23, -3, -128, 50, 5, 127, -128, 76, 101, -103, -112, 127, 103, 127, -128, -128, 13, 127, -52, -128, -128, 127, 127, -128, -38, 81, 127, 8, -68, -80, -79, 80, 127, 63, 81, -111, -128, -128, 127, 85, -11, -75, -52, 127, 103, -128, -6, 127, 54, -55, -76, -50, -21, -81, -21, 127, 52, -10, 95, -42, -128, 34, 127, 43, -128, 38, 127, -116, -128, 127, -2, -13, -31, 127, 60, 79, -64, -7, -128, 127, 17, 22, -128, 112, 127, -38, -128, -47, 127, 93, 32, -90, -128, -71, 18, 127, 10, 17, -128, 127, 127, -97, -81, 127, -128, -3, 86, -118, -128, 127, 3, -112, 127, -70, 91, -128, 127, -128, 42, -50, 127, -124, -13, -36, 127, 22, -70, -128, 127, 33, 127, -70, -128, -33, 127, 103, -63, -128, -31, -91, 5, 108, 127, -76, -128, 86, -15, 127, 2, 26, -76, 90, -124, 127, 33, -128, 10, 5, 43, 34, 42, 127, -75, -80, -34, -128, 37, 127, 127, -128, 59, -128, -34, 127, -90, -43, 29, -128, 87, 122, 116, 37, -128, -128, -2, 127, -95, -128, 23, 0, -37, 127, 81, -2, -48, -76, 127, 127, -52, -128, 29, -3, -65, 127, -34, 5, -2, -37, -32, -128, 108, 127, -128, -50, -3, 127, -74, 98, -128, -68, 118, -101, -91, 127, 69, -128, -49, 127, -112, 0, -76, -90, -87, 109, 95, -5, -76, 33, 127, -128, 6, 127, -60, -128, 36, -23, 127, -103, -69, 127, 36, -128, 39, -37, 111, -3, 33, 127, -43, -128, -5, 127, -128, -128, 96, 127, -128, -109, -57, 127, -33, 48, -128, 121, 28, 55, 24, -128, -128, 127, 96, 44, -128, 27, -8, -57, 86, -71, -48, -50, 59, -128, -1, 127, -93, -128, 102, 57, -26, -128, 47, 127, 127, -112, -93, 127, -73, -128, 127, 39, -128, -103, 127, 107, -117, -10, 12, 127, -128, -107, -75, 23, -60, 117, 127, 16, -128, 27, 127, 87, -128, -128, 71, 122, 5, 95, -128, -128, 127, -34, -128, -28, 27, 100, 127, -65, -128, -11, 74, -75, 28, 58, -128, 76, 95, -128, 15, 23, 1, 28, 127, 50, -15, -91, 1, -128, 58, -128, -128, -128, 127, 52, -128, 127, 127, -128, -128, 127, 28, 49, 76, -128, 7, 127, -90, -128, 95, 108, 116, 78, -92, -128, -17, 127, 113, -128, -37, 23, -97, 127, 127, -109, -103, 127, 68, -111, 29, -32, -68, 112, 127, -128, -5, 107, -48, 80, -128, 86, -11, -128, 57, 127, 127, -90, -101, -53, 36, -31, 76, -106, -128, -2, 127, 7, -128, -22, 119, -57, -2, 127, 38, -128, -13, -1, 98, 127, 127, -69, -128, -128, 114, 127, 81, -128, -6, 127, 102, -16, -128, -119, 127, -52, -86, 88, 27, -112, 101, 32, -21, 6, 127, -107, 26, 127, 127, -33, -128, -27, 127, -74, -128, 76, 66, 27, -128, 127, -26, 127, -90, -15, -5, 127, -95, 1, 37, -128, -53, 10, -45, 26, 127, -68, -8, -47, 36, -31, -11, 127, -128, 100, -128, 92, 31, 11, 21, -119, -128, 127, 127, -93, -128, 26, 127, -127, 127, 32, -15, -128, 102, 127, -68, -128, 98, 127, -65, -85, -6, -85, -68, 68, -68, -101, -11, 57, -128, -119, 127, 2, -128, 127, -59, 69, -7, -6, 28, 127, -128, 5, -57, -128, 65, 127, -113, 17, -90, -38, -45, 127, 127, -36, -128, -86, 127, 55, -128, -87, 127, -21, 8, -95, 127, -128, -31, 127, -101, -128, 127, 127, -128, -128, 100, 127, -44, 85, -128, -65, -91, 58, -52, 103, 127, -108, -128, 87, 45, 90, 63, -128, 65, 127, 70, -128, 0, 112, -11, -32, -43, 127, -55, -8, -102, -12, 66, 127, -128, -63, 127, -43, -78, -69, -128, 100, 12, -74, 127, 127, -128, -71, 127, -60, -96, 47, 127, -24, -11, -18, -50, 3, 54, 15, -59, 97, -128, 24, -128, 34, 127, -11, -128, -81, 127, 127, -118, -128, -50, -47, 44, 127, -80, -49, -37, 98, -128, 23, -75, 78, 127, 121, -74, -128, -79, 60, -12, 45, 127, -92, -18, -74, -64, -42, 118, 127, -81, -113, -128, 97, 127, -50, -128, 127, 44, -90, 45, 127, 102, -128, -81, 127, -74, -128, 114, -24, -128, 127, -44, -113, 21, 54, 97, -128, 127, 8, -128, 85, -88, 127, 37, 18, -128, 127, 48, -128, 127, 33, -128, 127, -79, 31, 127, -128, -37, -1, 112, -36, 24, -128, 127, -2, 127, -118, 127, -42, -128, -27, 127, -58, -17, 10, 127, -27, -128, 50, 31, 66, -17, 87, -53, 68, -93, -87, -22, 66, -75, 88, 123, -75, 113, -17, -128, 71, 127, -128, -39, 52, -109, 86, 42, 11, 106, 24, -73, 116, -107, 28, 124, -128, 121, -81, 108, 22, -128, -76, 127, 88, -128, -128, 90, 127, -78, -128, 71, 127, 90, -128, -11, 29, 101, -79, -128, 127, -128, 127, 1, -80, -128, 127, 127, -122, 86, 127, -98, -73, -58, -79, 127, -49, -128, 48, 106, 28, 100, -128, -128, -29, -7, 117, 127, -22, -128, 127, 76, -128, 52, 13, -85, 103, -48, -49, 127, 116, -128, -128, 109, 123, -65, 11, -86, -21, 127, 63, -128, 42, 81, 66, -128, 21, -43, 127, 92, 58, -128, 127, 127, -102, -18, -128, 116, 127, 52, -121, -88, 21, -57, 127, -37, -128, 111, -7, 122, -23, 18, -108, 38, 127, -116, -128, 55, -80, 118, 98, -128, 5, 127, 127, 24, -45, -93, -128, 90, 48, 58, -65, -50, 123, 127, 78, -128, 27, 1, -128, 124, 42, 109, -33, 12, 127, -69, -128, -128, 127, 78, -13, 127, -128, 58, -54, -128, -7, 127, 91, -128, 118, -66, 5, -45, -34, 86, 127, -128, 127, 26, 12, -23, -117, -38, 127, -28, -128, -26, 97, 31, 12, -100, -24, 34, -128, -13, 38, 74, -124, 64, 119, -11, -31, -6, 23, 13, -7, -43, 0, -32, 127, -33, 55, 127, -123, -81, 127, -22, -128, -37, -57, 96, 32, -54, 27, 28, 111, -5, -57, 43, -13, -128, -98, -128, 73, 127, 7, -100, 127, -128, -114, 92, 127, -73, -128, 60, 127, 2, -128, -57, -106, 127, 47, 95, -5, 98, -128, -63, -128, 127, 127, 50, -44, -38, 8, -111, -128, -128, 127, -6, 18, 2, -21, -128, 76, 127, 45, -128, 127, 74, -114, -128, 127, 107, 127, -128, 0, 37, -128, 109, 17, -68, 127, 74, -128, -90, -3, 81, -58, 29, 123, -128, 29, 0, 86, 34, -39, -128, 85, 127, 127, -128, -111, 127, 127, -128, -128, 15, -107, 127, 13, -71, -73, 118, 47, -28, 76, 15, -7, -42, -76, 50, -128, 127, -60, -52, 91, 127, -128, -128, 91, 127, 76, -128, 59, -52, 121, -60, -28, -119, 113, 86, 127, -15, 21, -7, -128, 70, 65, 66, -58, -128, 127, 98, -127, -118, 60, -71, 127, -48, 127, -128, 101, -87, 127, -128, -128, 70, 118, 90, -128, -128, 100, 127, -76, -128, -69, 127, 8, -128, -73, 112, 119, 32, -98, 127, 119, -36, 5, 59, 0, -128, -118, 127, -75, -128, 58, 127, 71, -128, -128, 127, -21, -5, -16, 127, -100, -128, 26, 39, 80, 127, -128, -87, 100, 57, -118, -59, -52, 122, -12, 109, -79, 119, -128, 100, -128, 127, 13, -121, -85, 127, 36, -97, -21, -16, 78, 1, -128, -26, 124, -71, -128, 127, 63, 38, -86, 57, -100, 88, 78, 23, -128, -128, -96, 127, 95, -21, 16, -22, -70, -128, 69, -66, 80, 8, -128, -39, 127, 127, -128, -128, -48, 127, 59, -128, -128, 114, 71, -22, 31, 59, -45, 127, 1, 65, 95, -117, -48, 95, 5, 127, -128, -11, 127, -63, 49, -128, -1, -128, 127, -111, 93, 50, -128, -42, 127, -93, -37, -93, -53, 22, 8, 24, 58, -128, 127, 87, -23, -128, -10, 127, 127, -128, -128, 93, -93, 127, 5, 90, -128, 3, 127, -42, -128, -108, 127, 5, -91, -27, -65, 100, 127, -57, 24, -15, -50, -85, -11, -29, 121, -98, -119, -27, 127, -128, -59, 112, 76, -128, 81, -47, -128, -16, -70, -18, 127, 124, 71, -128, -128, -24, 71, 18, -59, -21, 18, -128, -96, -128, -50, 127, -8, -66, -8, 12, 52, 127, 81, 34, -128, -53, -78, 127, 60, -128, 86, 127, -128, -38, 36, -128, 81, 96, -34, 23, 71, -48, 44, -98, 127, 24, -26, -42, 124, 101, -128, 64, 111, 87, 7, 43, -128, 127, 42, -26, -49, -22, -70, 127, 90, 127, -88, -128, 66, 127, 98, -128, -90, 127, -21, -128, -68, 127, -49, -18, 1, 7, -5, -32, -128, -124, 28, 55, 0, -128, -86, -128, 127, -39, -32, 124, 71, -54, -128, 127, -53, -128, 127, -29, 39, 36, 127, -128, -128, 119, 127, -128, 112, -33, 26, 44, 127, -7, 7, -128, 47, 57, 49, -128, 52, 91, -128, 70, -68, 68, 11, 127, -128, -123, -81, 29, 127, -21, -128, 127, 24, -128, -128, 127, 26, 127, -12, -128, 43, 10, -24, 127, 52, -128, 86, -108, -44, 92, 127, -64, -69, 127, -31, -128, 37, 98, -55, -18, 127, 127, -1, 28, -128, -57, -5, -1, 127, -33, -128, 103, 127, -128, -103, 93, 127, 48, -16, -101, -128, 96, 69, 88, 50, -113, -102, -43, 127, 49, -63, -44, 119, 13, 127, 13, -7, 127, 39, 2, -8, -101, -13, 127, 97, -128, -128, 97, 114, 122, -111, -118, -44, -58, 127, -22, -85, 0, 6, 21, 23, -11, -11, 127, -128, -128, 116, -3, 127, -121, -128, 63, 127, -128, 49, -59, 43, -29, -48, 127, -128, -48, 127, -128, -128, 116, 27, -45, -76, -128, 86, 127, -7, -102, -128, 109, 127, -121, -128, 74, -1, 8, 127, 92, -128, -128, 31, 65, 22, 57, 79, 7, 70, 127, -128, 60, 54, -71, -118, 127, -22, 49, -64, 12, 47, -15, -49, -128, -13, 101, 55, -7, 37, -45, -128, 3, 127, 34, -128, -29, 127, -6, -128, -107, 127, 127, 16, -128, -128, -128, 127, 127, -45, -44, -65, 109, -32, -128, -23, 127, 69, 54, 58, -128, -128, 3, 127, -68, -90, -97, 76, 74, -128, 98, -107, 60, 7, -128, -47, 127, -86, -128, 127, 80, -128, 127, 73, -128, -65, 55, 127, -21, -11, 127, 127, -128, -128, -6, 91, 127, 18, -128, 63, 6, -128, 102, -29, 58, 12, -74, -128, 127, -108, 0, 127, -87, -96, 127, -96, 59, -6, -44, -128, 127, 58, -128, 117, 87, 63, -10, -128, -34, 33, 127, -81, -98, 74, 101, -87, 79, -128, -36, -86, 2, 39, 54, -92, 63, 98, -15, 10, 127, -57, -128, 1, -17, 127, 16, -128, 69, 127, 42, -128, -128, 92, 127, 11, -107, 106, 34, 127, -128, -54, 127, 29, -106, 127, -63, 0, 59, -81, 60, 127, -58, -85, -74, -128, 127, 64, 96, -128, 24, 28, -52, -128, 127, -93, 29, 127, -17, -128, 78, 29, 28, 127, -128, 0, -43, -2, -114, 127, -58, 38, 127, -93, -76, -1, -81, 24, 127, -90, -119, 127, 127, -107, -128, 117, 127, -32, -128, 65, 52, -33, 44, -28, 68, -128, -33, 127, -128, 36, -128, -44, 127, -128, -22, 11, -6, -95, -31, 91, 29, 26, 73, 122, -128, -128, -5, 127, -128, -36, 123, 66, 127, -108, -128, 127, 90, -34, 1, -11, 78, -106, 43, 31, 59, 127, -128, -93, -28, 54, 127, -128, 42, -102, -60, 15, 112, -128, -55, 127, 76, -127, -81, 52, 6, 127, 27, -128, 98, -101, 103, -48, -44, 127, 39, -75, -128, 127, 127, -44, -128, 121, 57, 66, 81, 48, -128, 36, 45, -10, -60, 17, 88, 22, -68, 100, 127, 111, -108, 32, 45, -128, 42, 66, 52, -43, 123, -80, -114, -128, 7, 127, 73, -128, -47, 127, 98, -128, -128, 8, 121, -6, 0, 127, 18, -128, -78, 127, 75, -12, -21, 127, -128, -63, -128, 18, 127, 127, -128, -98, -48, 54, -78, -128, 38, 127, 71, -90, -128, 10, -39, 21, 127, 127, -116, -128, 90, 90, -52, -106, 127, -58, 24, -116, 69, -79, 127, -21, -128, -54, 127, -38, 39, -113, -111, 36, -7, -43, 127, -33, 74, 31, -128, -80, 127, -95, -53, 127, 127, 13, -128, -128, 127, 60, 65, 114, -128, -93, 107, -37, -128, 24, -50, 73, 112, -88, -108, 127, 26, -116, 127, -53, -128, -16, -8, 71, 127, -65, -128, 34, 127, -98, -23, -54, -128, 127, 127, -26, -114, 75, 103, 13, -43, -122, 87, 117, -128, -86, 12, -2, 127, -45, -128, 65, -37, -65, 75, 97, -128, -31, 127, -79, -111, 27, 113, 16, -109, -2, 127, -128, -128, 127, -128, -32, -50, 17, 101, -80, -128, 65, 74, -18, 91, -128, -128, 69, 102, -109, 33, -11, 47, 50, -128, -100, 66, 64, 112, 49, -128, 34, 18, -117, -128, 95, 127, -128, -101, 78, -60, -128, -91, 127, 127, -69, -66, 127, 127, -87, -24, -128, 100, 127, -12, -86, -47, -66, 127, 127, 44, -23, -42, -128, -128, 127, 127, -128, 7, 31, -100, -128, 27, 127, -85, -128, 114, -15, -101, 31, -54, 113, 47, -111, 73, -37, -36, -26, 65, -128, 111, 18, -23, -65, -38, 42, 48, -36, 127, 127, -128, -17, 122, -54, -128, 127, 73, -65, -49, 127, -86, 121, -93, 29, 43, -27, -128, 22, 42, 78, 127, -2, -128, -18, -23, 127, 63, -98, 63, 127, 127, -128, -98, -128, 116, 127, -7, -128, 127, -78, -18, -23, -33, 33, 93, -92, 95, 127, 127, -128, -66, 2, -24, 127, -107, 12, -123, 127, 18, -7, -17, -59, -27, -34, 127, -97, -128, -47, 127, -78, -47, 54, 127, -109, 1, 71, 60, -16, 44, -15, -128, -128, -88, 119, 127, -128, 127, 81, 17, -58, 18, 88, -128, 2, 68, 52, -109, -112, 127, 127, -128, -2, -111, 22, 52, -2, 28, -128, 12, -16, -128, 85, -38, 13, 43, -128, -128, 100, 101, 2, 55, 2, -102, -101, 1, 39, -64, 49, 127, -86, -117, -128, 127, 127, -75, -64, -128, 53, 127, 106, -18, -128, 97, -128, -53, -45, 127, -128, -13, -128, 127, 59, -80, -128, 108, -55, 90, 127, 70, -128, 114, 79, 74, -114, 21, -26, 52, -73, 69, 5, 2, 127, -7, -128, -95, 127, 48, -122, -128, 127, 127, -128, 113, -128, 8, 22, 127, -128, -2, -26, 23, -34, -12, -73, -33, 127, -86, 53, 119, -8, -87, 68, -45, 127, -128, -128, 2, 127, 92, 43, -128, -75, 127, -3, -71, -36, 100, -85, -13, -127, -74, 88, 97, 11, -128, -15, 127, 127, -128, -79, 127, -39, -65, -90, -111, 127, -86, 127, -122, -91, 58, 127, 85, -39, -128, -119, 17, 119, 22, 71, 60, -119, 0, 0, -53, 66, 127, 88, -128, -15, 127, -128, -63, 127, 31, -91, 29, -86, -66, 68, 11, 127, -24, -128, -39, 127, 98, -128, -128, 101, 75, 101, -116, 33, 127, 38, -116, -128, 37, 108, 127, -128, -128, 127, 1, -78, 68, 31, 50, -81, -128, 127, 127, -37, 55, -128, -5, 127, -27, -107, -45, 10, 21, -116, -23, 127, 49, 60, -128, -49, -12, -13, -128, 42, 127, 91, -111, -38, 116, 52, -39, -71, 100, -128, -128, 127, 78, 75, -128, -37, -128, 127, 52, 76, 37, -128, 88, 49, -128, 44, 127, -128, -128, 127, -26, -128, -37, -103, 127, 127, 6, -128, 78, -65, 112, -116, -128, 39, 127, -1, -121, 70, 29, 66, -106, 87, 12, 127, -87, -128, 108, 7, -13, 44, 33, 69, 127, -128, -22, 127, -44, -128, 28, 15, -71, 59, 127, 127, 17, -128, 13, 124, -66, -33, -64, 68, 127, -63, -128, -38, 57, 38, 28, 27, -11, 127, 88, 90, -88, -26, -128, 85, 13, 29, 127, -128, 38, -128, -5, 116, 127, -128, -68, 27, -128, 86, 5, -27, -52, 31, -33, 122, -128, -128, 69, 127, 53, -128, -32, 55, 24, -128, -10, 71, 127, 37, -98, -113, 78, 44, 73, -128, 75, -36, 122, -1, 100, -47, -101, 127, -128, -23, 127, -24, -128, -52, 21, -15, 42, 127, 127, -123, -128, 127, 11, 102, -128, 8, 127, 127, -128, -42, 1, 127, -74, -128, 88, 127, 70, -128, -44, 108, -128, -113, 45, -71, 3, 79, -36, 47, 75, -48, -128, 87, 127, 90, 28, -128, -28, -88, 32, 127, -114, 21, 87, -90, -128, 17, 127, 85, -91, -128, 28, 127, -12, -128, -52, 127, -18, -128, 127, 118, -22, -74, -7, 26, -36, 127, 6, -68, -2, -17, 27, 6, -2, 63, 108, 48, -128, -122, 13, 127, 18, -128, 101, 127, -128, -116, 127, 98, -128, 70, 0, -95, 39, -64, 93, 69, -18, 7, 49, -23, -34, 127, 86, -24, 49, 47, -128, 69, 127, 127, -102, -128, -60, -10, 127, 127, -80, -111, -60, 127, 22, -128, 3, -11, 53, 127, -90, 85, -11, -128, 60, 97, -66, 5, 97, 66, -88, -38, -128, -31, 127, 52, 26, -70, -119, -128, 127, 127, -12, -128, -81, 47, 58, -12, 66, -43, 71, -13, -45, -128, 127, -12, -75, -128, 127, 127, 103, -128, -52, 127, 2, -128, -52, 90, 127, -70, 49, -34, -128, 127, 54, 107, -86, -53, -22, 127, -123, -123, -65, 101, -13, 79, 69, 122, -123, -53, 58, 13, -128, -1, 118, 18, -58, -116, 127, 127, 63, -97, -58, -58, 127, 108, 38, -36, -128, -44, 127, -96, -38, 59, -44, 11, 127, -81, -50, 127, -80, 13, -128, 48, 92, -24, -18, -49, -32, 71, 38, -55, -36, 68, -128, 7, 127, -91, 10, -32, -128, 45, 127, 39, 37, -48, -128, -128, 127, 127, 66, -31, -49, -127, -38, 127, -45, -128, 48, 127, 74, -128, 78, -102, 127, 17, -128, -15, 127, 58, -128, -86, 127, 10, 58, -128, 44, -128, 34, 118, 47, -98, -128, 127, 127, -116, -128, 11, -29, 127, -58, -97, 36, 127, -80, 58, -128, -128, 122, 127, -39, -127, 24, -128, -13, -50, 127, 49, -128, 127, 31, 48, -128, 59, 127, 60, -128, -128, 112, 87, -103, -128, 73, 31, 12, 127, 127, -128, 60, 112, -128, 65, 15, -36, 59, 52, 31, 66, -128, 91, -33, 127, -108, -63, 127, 127, -128, -111, 50, -42, 127, -121, 7, -2, 43, -66, -102, 127, 53, -23, -52, -106, 6, 127, 87, 117, -128, -119, 48, 127, -128, 102, -128, 31, 95, 118, -128, -71, 127, -79, 0, 127, -26, -123, -128, -8, 127, 47, 5, -50, -128, 127, 109, 43, -106, -80, 95, 127, -128, -128, 127, -24, -128, 127, 11, -128, 124, 2, -60, -81, 127, -69, -74, -87, 127, -128, -33, 87, -87, -68, 119, -50, 65, -8, 107, -101, -128, 100, 127, -128, -13, 85, -91, -8, 127, -24, -128, 127, -33, -22, 124, -47, 33, -13, -128, 97, -128, 122, 43, 18, -128, -111, 127, 22, -18, -66, -128, 127, 127, -44, 65, -47, 103, -15, -49, -90, 73, -22, 127, 122, -128, -21, 127, -88, 50, -39, -128, -6, 38, 53, 116, 127, -70, -128, -109, 127, 66, -111, 33, 88, 98, 50, 28, -7, -13, 15, 1, -48, 127, -128, -34, 63, 122, -128, 1, -52, -32, 127, 10, 17, 5, 127, -102, -98, 24, -59, -26, -70, 127, 57, -7, -59, 2, 97, 127, -57, -5, -31, 50, -32, 127, -123, 55, 116, -98, 17, 59, -128, 0, 127, -128, -1, 66, -128, -75, 127, -87, 123, 33, -128, 85, -117, 127, 5, 78, -12, 33, -21, -128, -100, -128, 127, 127, -42, -128, -21, 127, 27, -73, 38, 121, -106, 16, 127, -92, -71, -12, 47, -33, -128, -32, 127, 88, -43, 71, -128, -128, 98, 127, 37, -128, -128, 127, 37, -13, -107, 75, 85, 127, -128, 17, 127, -13, -128, -128, 26, 127, 127, -128, -119, 100, -79, 78, -121, 71, -48, 91, -119, -2, -128, 127, 3, -106, -73, 23, 87, 0, 117, 122, 38, -29, -128, 37, 8, 36, 85, 127, -128, 11, -114, -26, 15, -128, 55, -64, 11, 127, -128, -32, -97, 60, 127, -128, -60, 38, -113, -123, 119, 127, 31, -128, -128, 90, 127, 44, -108, 127, -87, 12, -5, -95, -2, 38, 48, 29, -128, 32, -128, 121, 95, -128, -108, 127, 16, 48, -128, -22, 118, -29, -18, -128, 1, -90, 90, 127, -33, -128, 63, -10, -34, 101, 127, -128, -13, 44, 107, -128, -109, -36, 58, 127, 91, 0, -128, 2, 8, 5, -97, 76, 60, -8, 88, -23, -106, 103, -34, -22, 71, -2, -128, -128, 26, 127, -43, -29, -22, -128, 101, 127, -128, -39, 127, 76, -24, -103, 3, -38, 95, -106, 22, -128, 74, 127, -91, 11, 79, -10, -71, -47, 39, 127, 16, 96, -73, -128, 11, 127, -34, -128, -60, 95, -38, 31, -128, 48, 112, 118, -108, -32, 121, -107, -27, 114, -101, -128, -66, 127, -44, -128, 34, 102, -128, -7, -18, 127, -128, -128, -5, 127, 68, -49, -28, -1, -58, -128, -1, 127, -69, -128, 127, 7, -128, 78, 0, 66, -80, -101, 34, 127, 65, -128, -32, 10, -85, 127, 127, -128, -34, 127, -37, -128, -93, 127, -98, -66, 122, -128, 69, 106, 88, -78, -128, 36, 127, 0, -57, -87, -42, 127, 127, 102, -128, -128, 97, -22, -10, 127, -3, -36, 60, -6, -17, -91, -42, 53, 38, -33, -37, 127, 29, 100, -128, 52, -128, 26, 118, -107, -43, -5, -42, 127, -108, -128, -43, 70, -10, 127, 10, -118, 5, 123, -128, -81, 122, 97, -58, -128, 63, -54, 36, 127, -87, -128, -119, 127, 7, -128, -33, 17, 109, 15, -128, 127, -7, 127, -128, 70, -7, -128, 52, 123, 8, 66, -1, -128, -66, -36, 80, -36, 102, 127, -124, -31, 124, -128, -1, 5, 97, -21, 100, 23, -128, 28, 7, 22, 50, -34, -114, 71, 127, -78, 59, 127, -60, -118, -29, -2, -128, 127, -8, -63, -78, 127, -128, 127, -96, 127, -18, -127, 103, 39, 76, -75, -128, 118, 127, -43, -124, 15, 33, 18, 1, 49, 106, -96, -128, 43, -17, 127, -31, 66, -63, -101, 36, 59, -10, -128, 3, 50, -39, -128, 127, 100, -128, -128, 127, 127, -12, -74, 54, 45, -128, -128, 3, 127, 127, -128, -128, 127, 57, -80, -128, 17, 74, 58, -119, -96, 6, -128, 53, -117, -5, 102, -113, -128, 127, 0, -8, 42, 114, -3, -128, -128, 68, 34, -36, 127, 8, -128, -128, 127, 127, -128, -128, 111, 127, -128, -15, -15, 122, 101, -68, -128, -5, 127, -70, 23, 127, 33, -21, -47, 43, 53, 2, -128, -59, 113, -128, 86, -47, -128, 127, 42, 38, -60, 44, -128, 74, -128, 23, 121, -88, 0, -122, -117, 127, 95, -79, -95, -10, 59, -59, -37, 127, -15, -128, 91, 54, -18, 6, -111, -122, 127, 15, 27, 57, 12, -24, -87, 127, 60, 127, -128, -76, 127, -128, -68, 127, -128, -111, 127, 33, -128, -128, -47, 127, -5, 13, -5, 127, -5, -103, -128, 122, 127, 6, 127, -29, -128, 65, 112, 11, -60, 47, -128, 127, -73, 44, 34, -29, -111, 127, 66, -109, -128, 127, -18, -90, 60, 127, -49, -109, 0, 45, -128, -66, 36, -29, 113, 50, 122, -128, -54, -64, -68, 59, 122, -114, 0, 111, 127, -128, -119, 127, 12, -128, 127, -18, -100, -106, 127, -15, -98, -15, 127, -75, -128, -54, -81, 127, 100, -64, 15, 45, -7, -128, 127, -78, 79, -107, 127, -128, 79, -39, 127, -12, -128, -50, 127, -48, 3, -18, 127, 127, -128, -73, 43, 80, -128, 102, 43, 71, 98, -113, -44, 86, 111, -128, -98, 127, 112, -128, 118, -42, -22, 97, -87, 42, 13, -38, -85, -128, 102, 55, -81, 24, 127, -128, 36, -24, -113, 31, -24, 127, 43, -32, -103, 127, 100, -128, 2, 127, -75, 5, -64, -68, 11, 127, 88, -8, -128, -128, 127, 64, 60, -55, -13, 74, -128, -48, 127, -128, -6, -7, 44, -49, 127, -111, -128, 78, -1, -106, 127, -100, 78, 122, -128, -128, 127, 127, -128, -128, 92, 127, -1, -55, -29, -37, 127, 26, 18, -17, -128, -5, 37, 21, -81, 26, -12, 32, -32, -106, 127, 6, -128, 127, 39, -49, -42, -59, 80, 127, -128, 2, -66, 8, 10, 50, 37, 75, -75, -85, 127, -8, 36, 22, -116, -45, 52, 93, 127, -128, -102, -127, 85, 5, -18, 60, -64, -15, -128, 127, -93, 65, -50, 127, 63, -124, -128, 127, -3, -6, 71, -45, 71, 127, -128, -128, 55, -26, 78, -88, 127, -2, 8, -128, 93, 127, 80, -85, -128, 53, -121, 75, 127, 36, -73, -57, -52, -91, 13, -103, 11, -88, 59, -116, -65, 85, -128, 118, -106, 3, -6, 33, -6, -43, -75, 127, 17, -60, -128, 127, 27, 98, 43, 12, -119, -49, 22, 80, -101, 76, 65, -90, -22, -16, 34, 127, -12, -96, -114, 127, -128, 22, 127, -75, 49, 103, -128, -128, 127, 29, 15, -45, -34, 124, -59, 95, -1, 43, 18, -128, -33, 95, 55, -128, 8, 39, -2, -88, 78, 47, -21, -69, -50, -16, 69, -100, -128, -128, 45, 127, 76, -128, 127, -108, -55, 127, -29, -128, 127, 66, -17, 78, 68, -128, -128, 90, 17, -128, -21, 127, 29, -128, -128, 95, 127, -2, -18, 100, -87, 53, -128, 71, -43, -21, 127, -128, -36, 127, -42, -128, 69, 106, -38, 127, -128, 43, 43, 127, -37, -128, -97, 127, 90, 12, -128, -127, 34, -18, 37, 78, 15, 87, -39, -118, -3, -42, -128, 127, 119, -128, 52, 127, -118, -76, 52, -42, 44, -1, -122, -47, 127, 112, -116, -73, 127, 18, -18, -66, 127, 127, -128, -128, -18, 127, -31, 24, -92, -128, 55, 127, -98, -128, -109, 63, 119, 112, 123, -128, -128, 111, 73, 127, -128, 85, 107, -128, -57, 127, 21, -128, 118, 36, 6, -42, 127, 15, -90, 71, -13, -48, -128, -7, -106, 127, 127, -74, -81, -103, 32, 127, 59, -128, -87, 109, 34, -128, 127, -79, 85, -42, -128, 127, -43, 11, 93, 127, -109, -112, 10, -6, -128, -128, 112, 42, 42, 0, -128, -128, 127, -43, 121, 31, 11, -128, 127, 127, 0, -88, -70, 118, 118, -57, -81, 73, -128, 47, 127, 106, -128, 69, -6, -128, -34, 127, 127, -128, -13, 65, -103, 26, 127, -103, -128, 127, 109, -88, 13, 127, -128, -128, 65, 127, -128, 5, 127, -128, -15, 127, -76, -128, 80, 127, 66, 127, -128, -119, -76, 53, 11, 127, -97, -128, -53, 127, 102, -128, -121, -64, 69, 127, -92, -128, -78, 2, 127, -118, 37, 75, -90, -128, 127, -114, -95, 117, -47, 70, -34, -23, -128, 85, 18, 127, -128, -81, 13, 43, 98, -128, -113, 127, -121, -128, 127, -10, -98, -34, 107, -92, 92, -128, 85, 117, -93, 87, -80, -29, -102, 127, 107, -128, -128, 6, 127, -13, 93, -128, -128, 127, 29, -128, -11, 75, -10, 64, 118, -127, -117, 42, 68, 86, 38, -1, -98, 68, 73, -28, -100, 34, 108, 10, 108, -98, -123, -128, -48, 127, 127, -29, -80, -59, -81, -18, -34, -27, -37, 23, -10, -69, 66, -128, -38, 5, -21, 11, -12, -52, 66, -128, -128, -32, -127, 1, 127, 127, -128, -96, 127, 65, -112, -128, -53, 127, 49, -37, 32, -86, -18, -43, 127, -80, -128, 92, 37, 29, 12, 127, -128, -65, -55, 3, 88, 64, -17, -128, 47, 86, -128, -49, 127, 95, 48, -42, -128, 42, -28, -128, 79, 127, -128, 0, -109, 29, 26, 127, -128, -128, -43, 53, 102, 26, -128, 66, 49, -6, -69, 79, 122, -36, 6, -48, -3, 85, 81, -68, -17, 37, 96, -128, -117, -122, -16, 127, 93, -31, -70, 5, -23, -34, 127, 22, -128, 93, 45, 78, -1, -128, 10, 103, -42, -12, 127, -128, -53, 127, -64, -128, 64, -48, 127, 127, -42, -128, 122, 109, -65, -103, -73, 60, 127, 96, -128, -63, 127, -47, -128, 109, 81, -43, -13, 127, 39, 127, -65, -42, 71, -128, 127, 57, 29, -128, 63, 80, 55, -128, -37, 23, -98, 91, -128, -54, -71, 127, -37, -10, -88, 32, 127, -127, -108, -128, 127, -68, -50, 127, -75, -91, -5, -45, 36, 127, -113, 79, 127, -12, -128, -128, 127, 68, -23, 48, -11, -8, -22, 127, 127, 79, -128, -12, -78, 52, 127, 42, -128, -15, 111, 10, 2, 0, 112, 127, -128, -114, 69, -60, -24, 0, 21, -55, 124, 48, -118, 127, 26, -7, 127, -63, -128, -6, 127, 127, -128, -101, 127, -128, -81, 127, -118, -71, 95, -49, 38, -23, -80, -128, 127, 127, -97, -128, 95, -36, 127, -121, -128, -11, 108, 48, -5, -12, -42, 37, 127, 127, -22, 21, -15, -128, -128, 119, -54, 127, -69, 21, -128, 59, 78, 26, -128, -17, 33, 48, -16, 74, -68, 65, -80, -79, 119, 74, -128, -114, 98, -69, 86, -17, 127, 66, -128, 0, 5, 93, 65, 127, -113, -128, -37, 8, 114, 91, -128, -128, 0, 57, 122, -106, -5, 93, 12, -128, 68, 68, -68, -128, -64, 49, 127, 76, -128, -3, 127, -128, 21, 13, 7, -73, 73, 127, -128, -87, 101, -32, -39, -78, 71, -102, 22, 118, 127, -128, -63, -118, 52, 74, -128, -38, 127, -109, -128, 127, 93, -128, 63, 103, -108, -128, 127, 113, -128, 70, 127, -59, -128, 127, 95, 127, -97, -80, -117, 87, 109, -5, 34, -71, -107, 65, 27, 29, -128, 0, 127, 87, -128, 12, 38, 52, 45, -111, 92, 101, -91, -15, -63, 112, 127, 90, 71, -128, -80, 127, -128, -128, 127, 1, -31, -44, 98, 70, -128, 18, 37, -24, -36, 26, -26, 127, -58, -74, -8, -44, 127, -128, -55, 116, 24, -128, 10, -92, 8, 74, -29, 18, -10, -102, 127, 18, -128, -10, 127, 69, -128, -114, 80, 127, -128, 127, -128, 102, 6, -3, -98, 98, 47, -90, 8, -128, 107, -6, -128, -121, 127, 16, 5, -39, 26, 113, -44, -95, -128, 127, 113, -128, -128, 85, 44, 127, 48, -15, -128, 96, 3, -128, 124, -38, -128, -128, 127, 127, 127, 21, -100, -128, -28, 127, 11, 76, -114, 15, -54, 98, 88, 49, -37, -128, 73, -6, 127, -128, -32, 32, -113, 52, -15, 79, -81, 34, -54, 81, -128, -16, -75, -43, -128, 127, 116, -36, -87, -69, 55, 127, -43, -128, 127, 47, -36, 127, -128, -116, 38, 2, -128, 127, 1, -128, -10, 119, -128, 101, 127, 3, -101, 127, -128, -12, 58, -88, -91, 127, -7, -12, 22, -6, -55, 22, -37, 109, 7, 127, -27, 17, 28, -36, -58, 17, 112, -66, -28, 111, 22, 75, 127, -128, 23, 17, 0, -128, 127, -42, 96, -93, 48, 101, 31, -10, -15, 32, -87, -96, -57, 45, 42, -128, 127, 127, 127, -128, -128, 31, 127, -79, 28, -32, -45, -128, 32, 127, -15, -128, 127, 12, -128, -1, 101, 127, -128, -6, 86, -128, 54, 127, -128, -24, -26, 127, 65, -66, -55, 65, -39, -93, -10, -7, 54, 101, 127, -128, -36, -28, 15, -44, -97, 127, 127, -3, -74, -43, 127, 127, 70, 44, -28, -128, -106, 112, 1, 34, -116, 127, 85, -128, 0, 127, -128, -123, 29, 127, -128, -43, -98, 29, 123, -11, -32, -124, 12, 12, -65, 127, -128, 57, 53, -116, -5, 127, -70, -128, 127, -27, 127, -92, -65, -86, -95, 121, 127, 38, -98, 64, -128, -117, 127, -97, -128, 91, -16, 5, 101, -65, -128, 57, 127, -128, 55, 34, -68, 42, -27, 34, 127, -127, -107, -128, 34, 54, 64, -87, 44, 27, 26, -28, -128, -108, 127, 55, -128, 3, -124, 127, 127, 73, -128, -80, 113, 24, 78, 92, -128, -42, -12, 109, -12, -128, 127, 2, -13, 24, -114, 123, 22, 3, -113, 127, 127, -1, -128, 5, 127, -71, -128, -57, 121, 10, -128, 70, 127, -57, -43, -39, -37, 96, -128, 2, -101, 117, -17, 49, -80, 16, -74, -128, 127, 74, -10, -128, 127, 127, -112, -2, 107, -128, 29, 74, 6, -27, -50, 0, 73, 112, 60, 33, -103, 122, 127, -128, -18, 13, 47, 5, 36, -128, 102, -124, 88, 88, 48, 26, -93, -66, -15, -57, 100, -23, 127, -53, -128, -26, 127, 74, -43, -17, -128, -34, 13, 28, -128, -32, -33, 122, -3, 2, -68, -59, 127, 16, 95, 15, -80, -44, 13, -55, -42, 127, 127, -29, -73, -128, 118, 127, 78, 16, -123, -87, -3, -116, 12, 127, -122, 74, 5, 127, -128, 44, -10, 11, 5, -29, -27, 27, -28, -21, -128, -21, 127, 121, -109, -128, -128, 114, 127, 101, -47, -68, 65, 43, -2, -128, 107, 127, 1, 31, 85, -65, -63, -48, -106, 127, -103, -128, -102, 122, 42, 127, 7, -59, 81, -78, -6, 59, -80, -128, 127, 75, -11, -128, 93, 21, 123, -128, 45, -59, 127, -128, 119, -12, -85, 13, 127, -128, -128, 87, 90, 5, 13, -32, -128, -42, -43, -78, 108, 68, 127, -90, -128, -128, 127, -85, 78, -13, 113, -117, -128, 106, 109, 26, 127, -128, -74, 127, -128, -38, -112, 18, 38, 49, 101, -128, 47, -63, -107, -75, 127, -127, 127, -86, -21, 127, -37, -73, 8, 127, -128, -128, 42, 122, -57, -88, 127, -23, 39, 57, 127, -50, -128, -42, 127, 76, -128, -15, 80, -24, -49, 31, 55, -128, -128, -79, 127, 127, -70, -128, 127, 75, 44, -128, 69, 2, 58, 55, -128, -109, -103, 116, 49, 68, 74, 39, -128, 127, -64, -70, 53, 127, -128, -17, -108, -39, -36, 32, -69, 127, -128, 80, -128, 24, 127, -128, -85, 127, -50, -128, 0, 127, 68, -58, 47, 92, -101, -18, 127, 127, 5, -128, -128, 127, 49, -64, -16, 122, -80, -90, 21, -128, 127, 127, -128, 31, 127, -7, -102, 114, -112, -52, -102, 127, -70, -33, 57, -27, 127, -80, -128, -54, 87, 39, -66, 127, 127, -57, -128, -8, 127, 127, -128, -128, 117, 101, -11, -47, -45, -91, -128, 102, 55, -91, 96, 44, -128, 59, 73, 111, 97, -128, -92, -128, 127, -44, 43, 10, -26, -5, 127, -2, -128, 0, 73, -13, -107, 114, 127, 81, 16, -128, -128, -98, 127, 50, -128, 38, 37, -91, -17, 127, -53, -32, -95, 127, 43, 127, -128, -128, 54, -98, -2, 106, 127, -69, -33, -42, -58, 127, -37, 5, -59, 127, -91, -128, 79, 127, -128, -128, 52, 21, -8, -128, 127, -18, 58, 127, -69, -128, 37, 127, -78, 29, -87, -128, -5, 95, 15, -98, 119, -86, 97, 127, -128, 37, 88, -68, -93, -8, 23, 127, 44, -69, -128, 39, 127, 127, 64, -128, 45, 3, -113, -2, 3, 69, 127, -2, -128, 11, 119, -128, -63, 1, 44, -128, 98, -34, -128, 106, 127, 0, -37, 52, 127, -128, 66, 127, -100, -128, 127, -70, 66, -44, -128, -52, 127, -26, -128, 43, 127, 96, -128, -22, 49, 127, -128, 101, -128, -10, 57, 123, -74, -128, 87, -21, -113, -2, -16, -5, 12, 108, 66, -122, -90, 127, -71, 54, -33, -13, 0, -45, -64, 38, 16, 118, 108, -128, -60, 109, -128, 127, 127, -101, -86, 91, 92, 102, -128, -78, 107, -16, -5, 92, 50, -128, -128, 55, 127, -124, -74, -128, 116, 87, -128, -34, 78, 127, -128, -42, 63, -27, 1, -90, 18, -32, -119, 59, 58, 52, -117, -5, -8, -128, -128, 76, 97, -8, -128, -32, 63, 8, 127, -68, -114, -75, 70, -86, 75, 127, 73, -128, 76, -128, -119, 127, 108, -128, -108, 23, 127, 31, -128, 87, 103, -52, -106, 87, 53, -128, 127, -34, 17, 74, 0, -128, -5, -112, 107, 52, 18, -128, 59, 127, -15, -128, 73, 81, -39, -22, 26, 42, 70, 2, -114, -68, 48, 127, -45, -29, -32, 59, 127, -128, 103, -109, -122, 55, 127, -128, -88, 23, 98, 5, -128, 100, -18, -64, 68, 124, -13, -96, 127, 44, -128, 55, 53, 79, -128, -64, -53, 127, -113, -65, 87, 66, -13, -107, 127, -69, 127, -78, -11, 127, 33, -124, 27, 45, -59, -24, 93, 24, -15, -128, 6, 127, 2, -128, 127, -65, -42, 108, 36, -33, -128, 127, -71, 127, -128, 34, 127, -90, -48, 22, -1, 0, 42, 114, 127, -128, -63, 17, 116, -128, 1, 127, 116, -128, -33, 73, 81, -117, 43, -96, 127, -76, -42, 10, 127, -128, -102, 127, 34, -128, -128, 127, 127, -96, 70, -24, 96, 22, -108, -86, -80, 12, 127, 127, -128, -2, -128, 127, -123, -86, 42, 13, -16, 78, 47, -128, 6, 65, 127, 11, 73, -128, -128, 127, 92, -127, -90, 127, -29, 127, -128, 127, -68, -74, -42, 127, -127, 43, -75, 29, 127, -128, -100, 88, -128, -43, 127, 50, -128, -106, -31, 116, 116, 38, -128, -128, 106, 127, -128, -15, 109, -128, -68, 127, -45, -57, 75, -103, -1, -57, 58, -128, 54, 79, -12, -128, 5, 127, 12, 66, -21, -128, 52, 124, 48, -128, -43, 86, 65, 112, -128, 127, -39, 127, -52, 6, 92, 39, -108, -54, -93, -102, 33, 127, -58, 10, -52, 57, -128, -33, 127, 39, -128, -95, 127, 88, -128, 86, 68, -78, 33, 32, -44, 11, 127, -26, 66, 127, -43, -128, 116, 57, 36, 50, -107, 95, -38, -128, 27, 127, -71, -47, 127, -95, -128, -108, 127, -80, -128, 127, -23, -64, -113, 66, -60, 127, 117, -128, -101, 70, 127, -63, -29, -57, -128, 13, 127, 53, -2, -26, -128, 69, 69, -24, 127, -119, -7, 127, 23, -128, 55, -68, -128, 127, 42, -47, -91, 127, -52, 0, 98, 26, -10, -128, -13, -13, 127, 17, -128, -27, 91, 69, 11, -78, 79, -54, -86, 52, -26, -18, -128, 127, 127, 42, 0, -128, 118, -128, -128, 127, 100, -128, 27, 127, -87, -128, 127, 54, -128, 36, 27, 12, 127, -45, 93, -87, 127, -60, -65, -38, -43, 75, 127, -70, -75, -86, 111, 106, -45, -128, 127, 57, -2, 127, -38, -128, -85, 127, 60, -128, -27, 127, -106, -128, 127, 79, -128, 24, 127, -78, 12, 98, -128, -88, -66, 106, 127, -128, 16, -50, -128, 50, 127, 57, -128, -119, 127, -3, -128, 88, -87, 11, 127, -128, -128, 127, -107, -17, 57, -128, -55, 88, 127, -108, 6, 45, -69, 54, 15, -128, 127, 55, -55, -128, 112, 127, 91, 127, -128, -128, -17, 92, 92, 8, -128, 73, -128, 39, -87, 60, 96, -128, -43, 106, 0, -128, 21, 127, -28, -128, -73, 127, 52, -66, -23, -108, 127, 69, 38, -45, -128, 127, 127, 113, -65, -128, 127, -90, -119, 53, 102, 127, -128, -128, 127, 11, -50, -128, 127, -32, 127, 11, -128, 121, 11, -11, 98, 123, -128, -128, 55, 127, 29, -15, -79, 127, 127, -128, -128, -6, 47, 127, 22, -128, -81, -128, 127, -44, 127, 71, -65, -128, 119, 127, 71, -128, -65, 5, 57, -8, -93, 33, -28, 127, 45, 124, -54, -128, 3, 60, 101, 59, -128, -80, 71, 75, -74, -128, -8, 127, 127, -128, -103, 68, 127, 63, -128, -128, -34, 24, 119, 127, -119, 127, 119, -34, -66, 8, 114, 65, -100, -68, 97, -32, 92, 127, 15, -128, -113, 127, 53, 31, 64, -128, -96, 127, 90, -128, -21, 127, -28, -3, 95, 26, -79, 8, 100, 127, -88, -92, 31, -37, -24, -124, 50, -107, 127, -128, -3, 88, 127, -26, -128, -97, 0, 90, 127, 7, -128, 31, 119, 127, -128, -15, -128, 103, 5, 111, 24, -93, 47, 6, -103, 29, 22, -128, 23, 48, 34, -128, 63, 127, -128, -5, 127, 3, -128, 70, 5, -101, 127, -28, 32, 39, 28, -28, 23, 70, -65, 96, 127, -74, -128, 127, 60, -128, -28, 127, -113, -86, -42, -32, 71, -11, 127, -44, 127, -3, -128, -50, 108, -27, -29, 107, 127, -29, -88, -34, -38, 53, 6, 121, -17, -128, -23, 57, -116, 45, 121, -71, -128, -60, 127, 52, -127, -57, 65, 127, -22, -36, -128, 127, 26, -47, 123, -95, 11, 127, 18, -128, 8, 127, 87, 57, -66, -128, 55, -29, 127, 101, -6, -90, -128, 127, -22, 33, 85, 80, -128, 53, 43, 49, 95, -128, -109, 112, 29, 68, -75, 10, -128, 33, -8, -128, 127, 127, -48, -92, 10, -17, 32, 31, -11, 127, -112, -74, -128, 42, 127, 49, 33, -128, -36, 57, 22, -102, 29, 127, -42, -128, -119, 88, 127, 33, 88, -119, -128, -128, 127, 127, -128, -128, 23, 108, 54, -128, 121, 88, -128, 103, 15, -7, 23, -66, 65, 60, -128, 127, 92, -128, -39, 127, -128, -75, -128, 96, 127, -128, -128, 127, -103, -71, -39, 100, -23, -117, -36, 13, -117, 95, 45, -122, -45, 127, 18, -59, 121, -8, -128, 127, 17, -128, -123, 127, -34, 74, -21, 107, 3, 7, -66, -97, 2, -73, -42, 54, -128, 44, 80, 49, -43, -128, -1, 127, 15, 75, -106, -128, 52, -1, 70, -24, -97, 24, 70, 2, 127, 43, 59, -128, 100, 73, -57, -81, -2, 127, -34, 127, -78, 113, -42, 57, -70, -128, 36, 127, -121, -108, -64, 127, -128, -11, -21, 86, -128, 127, -8, 127, -128, 5, -128, 87, 70, 127, -128, -117, 127, 48, -128, 127, -116, 12, 75, -55, -128, 6, 127, -42, -128, -128, -128, 121, 127, -64, 127, -59, -128, 127, 64, -75, 13, -13, 8, -123, 34, 127, -93, -128, 127, 123, -75, 116, -1, -117, -128, 124, 127, 33, -128, 112, 33, 127, -128, 39, 123, -17, -128, -90, 58, 127, 127, -22, -128, 127, 59, -75, 24, 127, -70, -80, 127, -87, 127, -128, 32, -118, -7, 1, 127, -45, -34, 23, 101, -128, -49, -98, 127, 127, 57, -128, -23, 127, -8, -2, 91, -97, -128, -37, 127, -36, 78, 7, -128, 58, 127, 21, -118, 87, -38, 75, -50, -102, -42, 127, 108, -106, 26, 57, -128, -60, 127, -55, -16, 0, -101, 2, 17, 90, -128, -76, 127, 127, -128, -128, -44, 7, 52, 127, 75, -128, -127, 47, 127, -74, -128, -85, 0, 109, 70, 100, -121, -117, 101, -38, 23, -128, 32, -128, 28, 88, 127, -78, -128, -54, 127, -108, -128, 127, 127, -128, 127, -128, -53, 127, -128, -108, 26, -6, 37, -1, 127, -128, -128, -113, 127, -7, -43, -113, 6, 13, 50, 106, -128, -128, 28, 127, 5, -18, -128, -128, 127, 98, -28, -109, -128, 127, 98, -128, 101, 63, -66, 23, -32, 65, 109, -128, -71, -3, 26, 97, 1, 108, -36, -128, -50, 127, 86, -128, 79, -92, 90, -76, -128, 127, 38, -18, 17, -8, -64, 112, -93, 106, 88, -128, 53, -75, 103, 116, -113, -53, -55, 53, 127, -95, -128, 10, -3, 127, -128, 113, 106, -101, -11, -33, -7, 75, 127, 123, -128, -121, -37, 127, -76, -1, 39, 7, 29, -22, -50, -108, 90, 93, -128, 107, -45, 127, -128, 59, 108, -39, -52, -26, 15, -60, -43, 6, 63, 127, 52, 31, -52, -70, -10, 127, 113, -86, -128, 127, -45, -98, 57, 50, -86, 118, 33, -38, -128, 8, 127, -123, 58, 127, -103, 21, 16, -128, -69, -23, 127, 58, -128, 58, -2, 93, 52, -124, 58, 79, 80, -128, 63, 98, 27, -128, 100, -65, -128, 127, 127, -75, 11, -128, 127, -11, 8, 92, 1, -112, -128, 127, 127, -112, -128, 127, 53, -60, -26, 74, 59, 70, 127, -34, -128, 78, 127, -13, -1, -28, -85, 37, -123, 88, -128, 92, -26, -37, -26, -55, 102, -2, -103, -101, 127, 127, -52, -7, -128, 3, 127, 17, -128, -128, 127, 127, -128, 23, 109, 17, -128, 23, 127, 127, -128, -27, 106, -128, -29, -117, 127, -13, 101, -128, 127, -69, -92, 52, 127, -11, -36, -53, -128, -43, 127, 127, -128, 36, 73, -128, 48, -27, 127, 43, -32, -128, 113, -55, 123, 38, 57, -128, 127, -15, -60, -32, 38, 33, -57, 6, 11, 127, -43, 27, -44, 23, -57, -2, -128, 127, -128, -128, 29, 88, -128, 122, -48, 127, -128, 101, 127, -58, -97, 127, -24, -128, 33, 90, 127, -128, 117, 36, -101, 101, 86, -79, -121, 127, -86, -97, 127, 70, 6, -128, 91, -128, 92, -18, -76, -32, 127, -39, -114, 6, 118, 103, -42, -128, 59, 36, -49, -90, 11, 34, 127, -128, -38, -33, 91, 55, -69, 36, 26, 17, 48, -128, -79, 117, 127, -121, 3, -1, -128, 64, -27, 127, -128, -2, 127, -91, -128, 127, 127, -128, -81, 98, 127, -128, -128, 2, 127, 1, -128, 102, -80, -3, 127, 36, -59, -96, -128, 127, 127, -128, 127, 85, -128, 68, 127, -128, -92, 70, 127, -128, 54, 127, -22, -32, -48, -128, 127, 127, -128, -128, 127, 127, -101, 69, -124, 27, -5, 55, 31, 112, -128, -128, -128, 101, 127, -13, -54, -106, 127, 12, -60, -16, 48, -33, 127, 34, 32, -128, 64, 127, -128, 38, 11, -45, -60, 12, 127, 1, -128, 113, 127, -60, -128, -34, 127, 127, -107, 81, 47, -128, 6, 127, 127, -128, -128, -1, 127, 127, -128, -128, -68, 127, 127, -98, -128, -53, 0, 127, 43, -93, 93, 73, -27, 124, -45, -128, -86, 127, -114, 11, 34, -100, -128, 127, -15, -12, -128, 127, -116, 114, -57, 63, 27, 15, -128, 57, -128, 79, -18, -57, -75, 111, 127, -58, -5, -92, -74, -21, 34, -108, 127, 81, -63, -74, 127, -128, -24, 127, -79, -15, -27, -73, 8, 55, 69, 52, 2, -11, 16, 127, 127, 53, -88, -124, 127, -97, 38, -44, 50, 22, 24, 79, -31, -50, 127, -124, -128, -127, 117, 127, -128, -128, 127, -37, -11, 123, -43, -128, 108, 127, 127, -128, -49, 16, 37, -128, 114, 13, -26, -80, -116, 50, 127, 10, -128, -128, 11, 92, 97, 92, -78, 50, -128, 23, 113, -128, -2, 127, -29, -90, -18, -5, 48, 24, 13, 7, 127, -21, 127, 127, -22, -112, 45, 54, 88, 127, -128, 1, -36, -55, -95, 127, 127, -128, -121, 127, 127, -128, -60, -36, 69, -103, 113, -75, 55, 71, -42, -128, 22, 87, 15, -128, 71, 127, 96, -106, 2, -63, -128, 59, 29, -128, -13, 42, 91, 127, 37, -128, 76, 127, -13, -128, -10, -98, 127, -38, 85, 127, 37, -128, 76, 127, -118, -103, 111, 57, 79, 33, -69, -39, 127, -128, -128, 55, -26, -7, -73, 79, 127, -74, -55, -39, -90, 3, 91, -37, -76, -27, 106, -128, 69, 79, 103, -53, -76, 70, -128, -128, 116, 71, -87, -65, -6, 93, -128, -10, 96, 71, -75, 6, -73, -128, -34, 127, 127, -112, -128, -50, 127, 44, 28, 27, -59, -128, -97, 127, 24, 74, -52, 3, 53, 10, -87, -102, -118, -31, 127, 96, 59, 28, -88, -128, 60, 64, -128, 59, -52, -128, 127, -63, -22, 60, 127, -119, -66, -128, 32, 53, 90, 71, -65, 74, -128, -101, 124, 70, 0, -71, -95, -128, 127, 127, -113, -128, 58, 39, 127, -128, -128, 93, 127, -128, 63, -112, 34, -55, -37, 127, -128, 24, -128, 53, -79, -2, 108, 45, -74, 91, -128, -6, -70, 66, -128, 124, -90, 54, 127, -128, -128, 127, 87, -128, -60, -48, 122, 127, 85, -92, 93, -117, 109, -21, -87, 113, -50, -128, 80, 107, -128, 0, 127, -128, -38, -106, 121, 17, 127, -128, -76, 127, -11, -128, -34, 13, 127, 127, -112, -26, 81, -74, -44, 95, 127, 59, -128, 21, 127, 112, -128, 60, -119, -128, 127, -52, -128, 127, 24, -128, -26, 59, 127, 6, -128, -128, 127, -128, 73, 127, -43, -128, -128, 127, 98, -45, -3, -38, 69, 107, -28, -118, 74, -128, -29, -15, 101, 27, -81, 96, -128, 47, -54, 22, 43, -49, -87, 127, -107, -34, 127, 1, -128, 53, 127, -87, -128, -1, 127, -5, -11, -23, 103, 59, -90, 5, -16, 16, -128, 16, 27, 48, -48, 43, -85, 100, 2, -128, 111, 127, -78, -128, 127, 127, -92, -97, 0, 48, 127, 123, -7, -127, 122, -123, -31, -57, 39, -50, 127, 10, 65, -47, 98, 2, -50, 44, 127, -128, -73, 102, 76, -128, 44, -45, -103, 98, 6, -128, 76, 117, 74, -42, -73, 58, -12, -128, -116, 127, 42, 127, -73, -128, -128, 127, -22, 86, 17, -27, -112, 127, -86, -28, 127, -90, -128, 69, 31, 74, -37, -27, -128, 127, 127, -22, 98, -128, -6, 0, -107, 98, 47, -75, 91, -92, 78, -52, 28, -71, -111, 71, 127, -128, 96, -128, 2, -36, 127, -23, -106, -117, 111, 127, 16, -128, 52, 18, 76, 31, -124, 60, 127, 127, -107, -128, -92, 85, 127, -65, -58, 47, -122, 127, 79, -107, 71, -29, -57, 127, -124, 26, -50, 23, -13, -5, -128, 127, 28, -33, 36, -21, 71, -87, -128, -38, 127, 23, -128, -128, 127, 127, 50, -128, -123, 97, 97, -16, -86, -122, 38, 127, -128, -116, 28, 60, 102, -128, -128, -37, 127, -128, 127, -17, 68, -128, 68, 127, 55, -128, 79, 5, -128, -91, -66, 81, 127, 127, -128, -128, -44, 127, 79, -57, 122, -128, -63, 1, -55, -123, 127, 116, 7, 2, -100, 69, 26, 127, -21, -128, -1, 18, 47, 57, -101, 127, 24, 127, -57, 69, -128, 54, -96, 127, 87, -78, -91, 127, -27, -128, 127, 17, -108, 15, 127, -128, -28, -122, 69, 0, 127, -128, -15, 127, 22, -121, 121, -55, -128, -128, 86, 127, -68, -79, 127, 6, -117, -36, 127, -49, 17, 127, -16, -128, 50, 127, -128, 121, 42, 127, -117, -128, 21, 127, -74, -128, 127, 127, -128, -7, 127, -11, -7, 127, -47, -128, -128, 127, 97, -15, 0, -50, -10, 127, -86, 39, -22, -128, -128, 127, 127, -66, -128, 127, 86, -128, 117, 74, -128, -100, 127, 100, -118, 2, -26, 42, -66, 22, -44, 17, -88, -128, 81, 127, 127, -128, -128, 127, 74, -86, -108, 65, 91, -95, 127, 100, 86, -64, -78, -128, 127, 127, -111, 57, 44, -128, -3, 127, -70, -76, 23, 88, -128, 37, 127, 103, -117, -128, 64, 8, -114, 63, 127, -128, -50, -54, 108, 2, -73, -128, 127, 127, -128, -50, 53, 7, -128, 127, 13, 127, -15, -101, -39, 18, 127, -119, 53, -128, -91, 75, 16, 127, -31, -128, 119, 54, -12, 10, -63, 27, 92, -17, -128, 119, 127, -118, -127, 127, -128, -18, 64, 87, -128, -48, -57, -8, 127, 86, -13, 127, -128, -128, 114, 127, -128, -128, 127, 127, 127, -119, -128, 10, 80, 127, -7, -57, -58, 127, -54, 0, 127, 49, -63, -128, 127, 127, -111, -116, 127, 16, -55, 93, -127, -128, 86, 127, 52, -81, -106, -16, -1, -64, 106, 127, -71, -22, 127, -47, -44, 13, 26, -69, 127, 45, -22, -69, 44, 127, -128, 26, -128, -22, 23, 127, -98, -128, 74, -2, -88, 2, 17, -29, -128, 48, -128, 127, -128, 127, -119, -85, 95, 59, 107, -109, -103, -109, 39, 32, 27, 53, 64, 127, -45, -63, 39, -92, 27, -22, 87, -75, -128, 127, 88, -29, -66, -123, 127, -76, 127, 98, 127, 10, -128, -15, 71, 127, -128, -119, 36, 127, -128, -2, -7, -85, -114, -113, 71, 127, 127, -33, -98, -60, 66, -23, -128, -128, 127, 124, -71, -128, 66, 113, 43, 38, -23, -128, -47, -121, 28, 127, -86, 102, 38, -128, -128, -1, 127, 127, -128, -45, 127, -90, -111, 44, 31, 33, -117, 91, 127, -87, 107, 17, 39, -45, -64, -128, 75, 90, -49, 17, 127, -118, 5, 127, -34, -128, -128, 78, 22, 127, -42, -79, 127, -128, -79, 1, 127, -73, 16, -128, -16, 127, 95, -91, 8, -128, -26, 127, 34, -108, -128, 127, -11, 92, 127, -71, -128, 114, 7, -16, -13, 75, 18, 55, 127, -95, 75, 43, -128, 111, 24, -124, 127, -106, 108, -79, -15, -24, -11, 10, 106, -128, 43, 122, 127, -92, -128, -45, 58, -128, 75, 107, 108, -128, 45, 48, 12, -55, -109, 44, 3, 2, 48, -36, -21, 34, 127, -74, -128, -24, 1, 68, 81, 73, -87, -128, 3, 88, -85, 33, 127, 71, -95, -65, -65, 127, 98, -128, 55, 127, -10, -128, 1, 70, 48, -128, -11, -10, 127, -32, -128, -16, 113, 127, -22, 8, -97, -47, 127, -49, 33, 127, -128, 18, 33, 64, -86, 116, -34, -128, 127, -70, 88, 87, -128, -118, 127, 65, -128, -7, 127, -128, 127, -33, 118, -57, -73, 26, 127, -128, -38, 76, 17, 85, -23, -128, -91, 31, 91, 86, -27, -128, 55, -64, -128, 127, 58, -49, -128, 127, 127, -69, -128, -8, 32, -119, 127, 15, 58, 28, 85, -128, -12, 127, -93, 5, 1, -128, 111, 127, 87, -128, 21, 127, 92, -128, -128, 117, 127, -60, -128, -75, 8, 127, -27, 65, 127, -6, -76, 1, -128, -93, 127, -123, 127, 66, -128, -43, 127, 11, -124, 127, -28, 11, -128, -124, 33, 80, 90, 32, -128, 127, 127, -128, 111, 37, 127, -128, 11, 10, 127, 11, -128, 18, -34, 127, -128, -48, 127, -102, -112, 102, 127, -128, -128, 53, 127, 66, 127, -128, -128, 31, 127, -128, -49, 127, 60, 27, -128, -102, -2, 34, -90, -7, 42, 44, 107, -55, -128, 127, -31, 107, 87, 66, -98, -109, 28, 127, -123, -18, -65, 18, 127, -128, -100, 96, -52, -128, -85, 98, 127, 127, -50, -117, -37, -87, 127, 127, 3, -113, -63, 71, 127, 15, 16, 127, -68, -128, -128, 127, 15, -95, -5, 111, 28, 93, -128, -128, 48, 127, -29, -128, -128, 127, 11, -81, -8, 127, -63, -93, -128, 127, -36, -81, 127, -80, 48, 8, 34, -78, -128, 127, 127, 42, 21, -2, -21, -128, -64, 127, 103, -33, -128, -128, 121, -2, -43, -1, 127, -63, -128, 127, 85, -128, -18, 127, -55, -33, -2, -7, -96, 60, 127, 73, -39, -122, -79, 127, 121, -114, -124, 78, 127, -128, 39, 127, 88, -128, 7, 127, -76, -128, -65, 54, 127, -48, -128, 43, 127, 127, -91, -128, -96, 127, 101, -128, 18, 127, -52, -128, -54, 37, 95, 29, -39, -128, 127, 127, -118, -18, 127, 118, -128, -68, -71, 127, 103, 127, -128, -128, -21, 127, 21, -128, 42, -75, 59, 127, 15, 52, -111, -47, -37, 60, 74, 127, -22, -128, 127, 60, 59, -128, 28, 121, -8, -71, 66, -29, -102, 90, 90, -65, -102, -128, 112, -54, -6, 127, -85, -128, 60, 122, -66, -7, -55, 13, 73, -107, -7, 1, 60, 127, -12, -45, 5, 65, -71, -128, -43, 127, -32, -63, 33, -128, 5, 76, -74, -128, 24, 127, 47, -44, -91, 127, 127, 101, -117, 48, -111, 71, -44, -128, 31, -22, 114, -12, 127, -93, -128, -26, 127, 111, -39, 44, 38, 28, -128, 122, -66, -108, -17, 127, 15, -69, 57, -128, -121, 127, -64, 52, -38, 21, -48, -7, 76, -79, 127, -37, -92, 79, 127, -128, -128, 53, 127, 29, -128, -128, 81, -91, 127, 71, -21, -3, 49, -124, 92, 1, -128, 65, 127, -128, -49, 127, 90, -12, -118, -128, -109, 127, 123, -128, -128, 123, 127, -127, -116, 114, -98, 127, -39, 7, -18, 88, -49, 127, -128, -128, 71, 95, -118, -116, 127, -12, 107, -128, 118, 24, 11, 68, -128, 116, -57, 29, 93, 26, -128, -16, -53, 127, 93, -36, 65, 39, -128, -57, 122, 60, -1, -96, 16, -116, 78, 8, 38, -118, -128, 44, 127, 127, 7, -128, -66, 127, -73, -17, 23, 50, -32, -116, -50, -48, 127, 49, -54, -27, -37, -31, 127, 121, -103, -122, 0, 48, 127, -73, 127, -15, -88, -27, 127, 6, -32, -7, 33, 127, 127, -111, -39, -15, -87, -97, 57, -58, 47, -128, -76, 88, 127, -128, -128, 53, 39, 60, 23, -80, -31, 44, 32, -33, -128, 127, -33, 39, -113, 114, -86, 108, -107, 127, 5, -63, -78, 111, 117, 127, -93, -34, 88, -102, -128, 127, 127, -128, 44, 88, 37, -58, -92, 127, -128, -81, 58, 127, -12, -81, -8, -79, -128, -38, -5, 71, 95, -128, 0, 121, 12, -76, 26, -128, -11, 127, -15, -85, -128, 81, 127, -128, -44, 58, -39, 127, -128, -31, -7, 53, -2, -59, -45, -128, 116, 127, 53, -111, -90, -3, -26, 127, -70, 31, -80, -128, 127, 127, -76, -12, 100, -95, 107, 16, -29, -91, 88, 75, -113, -37, 5, 69, 127, -128, 53, 60, -52, -128, 127, 91, -128, -118, 127, 95, -31, 52, -45, -85, -12, -45, -128, 44, 96, -63, 75, 127, -119, 43, -21, 127, -97, -53, 74, -127, -111, 127, 43, -128, 113, -75, 18, 124, 6, -45, 6, 91, -128, 21, 86, -38, -128, -31, 127, -16, -90, 70, -57, -128, 21, 108, -93, -5, -96, -118, -58, 1, 127, 36, -101, 44, 127, 116, 102, -128, 121, 26, -102, 36, -49, 98, 127, -26, -128, 98, 127, 127, -128, -52, 119, 87, -114, -128, 127, 23, -66, -128, 127, 11, 127, -76, -16, -5, -128, 48, 127, 34, -128, -5, 78, -109, 93, 3, -54, -88, 96, -16, -128, 27, 127, -54, -128, -123, 121, -39, -128, 127, 97, -27, 76, 98, -128, -37, -1, 3, -10, -5, -128, -70, 70, -13, -128, 127, 18, -114, -128, 127, 55, -42, 24, 127, 127, -128, 97, -64, -55, 80, 127, -26, 44, -128, 101, -97, -128, -32, 81, 47, -114, 127, -28, 39, -31, -106, 63, -73, 78, 127, 22, -128, -103, 127, 96, -128, 63, 15, 88, 103, 79, -128, 32, -96, 11, 127, 101, -128, -74, 92, 50, -128, -93, 5, 71, 127, -127, 54, 92, -128, 109, 17, 127, -23, -63, -6, 68, -113, -53, 127, 127, -128, -100, 103, 31, -13, -54, -128, -38, -52, 111, 2, -22, 15, -79, -128, 27, 121, 117, 66, 97, -128, -128, -54, -43, 127, 90, 31, 37, -128, 55, 7, -128, 75, 127, 127, -117, -128, 127, 127, -87, -13, -85, 0, 53, 114, -102, -128, 127, 127, -128, -88, 127, 16, 127, -52, -122, 93, 45, 70, 80, -128, 54, 79, -128, 127, 31, -45, -103, 127, 127, -106, 69, -64, -5, -128, 127, 127, -64, -128, 127, 124, -74, 127, -18, -128, -53, 127, 98, -38, -108, 37, 81, -128, 106, 101, -11, -128, 47, 127, -128, -39, 127, 22, -38, -128, -7, 127, 127, -123, -128, -112, 127, 127, -1, -128, -64, 127, -44, 33, -91, -45, -128, 48, 112, 116, 37, -97, -128, 127, -128, -49, 6, 127, -18, -116, -128, 127, 6, -127, 6, 113, -55, 70, 127, 92, -128, 37, -76, -127, 122, -42, 2, 118, -42, -66, -128, 127, -32, 127, -59, 92, -57, -128, -52, 127, 113, 16, 107, -31, -128, 127, 127, -26, -78, 88, 8, 127, -12, 90, 36, 24, -80, 127, 116, -128, 66, -113, 122, 127, 43, -7, -128, -128, 80, 127, 95, -128, -50, 107, -128, -128, -121, 127, 127, -127, -128, 80, 127, 0, -90, -128, -31, 55, -60, 85, -39, 114, 127, -58, -112, 42, 12, 32, 127, 28, -54, 50, -128, 127, 88, -5, 107, 3, -128, -128, 127, 39, -100, -128, 127, 106, -73, 127, -13, 1, 78, 91, -79, -128, -128, 127, 127, -128, -55, 127, 127, -128, -121, 91, -8, -128, 81, 127, 63, 8, -128, 39, 66, -128, 80, 5, -91, -98, 127, 12, 47, 28, -50, -128, -71, 50, 116, -11, -128, 0, 127, -39, -39, -123, 75, -6, 2, -116, 95, 127, 127, -100, -128, 0, 127, 127, -128, -23, -44, -42, 64, 43, -22, 127, 0, -58, -114, 26, 58, -45, -128, -18, 92, 124, -63, -64, -59, 95, -128, -128, -10, 127, 81, -128, -7, -15, 36, 17, 127, -128, -18, 127, -43, -128, 7, -29, 116, 16, -128, 85, 29, 124, -2, -44, 23, -87, -27, 127, 53, -91, -90, 45, 6, 80, -54, 32, -57, -13, -128, -128, 65, 127, -59, -128, 127, 117, -128, 0, 119, -57, -55, 16, 127, -74, -128, -93, 127, -87, 112, -128, 57, -26, 127, -128, -53, -128, 127, 42, -52, -128, 88, 127, 127, -128, -18, -76, 127, -97, 121, -128, 127, 0, -128, 17, 127, 29, -128, -58, 127, -128, 127, -76, 36, -121, 79, -54, 87, 58, -66, -28, 80, 76, -11, -128, -91, 127, -1, -128, -10, 127, -6, -128, 2, -13, 47, 127, 29, -128, 31, -22, 127, -50, -121, -54, 127, 127, -128, -65, -128, -3, 127, -78, -34, 27, 15, -128, -13, 97, -26, -73, 114, 0, -69, -128, 88, 49, 127, -47, 63, 17, -128, 111, -75, -128, 39, 127, 76, -128, 58, -70, -57, -60, 127, -27, -93, -123, 11, -128, 127, 98, 127, -122, -10, -66, -28, -101, 58, 127, 68, -21, 127, -128, -118, -78, 127, -128, 17, 42, 36, -128, 22, 127, -68, -39, 127, 26, -18, -128, -93, 127, 28, 57, -116, -128, 124, -23, 107, -128, -18, 127, -128, -128, 24, 1, -91, -8, 127, -45, 108, 42, -122, -21, 28, 127, -128, 58, 15, 8, -128, 127, -37, 74, -73, 3, 112, 78, 98, -73, -128, -2, 96, -128, 127, 31, -66, -52, 127, 32, -128, -73, 2, 97, 127, -36, -36, 127, -29, -128, -7, 66, 38, 26, -7, -80, -65, 28, 127, 127, -116, -128, 11, -70, 65, 70, -45, -74, 1, -88, 127, 34, 32, 127, -22, -128, 127, 127, -128, 74, 75, 95, -128, 52, 127, 22, -128, -100, 28, 111, 127, -121, -128, 102, 78, 42, -27, -65, 127, 118, -37, -128, 74, 127, -91, 24, 127, -65, -128, 58, -128, 127, 57, -96, -106, 93, 127, -128, -79, -5, 118, -128, 17, 127, 127, -114, -64, -87, 127, -31, -128, 0, 15, -45, 127, -26, -74, 11, 109, 92, -128, -42, 52, 21, -8, 2, -128, 38, 127, 127, 116, -128, -128, 63, 127, 32, -128, -128, -37, 127, 127, -128, 36, -128, 127, 3, -39, -22, 102, -128, 127, -38, 64, 86, -128, -128, 127, 127, -88, -128, 127, 112, -128, -29, 127, -113, 37, 127, -11, -128, -128, -23, 127, 127, -119, -97, 17, 50, -36, -128, -28, 127, -87, -3, 23, 5, 33, 127, -128, -128, 127, 23, 68, -113, -101, 127, 127, 10, -128, 127, -128, -31, 18, 95, 16, -128, 27, 127, -59, 127, -63, -128, 102, 127, -33, -123, 1, 78, 29, -128, -66, -45, 23, 127, 33, -128, -24, 127, -5, -121, -128, 127, 127, -18, -128, -128, 114, 127, 127, -128, 49, -73, 127, -78, -12, -74, 93, -29, 91, 127, -128, -71, -47, 80, 86, -68, -85, -48, 119, 38, -128, -33, 64, 92, -128, 127, 122, -128, -7, 127, -108, -31, -128, 69, 119, 6, -111, 54, -6, -60, -87, 127, -81, -128, 127, 95, -111, 23, -23, 127, 5, -2, -103, 117, -12, 124, 7, 76, 127, -128, 15, -38, -128, -6, 32, 127, -42, -26, -26, 73, 127, 60, -128, -107, 10, 127, -97, -3, 93, 60, -47, -128, -95, 22, 127, 76, -128, -108, 127, 1, -128, 127, 23, -112, 95, 76, -70, 127, -81, -88, 3, -128, 31, 127, -93, -23, -128, -69, 127, -128, -88, 73, 127, -121, -128, 53, 38, 112, 18, -128, 7, 127, 64, -128, -50, -90, 102, -32, 37, 127, -54, -128, 121, -79, 79, 75, -33, -128, 78, 127, -114, -21, 112, 127, -128, -128, 50, 2, 32, -11, -93, 78, -128, -42, 12, -39, -128, 127, -28, 66, 24, -5, -128, 108, 87, 98, -128, -98, 33, 85, -128, 8, 127, -58, -128, 12, 127, -68, -128, 127, 80, -52, -74, -39, 5, 127, 100, -33, 15, -118, -100, 127, 50, 3, 13, -54, -128, 31, 127, 127, -53, -128, 93, 10, -128, -70, 116, 24, 65, 31, -6, -128, 28, 127, 54, -128, 93, 50, -128, 50, 116, 44, -128, -8, 127, 1, -128, -7, 127, 32, 28, -97, -29, 127, 31, -102, 32, 85, 59, 101, -96, -128, 80, 27, -1, 58, -100, -128, 117, -34, -31, 57, 1, -70, -128, -39, 127, 127, -128, -122, 127, 0, -103, -128, 127, 3, -128, 3, 127, 13, -122, -128, 127, 50, -11, -118, 12, 60, 100, 31, 33, -128, -96, -128, 127, 74, -91, -128, 58, 127, 60, 16, 39, -128, 29, -27, 100, 7, -128, 95, 127, 28, -101, -2, -1, -109, 2, 49, -128, 95, -117, 122, -86, 71, 69, -76, -128, 127, 3, 70, -44, -55, 127, -128, -12, -78, 114, -79, -10, 73, -97, 127, -58, -128, 127, 10, -128, 95, 127, -128, -128, 12, 127, -102, 123, -128, -11, -118, -47, 127, -92, -18, 101, -90, 78, -97, -28, 106, -36, 2, 57, -11, 16, -8, -88, -38, 87, -12, -128, -3, 127, -23, -128, -66, 86, 10, 118, 85, 66, -128, -8, 127, -54, -128, 26, 127, -128, -37, 39, 127, -128, 10, 103, -71, -44, 59, -109, 127, 18, -128, -18, 127, -128, 127, -34, -73, -3, 127, -128, -88, 112, 101, -128, 118, 90, -100, -80, -44, 127, 127, -128, 7, -2, 108, -128, 127, 11, -3, -98, 79, 127, 10, -128, 127, -29, 23, 127, -86, -128, 127, -128, 71, -22, 45, -128, 70, -12, 127, -121, 34, -68, 31, -49, 54, -65, -128, 107, 127, -55, -128, 53, 71, 127, -79, -47, -109, 127, -31, -128, 127, 5, -128, -33, 127, -18, -75, 39, -96, 127, -23, 3, -128, -45, 127, -12, -128, 15, 116, 0, 42, 93, -128, 114, 31, -128, 127, 127, -128, -45, 68, 117, 127, -95, -128, 11, 127, -12, -128, 71, 33, -118, -70, 127, 75, -128, -102, 127, 8, 73, -128, 70, -65, -29, -113, 127, 17, 10, 64, -48, 127, -70, -18, 85, 68, -80, -128, 88, 127, -68, -50, -128, 127, 12, 127, -128, 1, -128, -3, 81, 127, -47, -92, 15, -63, -128, 74, 124, 2, 8, -24, 24, -55, -128, -128, 127, 70, 127, -55, -49, -128, 92, 127, -1, -128, 127, 48, -15, -27, 34, -128, 127, -38, 93, 1, -64, -7, 88, -29, 0, 103, -15, -128, 127, 127, 39, -58, -53, -34, 33, -3, -111, 47, -6, 97, 28, 113, -81, 11, 2, -96, -128, -96, 28, 127, 21, -128, 127, 127, -128, -87, 127, -128, -36, 127, 3, -81, 10, -128, -92, 127, 109, -102, -109, 75, 27, -49, 45, 57, -66, -128, 65, 93, 127, -54, -5, -31, 7, -68, 53, 8, -45, -36, -65, -3, 29, 34, -59, 127, 65, 21, -71, -128, 49, -26, 95, 103, -128, -26, 127, -5, -128, 127, 90, 5, -128, 119, 10, 127, -58, 12, -128, 127, 81, -128, -7, 127, -68, 7, 127, 116, -128, -128, 127, 127, -79, -98, 127, 127, -128, -128, 97, 127, 5, -59, 127, -112, -128, -128, 127, 127, -55, -128, 69, -21, 127, 27, -96, 38, 116, 43, -85, 32, -128, -3, 127, -128, -15, -15, 93, 3, -121, -128, 127, 127, 127, -128, -128, 122, 38, 47, -128, -128, 127, 0, 66, -86, 80, -128, -24, 127, -54, -128, 93, -128, 49, 127, -16, -128, 23, 127, -5, -117, 57, -128, 86, 107, -113, 66, -8, -28, -128, 38, 127, 73, 55, -44, -128, 116, -128, 17, 68, 13, -87, -118, 119, 113, 68, 91, -54, -59, 48, -12, -128, -128, 127, -95, 13, 116, -63, -128, 1, 127, 127, -112, 31, 71, -76, 127, -102, -128, 95, 127, -128, -65, 127, -21, -85, 65, 127, -63, -86, -128, 107, 127, 127, 112, -128, -128, -48, 103, -1, -128, 69, 127, -12, -128, 45, 127, -31, -128, 106, 118, 53, 75, -128, -121, -2, 127, 49, -128, 88, -12, 127, 127, -128, -73, 127, -24, -97, 43, 127, -98, -128, 127, -68, -92, 100, 88, -70, -128, -6, 127, -48, -24, -128, -52, 90, 50, 66, -116, 79, -128, -128, 127, 0, -79, 50, 42, 85, -49, -128, 47, 127, 127, -101, -128, -95, 106, -45, 97, 127, 127, -76, -128, 93, 1, 76, -66, -33, 127, -114, -32, -128, 111, 47, -63, 55, 22, 45, -128, -21, 127, -28, -76, 81, -37, -23, 98, -3, -52, 127, 0, -103, -15, 100, -33, -34, 127, -69, -127, 127, -47, -123, -118, 127, 42, -49, -75, -60, 107, 127, 44, -128, -12, 127, -128, 58, 73, -128, 101, 109, -65, -23, 6, 15, -31, 127, 112, 119, -88, -128, -128, 127, 76, -128, 28, 127, 13, -55, -49, 78, -119, -128, 12, 88, -76, 33, -32, 127, -78, -128, 95, -24, 124, -75, -128, -63, 93, 16, 127, 13, -128, -128, 127, -26, -55, -71, 127, -87, -128, -3, 127, -128, 7, -64, -128, 63, 127, -26, 5, 95, -128, -128, 122, 127, -128, -128, 127, -38, 21, -55, 127, -87, -128, 48, 43, 112, 59, -22, -128, 127, 39, 65, -128, 127, 75, -95, -128, 127, 127, -128, -93, -98, 127, 52, -128, 121, 127, 44, -128, 116, -87, 127, -66, -112, 66, 55, -128, 69, 127, 22, -96, 15, 57, -15, -87, 47, 127, -128, -21, -43, 68, 45, 52, -108, -128, -42, 127, 1, -36, 0, 127, -64, -49, 18, 79, -87, -128, 127, -42, 38, -39, -86, 23, 127, -93, 88, -31, 127, -128, 127, -98, -60, 22, 127, -128, 2, 21, -128, 18, 121, -7, 71, -128, 3, -5, 57, -95, 55, -16, 55, 0, -128, -11, -128, 36, 68, 127, -66, -128, -128, 127, 127, 127, -128, -39, -128, 127, 54, -64, 52, 45, -128, -50, 101, 127, -87, -24, 127, -93, -64, 54, 48, 66, -38, -39, -128, 127, 17, 127, -86, -128, -48, 127, 8, 127, -128, 17, -128, 127, -64, -128, 127, 95, -128, -74, 127, 31, -128, -85, 127, -24, -128, 38, 127, 38, -128, 44, -52, -3, -128, 121, 93, -54, 0, 81, -11, -91, 102, 54, -128, -57, -5, 127, -38, -44, -33, 103, -95, -123, 16, 7, 127, 92, -128, 127, -97, 64, 38, 127, -37, -128, -128, 15, 127, 58, -128, -18, 88, -101, 68, 127, 127, -57, -128, 93, 81, -121, -44, 31, -26, 127, 116, -58, -128, 55, -23, 111, -7, 69, 127, -128, -119, 29, 127, -128, 58, -128, -32, 58, 58, 75, -100, -128, 127, -36, 24, 32, 127, -69, -128, -18, 50, 93, 127, -96, 15, -128, 44, 53, 37, -128, 127, 127, -34, -98, -128, 127, 50, -87, 53, 31, 92, -128, -42, 117, 70, -128, -128, 127, 66, -128, -97, 127, 127, -86, -63, 58, -128, 127, -111, 114, -31, -33, 65, -26, 12, 55, 32, -128, 116, 127, -6, -128, -53, 7, 93, 127, 10, -128, -16, 12, 27, 81, 127, 31, 59, -128, -90, 127, 91, -114, -107, 32, 31, -113, -68, -128, 127, 127, -87, 5, -81, 47, 127, -128, -17, 106, 38, -128, -128, 127, 107, -47, 43, -45, 75, -73, 100, 48, -128, -29, 117, 33, -3, -128, 127, 96, 45, -64, -12, -128, 69, 127, -3, -78, 38, -50, 6, -128, 1, 76, -101, -79, 50, 127, -128, -69, 127, 12, -128, -5, 127, 11, 122, -128, 3, 127, -128, -53, 127, -80, -123, 127, 0, -128, -24, 127, 127, -128, -128, -15, 97, 127, -128, 6, -92, -118, 96, 113, -128, -13, 112, 22, 29, -85, -102, 54, 55, -54, -128, 1, -107, 127, 127, -65, -128, 10, 127, 127, -85, -128, -48, 60, 38, -75, -128, 127, -100, 80, 80, -60, -128, 127, 33, 76, -23, -59, 45, -43, -15, -23, -128, 58, -122, 81, -21, -128, -50, 127, 26, -128, -23, 127, 16, 106, -128, 15, 127, -13, -23, -128, 16, -42, 73, -128, 71, 127, 44, -128, 6, 127, 127, -128, -128, 127, -69, -3, -128, -37, 31, 119, 1, -128, 0, 127, -75, -128, 21, 127, 109, -128, -11, 127, -128, -108, 103, -128, -68, 58, 127, -91, 127, -123, -128, -128, 127, 44, -55, 127, 93, -75, 24, -128, -64, 127, -7, -15, -121, 100, 78, 127, -128, -128, 2, 108, 47, -31, -31, 38, -102, 127, 127, -128, 13, -79, 127, 2, 2, 57, -26, -128, -128, 127, -121, -128, 127, 101, -128, 21, 127, -85, -95, 44, -31, -128, 34, 92, -98, -53, 127, -128, -128, -6, -73, 127, 43, -7, 38, 127, -31, -128, 127, -23, 0, 3, 108, -34, -38, 15, -50, 127, -128, -128, 70, 36, -36, 127, -128, -128, 7, 127, -106, 49, 53, -128, 31, 6, 57, -79, -106, 107, 121, 127, -102, -128, -128, 109, 69, 127, -93, -128, -48, 127, 127, -128, -16, 71, -128, 15, -10, 3, -128, 68, 74, 127, -7, 2, -128, -98, 127, 78, -128, -74, 27, 113, 10, 95, -128, -102, 127, -26, -66, 60, -53, -128, 127, 1, -91, 57, 127, -128, -128, 127, 113, -113, 107, 52, -128, -116, 127, -27, 47, 127, -128, -114, -66, -37, 107, 127, 127, -102, -128, -128, 127, 80, -128, 127, 37, -36, 88, -78, -52, 127, 75, -128, -128, 127, 16, 60, 22, 127, -24, 15, -128, 96, 127, -128, -2, 70, 74, 86, -128, -128, 42, 117, -49, -74, -128, 127, 111, 24, -59, -63, 97, -124, -124, 127, 68, -128, -18, 127, 127, 102, -128, -23, 27, 8, -23, 18, -90, -79, -47, 117, 127, -108, 71, -128, -16, 71, 49, -128, -96, 127, 1, -109, 127, 80, -128, -87, 8, 76, 127, -97, -13, 91, 0, -128, 65, 80, -121, 107, 127, 7, -33, -70, -116, 127, -75, 78, 26, -128, 13, 127, -86, -100, 24, 127, -86, -11, 127, 22, -128, -80, -49, 127, 127, -109, 43, 12, 37, -70, -34, -7, -33, 127, 127, -74, -128, -32, 37, 79, 95, -70, 26, -128, 127, -31, -128, 127, 48, 127, -52, -128, -28, 127, 75, -7, -128, -73, 127, 127, 1, -63, -128, 90, -128, -1, 127, 103, -93, -53, 118, -128, -128, 101, 102, 57, -128, -85, -128, 127, 13, 11, -68, 90, -80, 60, 28, 36, 127, -128, -29, 69, 23, -69, 0, 0, 55, -71, 127, -53, -21, 127, 127, -128, -63, -102, 127, -43, 90, -12, -128, 127, 127, -47, 42, -128, 73, -33, 127, -128, -32, 114, 121, -34, -28, -128, -73, 57, -16, 54, -65, 55, -58, -128, -107, 69, -17, 102, 74, -69, -45, -113, 122, 127, -128, -48, -5, -49, -47, -24, 127, 124, 97, -128, -128, 93, 127, 76, -128, 18, -128, -21, -39, 100, 71, 127, -128, -128, 28, 122, -128, 127, 100, 66, -128, 7, 121, 116, -128, -57, 123, 33, -128, 100, 73, -128, 101, 93, 49, -128, -23, 2, 11, 60, -15, 69, -81, 38, -18, -127, -128, 108, 127, -111, -91, -54, -33, 16, 127, -64, 52, -128, 85, 100, -54, 68, -78, -42, -128, 103, 127, 13, -128, 119, 114, -128, -15, -49, 42, 70, 127, -128, -101, 22, -11, -37, 43, -91, 54, -1, -88, 96, 102, -97, -128, 73, 107, 7, -128, 34, 127, -8, -128, -49, 127, -63, 64, -69, 13, -128, 74, 127, -128, -12, 127, 64, -128, 11, 109, -92, 90, 127, -128, -10, 100, -47, -26, 12, 127, -88, 7, 127, 16, -128, 127, 55, -64, -28, 124, 87, 43, -5, -128, -66, 38, 8, -128, 127, -128, -29, -128, 87, -11, 127, -28, -59, -87, 127, 127, -102, -113, -63, 96, 87, 127, -128, -10, 85, -128, -12, 127, 127, -92, -128, -128, 127, -107, 127, 31, -128, 18, 127, -128, 127, -78, 70, -49, -95, 127, -37, -34, 52, 74, 13, -23, -128, -47, 127, -128, 18, -18, 36, 57, -128, -60, 107, 127, -109, -54, 92, -128, -55, 22, -13, -42, 91, -74, 127, -12, 22, 118, 127, -128, -128, 15, 127, -8, -128, -114, -26, 127, 17, 113, 70, -114, 127, 17, 127, -65, -127, 127, 121, -128, -128, 127, 69, 22, 34, -55, -28, 18, -24, -44, 44, -128, 49, 75, -86, 3, 117, 127, -128, -128, 127, -50, 48, 17, -57, 53, 34, 127, -128, -128, 27, 127, -16, -128, 90, -106, 127, 60, -2, -112, -29, 92, -31, -98, 127, 88, 69, -65, -121, -29, 22, 18, 16, 127, -3, -17, 124, 15, 6, 80, -28, -128, -10, 34, -43, -114, -8, -128, -103, 127, -34, -119, 8, 127, -5, -32, -103, 73, 127, -102, -63, -24, -7, 49, -128, -128, 127, 78, -88, -32, -27, -128, 127, 127, -128, -54, 127, 88, -128, -33, 111, -128, 31, 53, -108, 13, 24, 127, -128, -57, 127, 7, -122, -64, 127, 0, -91, 54, 42, -52, -85, 127, 59, -114, -102, 69, 127, 127, -128, -31, 49, 118, 5, -128, 34, 29, -57, -91, 127, -28, -81, -128, 101, 93, -47, 127, 96, -128, 70, 127, -107, -60, 81, -13, -32, -50, 76, 15, 70, 127, -118, -128, -128, 124, 127, -70, -50, 127, -92, -55, -13, 70, 16, 23, 95, 39, -97, -80, -128, -57, 45, 127, 103, 121, -128, -128, 7, 127, 93, -118, -80, 6, -5, 127, 127, -123, -108, 5, 95, -92, 127, -73, -74, -87, 97, 76, -8, 102, 38, -74, -73, 127, 55, 12, 3, 5, 45, 127, -100, -128, -37, 107, 10, 127, -128, -74, 76, -106, 49, -71, -69, -21, 2, 98, -128, 8, -90, -44, -33, 36, 55, 127, -54, -95, -128, 124, 91, 127, -36, -128, 63, 16, -66, 32, 127, 10, -128, 58, 54, -128, 92, 33, 74, 52, 6, -42, 73, -1, -45, 6, -88, -128, -8, 127, 127, -128, -60, 2, 117, 18, 22, -68, -58, -59, 127, 127, -44, -16, 50, 127, -128, 76, -15, -128, -74, 127, 127, -3, -49, 127, -119, 6, 127, -16, -128, 70, 127, -81, -70, -128, 127, -22, 93, 10, -128, -15, 127, 109, -44, -128, -87, -86, 127, -70, -2, -124, 127, -37, 1, 44, -88, -34, -16, -100, 6, 47, -128, -32, -1, 32, -64, 112, -127, -85, 60, -10, -128, 3, 127, 36, -95, -128, 39, 127, -114, -111, 69, -2, 127, -101, -57, 18, 127, -128, -128, 3, -69, 107, 107, 127, -128, -128, 127, -68, -122, 127, 58, 24, -128, 31, 64, -13, -127, -76, 44, 112, -100, 92, -11, 0, -36, -92, -96, 127, -24, -26, 27, -39, 116, -128, -128, 127, 18, -128, 68, 127, -15, -128, 127, 123, 93, -74, -90, 127, -128, -27, 57, 31, -128, -47, 127, -128, -71, -37, 3, 50, -13, -10, 127, 65, 0, -128, 70, 127, -107, -53, 127, -128, 36, 127, 88, 90, -128, -31, -39, -95, 119, 59, 18, 47, -45, -128, 42, 37, 96, 127, -128, -90, 88, -49, -111, 119, 50, -70, 16, 127, -100, 12, 127, -66, 47, 97, -31, -81, 127, -97, -68, 113, -128, 58, 127, -44, -85, -63, 63, 127, -101, -42, 97, 102, -128, 127, 52, -5, -58, 97, -2, -128, 119, 45, 78, 31, -3, -128, -16, -26, -12, 34, -128, -26, 127, -68, -68, 97, -128, 93, 127, -107, -128, -36, 127, 64, -22, -26, 21, -98, 38, -91, -34, 8, -75, -128, 106, 127, 108, -118, -112, 15, 12, 0, -128, 13, -91, 118, 80, -52, -93, 32, 127, -128, 15, -5, -128, -16, 106, 127, -92, -128, -74, 38, 127, -2, 55, -60, 127, -107, -98, 127, -128, 68, 13, -128, -116, 127, -31, 68, 27, -75, -55, 127, 124, -128, -52, 7, 127, -128, 118, -58, -22, -128, 127, 127, -39, -128, 127, 127, 50, -128, -2, 16, 90, -63, 43, 96, -48, 57, 17, -32, 127, 22, 1, 26, -58, -95, -42, 127, 122, -21, -128, -103, 76, 127, -128, -93, -48, -121, 127, 127, 27, -128, 59, -31, 8, -11, -128, 15, 127, -66, -128, 78, 127, -22, -50, 127, 107, -128, 28, -32, -59, 96, -91, 127, -23, -34, 75, 117, -128, -128, 16, 114, 6, 69, -92, 15, 127, 53, -128, 66, 127, -111, -121, -128, 127, 95, 45, -128, 43, 24, -75, 68, 127, -128, -38, -81, 34, 127, -107, -80, -91, -58, -50, 127, -6, 6, 111, -128, -49, 69, -2, 59, -33, 127, -66, -128, 109, 92, -122, 12, 98, 42, -128, 32, 117, 127, -74, -128, 31, -128, 10, 112, -12, -2, 57, -128, 116, 0, -128, 38, -65, 127, 93, -128, -79, 127, -15, 108, -21, -22, -97, -37, 127, 37, -53, 22, 127, -11, -118, -128, -44, 76, 63, 66, -53, 39, -128, 43, -26, 75, 93, 23, -128, -16, 127, 54, -123, 127, 8, 92, -29, -75, 42, -23, 127, -57, 34, 73, 50, -64, -107, -54, -75, 127, 1, 127, -47, -80, 26, 127, -85, 23, -79, -112, 43, 34, -2, -80, 114, 127, 106, -116, -15, -128, 127, -73, 16, 127, 28, -76, -113, 65, -128, 127, -91, 127, -17, -128, -11, 127, 127, -128, -128, -36, 27, 58, -88, 49, 127, -128, -128, 71, 33, 15, 43, -81, -128, 53, 127, -128, -102, 127, -29, -128, 33, -63, 127, 1, 109, -108, 73, 127, 8, -128, 114, 22, 48, 127, -107, -38, 7, 31, -97, 127, -128, -128, -50, 127, -26, 11, 127, -128, -128, 127, 106, -128, -124, 127, -24, -117, 88, 6, -128, 127, -68, -91, -86, -128, 127, 127, 91, -81, -128, -16, 3, 44, -15, -128, 0, 75, -128, -87, 127, -128, -42, 127, -78, -114, -45, 15, 5, 127, -97, -128, 127, 109, -102, 66, -49, -1, 55, -128, 26, 112, 127, 37, -31, -128, 44, 81, -128, 28, 32, 127, -128, 15, -76, -103, -44, 127, 48, -128, -128, 109, 127, -36, -93, -128, 109, 5, 80, 59, 32, -107, -93, -92, -22, 127, 39, -128, 90, -6, -64, 127, -45, -128, -1, -8, 127, 16, 42, -39, -13, -34, 127, 10, -54, -128, 127, 127, 18, -128, -90, -11, 36, 127, 127, -117, -128, 123, 127, -23, -128, -11, 127, 127, -118, -128, -121, 127, 127, 45, -128, -91, 127, -48, 50, 79, -53, -128, 90, 127, -128, 52, 42, 64, 127, -57, -128, -128, 127, -98, 127, -109, 7, -97, 127, -12, 28, -128, 68, -98, 24, -45, -44, 127, 54, -128, -11, 127, -27, -128, -24, 96, 127, -43, -114, 28, -49, 71, -10, 92, 15, 6, -128, 18, 31, 101, 43, 80, -95, 15, 127, -128, 17, 43, -29, -47, 121, 81, -22, 44, 86, 106, -128, -96, -128, 108, 127, 85, -47, -128, -11, -48, 127, 44, -128, 80, -37, 53, -60, -128, 79, 73, -78, -39, 68, 123, -48, 17, 121, 17, -128, 127, 127, -128, 34, 45, 96, 43, -128, -97, 127, 87, -23, -128, -2, 108, 12, -26, -10, 123, 127, 127, -128, -128, 8, 127, -128, -3, 76, -37, -43, 69, -81, 92, 91, -128, 47, 127, -92, -80, 78, 47, -128, 127, -11, -80, 44, -54, 57, 127, 0, -128, 31, 79, 43, -128, 127, 86, -128, -81, 127, -106, 127, 21, 6, 21, -78, -26, -22, -23, 127, -26, -117, 127, 8, -45, -121, 88, 90, -107, 0, 36, -66, 127, -5, 27, 48, 76, -91, 48, -16, -128, 10, 127, 91, -96, -50, 93, 48, -50, -101, -59, -85, 71, 29, 88, 127, 127, -128, -128, -109, 127, 107, 127, -2, -128, -52, 23, 127, -95, -119, 0, 53, -128, 64, -42, -118, -95, -36, 127, 127, 64, -118, 28, -128, 7, 127, 127, -128, -128, 44, 127, -100, 39, -31, -1, 24, -37, -128, 23, 127, 127, 66, -128, -128, 6, -33, 127, -15, 107, -54, 127, -128, -28, 127, -12, -119, 66, -128, -79, 127, -88, -119, -26, 113, 6, -85, 123, -34, -17, 127, -97, -128, -114, 127, -79, 121, 107, -42, -128, 73, 127, 37, 34, -128, -93, -63, 127, 37, -118, 26, 127, -85, 85, -128, -60, 127, -32, -128, 11, -88, 95, 60, 127, -128, 57, -128, 116, -3, -57, -13, -2, -128, 127, 127, 127, -45, -128, -50, -3, -93, 49, 127, -93, -128, 22, 54, 11, -81, 55, 119, 64, 24, -128, -100, 33, 45, 48, 11, -128, -128, 44, -90, 78, 127, -3, -93, 127, -128, 34, -64, 66, -39, 60, -18, -128, 127, 60, 127, -128, 0, 108, -11, -29, -109, -64, 127, -108, -21, -32, -21, 127, 44, -128, -48, 127, 6, -16, -112, 24, 2, -73, 28, -113, 92, -66, 22, 108, 127, -128, 101, 7, -69, 42, -74, 38, 127, 73, -128, -128, 127, 21, 112, -128, 59, 117, -50, -92, -5, 107, 76, -128, 73, 54, -128, -119, 127, -102, 53, 23, -48, -128, 127, -114, -73, 127, -37, -128, 127, 47, -128, 24, 127, -27, -33, 100, 53, -65, -128, -121, 127, -45, -107, 127, 109, -128, -128, 127, 37, -128, -102, 127, 27, -128, 42, 59, 24, -128, 55, 127, -10, -128, 112, -128, -128, 102, 127, -128, 11, 112, 86, 26, -128, -100, 78, 12, 45, -3, -128, -128, -39, 127, 127, -128, -128, 127, 28, 11, 26, -128, 26, 127, 127, -128, -66, 127, -34, 23, -128, -65, 102, -26, 27, -11, 31, -128, 127, 63, -128, -71, 127, 114, 116, -47, -128, -128, 50, 127, -32, -128, -54, 127, -23, -63, 22, 101, -79, -55, 49, 0, 127, 127, -101, -128, 70, 127, -43, -70, -42, -116, 127, 127, -111, -128, 102, 32, 86, -128, -78, -11, 71, 33, -65, 33, -128, -53, -127, 96, 17, 114, -43, -5, 52, -36, 127, -128, -118, 95, 127, -128, 16, -10, -26, -66, 68, -21, 93, 127, -128, -13, 12, 127, -128, -128, -22, 69, 23, 107, -26, 21, -66, -17, 68, 127, -128, -128, 100, 21, -128, -60, 127, -127, -5, 127, -96, 16, 121, -128, -76, 127, 127, -128, 48, -28, 88, -123, 127, -7, -128, 17, 27, -18, 127, 127, -36, -103, -128, 127, 0, -128, -71, 127, 7, -55, -128, -102, 127, -1, -13, -52, 127, -73, -128, -97, -95, 127, 127, 47, 98, -47, -128, -57, 101, 80, -49, 0, -39, -6, 122, -123, 24, 127, 127, -128, -128, 31, 119, 48, -121, -58, 71, -54, -95, 127, -102, 27, 18, -128, 2, 127, -11, -128, -97, 29, 127, -79, 122, -43, 3, -54, -87, -85, 127, 37, 68, 127, -128, -128, 1, 127, -50, 71, -128, -52, -123, 60, 107, 127, -128, -128, 88, 127, -114, 45, -128, -43, 127, -78, -128, -21, -91, 118, 16, 24, -112, -43, 27, 127, 22, -95, -26, 108, 96, -128, -128, 68, 127, -128, -80, 85, -59, -70, 127, 6, -107, -69, 42, 6, -48, -80, -128, 90, 34, 33, -28, -128, -38, 127, 59, -128, -24, -79, 44, 127, 2, 49, -128, -121, 27, 127, -107, 49, -3, -39, -75, 102, -128, 88, 6, -92, -111, 55, 39, -8, 33, 127, -102, 71, 127, -17, -128, 58, -21, 127, -128, -106, 3, 106, -26, -121, -66, 127, 59, 127, -128, -47, 92, -45, 16, -101, -88, 86, 66, -86, -6, 71, -128, -112, -23, -18, 75, -76, 127, 127, -128, -47, 127, 64, -65, 17, -128, 33, -65, 52, -128, 127, -101, 80, -10, 127, -26, -128, -6, 69, -128, 127, 127, -128, -75, 124, -13, 33, 7, -1, -60, -128, 38, 0, -88, -96, 127, 37, 23, -128, -48, 127, -80, -128, 127, -95, -79, 112, 127, -101, -128, 127, -47, -17, -128, 81, 127, -21, -128, -92, 127, -128, -5, -24, 68, -128, 127, -52, 58, -128, -12, 103, 127, -102, -74, 27, 52, -34, -26, 127, 101, -128, -29, 73, 127, -98, -128, 93, -48, 55, 127, -53, -128, -79, 127, 60, 88, -95, 29, 127, -47, -128, 24, 103, 31, -128, 75, 127, -29, 43, -68, -128, 127, -98, 6, 23, -55, -128, 111, 127, 39, -128, 90, 127, -128, -15, 16, 127, -60, -128, 11, -75, 127, 59, 127, -128, -1, 127, -128, -16, 96, 24, -93, -111, 0, 127, 6, 118, -16, 22, 8, -28, 45, -8, -103, 127, -3, -128, 114, 127, -128, 59, -49, -55, -15, 127, 5, -64, -39, -106, 127, 10, -128, 127, 81, -128, 81, -8, -92, -2, 127, 39, -128, -5, 127, 5, 127, -36, -73, -5, 17, -47, -42, -70, 127, 127, -63, 64, 12, -113, 87, 28, -128, -92, -39, 96, 127, 127, -128, -128, 53, -11, 127, 127, 18, -128, -70, 127, 58, 29, -128, 38, 127, -128, -128, 91, 127, -75, -75, -128, 127, -32, 55, -55, -59, -69, 114, 127, -128, 3, 22, -98, -97, 127, 127, 118, -128, -70, -69, 80, 26, -128, -122, 127, -11, 112, -128, 60, -48, -26, -128, 60, 111, -90, 32, 47, -128, -128, 127, 127, -128, 127, 69, 65, -24, -103, -128, 127, 127, 26, -128, -76, -128, 127, 76, -63, -12, 47, 127, -128, 2, 15, -128, -128, 127, 127, -128, -128, 127, 65, 0, -128, -38, 127, 127, -128, -24, 71, -24, -128, 37, 127, 112, -127, 10, -90, -26, -70, 27, 24, 32, -101, 127, 29, -116, -76, 127, 28, 65, 103, -128, -66, 127, 24, -128, 55, 127, -49, -7, 53, 45, 45, -16, -128, -117, 13, -38, 124, 75, -90, 127, 127, -29, -88, -128, 127, -27, 119, -31, -128, 22, 92, 33, -22, 68, -66, -128, -128, 59, 63, -5, 127, 106, -55, -7, 95, -15, 127, -128, 55, 73, 59, 59, -128, 22, -85, -128, 64, 127, 127, -128, 48, -128, 21, 127, -78, -57, -54, 127, -106, -106, 127, 26, 2, -108, -75, 18, 127, 127, -128, -81, 127, -65, -74, -128, 48, -85, 101, 44, -76, -36, 127, -128, -13, 0, -128, 116, -91, 96, -87, 127, -128, 44, 28, -96, 26, -11, -79, 127, 85, -128, -50, 100, 33, -18, -128, 47, 38, 8, -98, 127, 10, 95, -128, -49, -11, -97, 42, -8, 93, -54, -128, 58, 127, -127, -128, 86, 18, 64, 22, 127, -55, 3, -32, -128, 127, 127, -37, -128, 127, 127, 114, 127, -128, -13, -15, -128, -8, 127, 50, -128, 127, 68, 32, -128, 92, 127, 22, -128, 16, -75, 127, -53, -128, 127, 93, -3, -16, 90, -48, -128, -55, -64, 127, -63, -8, -59, 127, -93, -128, -3, 127, -44, -128, 127, -21, -36, 127, -128, -13, -23, 114, -55, -128, -53, 127, 32, 92, 87, -128, 33, 49, -128, 5, 127, 127, -128, -47, 66, -12, 34, 127, -13, -128, -55, 127, -24, -128, -78, 118, 127, -128, -44, -75, 127, -63, -128, 109, 78, 127, -128, -128, 127, 52, -128, -54, 12, 127, -119, 16, 80, -73, -22, 16, 58, -23, -55, -54, -106, 127, 24, 5, 127, 44, -128, -39, -92, 75, 127, -5, -38, -127, -32, 127, -50, 123, -69, -27, 127, 29, -108, 103, -66, 127, -15, -5, -128, 127, -44, -32, 118, 23, -111, -128, 127, -7, -47, 127, 37, -128, 63, 109, -128, -10, -37, 36, 127, -121, -116, -44, 31, -52, 127, -33, -128, -59, 95, 24, -122, 2, 127, -128, -116, -37, 127, -12, -128, 107, 127, 79, -37, -128, 15, 23, -37, -2, 101, 53, 44, -80, -68, 127, 0, 12, -128, -34, 45, 92, -87, 73, 66, -116, -128, 15, 127, 5, -78, -128, -96, 127, -96, 119, 37, -128, 39, 127, -68, -114, -59, 29, -111, 127, -11, 32, 93, 127, -108, -103, 29, 18, -97, 8, 127, -65, -128, 101, -48, -128, 98, 114, -50, -64, -24, 0, 127, -128, -34, 127, -47, 13, -81, -128, 127, -75, 38, -11, 27, -1, -86, 42, 127, 76, -128, 85, 1, -55, -87, -34, 127, 102, -73, 33, 127, -128, -128, 123, 127, 79, -128, 103, 127, -85, -128, 17, 127, 1, -128, -15, 127, -36, -64, -100, 127, 86, 39, -128, -13, 60, 127, -37, -128, -70, 127, -39, 85, 36, -64, -128, 81, 127, -128, 47, -37, -128, -29, 127, -49, -128, 33, 127, -128, -124, -96, 37, 106, 29, -7, 37, 81, -108, -64, 23, -34, -68, -128, 118, -128, -114, 95, 43, -15, -128, 7, -2, 109, -128, -118, 127, 6, -128, 60, 127, -58, 33, -42, -121, -18, 55, 127, -38, -128, 117, 127, -91, 47, -108, -38, 52, 45, -23, 65, 73, -32, 57, -111, -128, 127, 102, -128, -117, 127, 127, -128, -128, -28, 127, 127, -44, -79, -128, 5, 127, 127, -128, 127, -69, 57, -90, 127, -15, -87, 75, 5, 68, -128, -27, 127, 102, -128, -45, -24, 103, 64, -7, -23, -48, -106, 15, -52, 127, -28, 127, -55, 90, -117, 37, 10, 87, -8, -128, 127, 64, 74, 27, -80, -81, 52, 127, -128, 28, 55, -91, -43, 64, 123, 39, -1, -107, 112, 38, 23, -91, -18, 95, 65, -95, 73, -63, 107, -128, -44, 57, 127, -128, -128, 127, 17, -5, -11, -18, -57, 5, 52, -21, 27, -53, 87, -128, 2, -128, -57, 127, 73, -90, -128, 91, 127, -32, -128, -90, 127, -5, 12, 6, 127, 48, -128, -128, -23, 127, 70, 45, 86, -128, -60, 97, 63, 55, -128, -128, 127, -92, -128, -119, 127, -27, -128, 119, 13, 78, -54, -66, 15, 70, -27, -128, -24, 127, -128, 0, 63, -75, -128, 127, 127, -128, 36, 43, 33, -128, -3, 60, -52, 66, 48, -128, 127, 44, -128, 127, 26, -128, 127, 127, -128, -128, 127, 106, -16, -63, 124, -119, 81, 112, 127, -65, -128, -53, 127, -128, -128, 124, 127, 63, -128, -81, -66, 127, 87, -118, 13, 127, -92, -76, -68, 93, 119, -32, -119, 48, -128, -128, 79, 127, -128, -71, 38, 34, 3, 74, -52, 58, -128, 70, 5, 38, -22, -59, -128, 127, 69, -128, 0, -7, 108, 64, 58, -12, -128, 127, 45, 33, -8, 54, -60, -2, -119, -52, -1, 127, -128, 64, 100, 27, -127, 47, 108, 15, -55, 127, -53, -97, 127, 69, -128, 1, 127, 39, -123, -75, 58, 127, -102, -128, 15, 76, 36, 98, 0, -128, -11, -22, -57, -113, 74, 127, 24, -74, -117, 127, 80, -13, -128, 17, 5, 103, -71, -26, -76, -53, -17, -39, -52, 127, -50, -109, 63, 124, -76, -128, 109, 12, 42, 127, -128, -128, -53, 127, 26, -128, 85, -128, 12, -44, -5, 127, 33, -127, -80, 127, -52, 127, -23, -128, -8, 50, 127, 39, -113, 1, -18, 0, 68, 127, -128, -102, 127, -128, 5, 127, -128, -128, 127, 26, 65, -74, -27, -23, -16, -42, -128, 127, 127, -128, -113, 127, -64, -88, -128, -1, 111, 127, -66, -128, -49, 21, -128, 117, 127, 127, -109, -128, 124, 17, -128, 127, 81, -87, -53, -33, 101, -128, 127, 127, -128, 15, 54, -87, -66, 97, 127, -128, 5, -42, -87, -88, 127, 17, -128, 127, 127, 15, -128, 0, 98, -31, 100, 96, -2, -7, 18, -128, 102, -6, -128, 44, 17, -3, 39, 127, -101, 31, 10, 55, -31, -7, 127, 118, -128, -128, 92, 124, 10, -12, -54, -6, 49, 127, -32, -6, -37, 75, -42, 7, -128, 127, 127, -128, 127, 22, -22, -10, -128, 123, 127, -58, 8, 127, -90, -128, 68, 43, 127, -74, 34, -1, -28, 42, -128, 47, 127, -69, -47, -11, -65, 127, 57, 24, -52, 112, -17, -128, -128, 127, 127, -44, -128, 102, 127, -128, -122, 127, 127, -90, 127, -128, -108, -45, 127, -68, 38, -95, 127, -12, 47, 37, 78, -128, 96, 43, 127, -128, 81, -74, 127, -36, -128, -24, 127, -112, 121, -119, -80, 21, 113, 34, -85, -91, -128, 127, -1, 27, 48, 80, 29, -128, 22, 52, -73, -101, 127, -17, -58, -75, 31, 127, 97, -128, -57, 127, 127, -128, 2, -6, 42, -70, -128, 127, 127, -18, 45, 6, -79, -32, 80, -58, -128, 52, 127, -87, -32, 0, 90, 87, -128, 100, -100, 3, 93, 127, -128, -128, -16, -22, 127, 127, -102, -24, 127, -128, -128, 81, 127, -128, -128, 23, 16, -93, -34, 21, 60, -128, -128, 36, -65, -18, 127, 42, -128, 95, 86, 123, -128, -128, 119, -32, -6, -80, 37, 36, -80, -128, 60, 127, 16, -128, -17, 29, -68, 48, 101, -128, -80, 85, 17, -128, -128, 68, 127, 127, -128, -128, 68, 127, 127, -128, -128, 55, 118, -38, -87, 127, 42, -128, -73, 127, -79, 95, -101, 114, -42, -111, 102, -69, -128, 127, 127, -128, -128, 7, 127, 33, -128, -74, 116, -10, 91, -96, -90, 127, -91, -69, -79, 42, -128, 96, 127, 113, -128, -128, 88, 119, -74, 1, -71, -52, -5, 24, -32, 127, 10, 122, -117, -128, 127, 2, -33, 127, -128, -31, -71, -54, -2, 127, -69, -128, 112, 6, -128, 63, 17, -128, -128, 109, 127, 112, 37, -128, -128, 127, 91, -128, 127, 44, -7, -128, 127, 124, 36, -32, -127, 86, 17, 127, -128, -42, 37, -31, -34, 70, -78, -128, -52, 86, 127, 69, -101, -102, -128, 114, 127, 55, 59, -128, -42, 52, -106, 91, -128, -10, -90, 98, 0, -70, -128, 127, 127, 127, -87, -128, -124, 127, 29, -26, 15, 68, 6, 43, 64, 127, -76, 11, -122, -3, 38, -98, -113, 66, 22, 78, -88, 85, -38, -128, -65, 127, 59, -128, -100, 54, -128, 86, 127, 0, -128, 68, 15, -34, 32, 127, -122, -128, -17, 97, -6, -97, 127, 75, -128, -55, 127, 33, -91, 13, 127, -7, 1, -128, 127, 88, -92, 127, 52, -128, -42, 127, 42, -128, -7, 127, -128, -63, 109, 26, -128, 127, 119, -128, -32, 24, -27, 127, 8, -7, -128, 27, 127, -44, -48, 86, 0, -16, -107, 44, -128, 127, -12, -73, 98, 127, -76, -128, 127, 78, -91, -43, 74, 60, 45, 31, -26, -88, 11, 47, -39, -71, -92, -101, 127, 15, -42, 15, 1, -17, -22, -36, 60, 39, -90, 127, 127, -74, -128, 127, 95, -107, 70, -11, -128, 124, 100, -49, -33, -116, 16, 80, -52, -22, -42, 2, 39, 127, -103, -24, 28, 15, -118, 80, 75, -58, -101, -128, 127, 5, 127, -57, 127, -128, 1, 127, 13, -128, 100, 39, -31, 50, -53, -91, -97, 127, -95, 33, -59, 88, -1, 69, -60, 44, 37, 3, 47, 127, 7, 18, -128, 29, -39, 68, -60, 58, -26, -26, -112, 114, 0, 127, -58, -37, 0, -3, 29, 127, -81, -24, 118, -21, 86, -128, -128, 71, -91, 127, 60, -88, -33, 13, 2, 111, 127, -122, -128, 12, 55, 102, -128, 1, 127, -128, -128, 45, 127, -73, -57, -85, 3, 127, -49, -71, -128, -71, 127, 127, 63, -80, -128, -73, 0, -18, 127, 32, 127, -34, -128, 27, 90, 127, -76, -96, -36, -23, 80, -64, -128, 127, 33, -33, -18, 127, -128, -108, 127, -39, -15, -29, -53, -6, 80, -128, 52, -75, -3, 95, 21, 29, -38, -17, 60, -128, 6, -38, -16, 88, -1, -1, 3, -128, 127, 127, -128, 81, 22, -17, -103, 90, 75, -34, 91, 33, 127, -49, -64, -71, 8, -23, 100, 18, -128, -116, 127, -86, -23, 69, -58, -128, 127, -63, -3, 127, 127, -128, -128, -103, 118, -8, 74, -18, 95, 29, 90, -97, -128, 127, 22, -8, 42, 127, -48, -124, -92, -128, 127, -69, 127, -42, -102, -79, 124, 74, 119, -13, -128, 38, 127, -47, -57, 127, -108, -54, -43, -106, 88, 63, -114, 10, -7, -28, 127, -75, 93, 118, -60, -128, 119, 127, -128, 16, 127, -107, 127, -36, -128, 127, 33, -71, 1, 12, -123, 127, -128, -68, 24, -37, 43, -37, 100, -60, 127, -49, -100, 127, 73, -13, 71, -85, -114, 18, 80, 87, -81, 37, 16, -128, 93, -88, -90, 102, 127, -128, -98, -23, 11, -128, 127, 127, -127, -101, 7, -121, 127, 127, -38, 17, -128, 48, -36, 68, 15, 127, -128, -128, -107, 127, 127, 69, -128, -128, 127, -64, 109, -59, 59, 127, -124, -32, -49, -128, 93, 127, -42, -10, 55, 7, -128, 74, 127, 49, 66, -128, 32, -100, -5, 127, -68, -128, 127, -10, -128, 86, 127, 18, -102, -3, -128, -128, 127, 32, -128, 6, 91, 127, -90, -128, -10, 15, 127, 123, 116, -128, 90, 3, -128, 69, 106, -128, 49, 127, 53, -58, -55, -128, 127, 127, -128, -79, 127, -116, 26, -57, 111, -128, 10, 111, 127, -128, -17, -95, -102, 127, 50, -128, -18, 127, 16, -114, 18, 13, 22, -118, 103, 112, 85, 8, -24, 13, -114, -128, 15, 127, 91, -128, 22, 127, 29, -128, 127, 127, -5, -128, -112, 86, 127, 21, 54, -124, -128, -43, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 55, -128, -128, 127, 127, -100, 85, 17, -113, 127, -6, 13, -97, 127, 0, 96, 26, -128, -128, 78, -92, 127, 127, -128, -119, 127, 88, -128, 127, 8, 54, -6, -15, -121, 127, -119, -65, 127, -26, -128, -128, 127, 127, 33, -128, -124, 127, 127, -114, -106, 43, -18, 112, 127, -88, 127, -6, 13, -73, 68, 127, -107, -38, 79, -103, -128, -39, 127, 127, -69, -128, 1, 127, 0, -78, -87, -128, 127, 127, -21, -95, 127, -28, 16, -96, -128, 127, 117, -128, -44, 100, 127, -128, -128, 127, -26, 36, -69, -128, 127, 42, 26, 127, -128, -128, 127, 80, -128, -128, 34, 127, -107, -6, 127, -26, -128, -119, 127, 127, -93, -128, 127, 24, -128, -10, 127, -91, -2, 92, -128, -10, 27, 69, -128, 87, 0, -71, -28, 97, 127, -18, -128, 117, -53, 66, 27, 127, -119, -128, -13, 127, 5, 8, 22, 21, 87, -119, -128, 127, 127, -128, 109, 38, 74, -22, -128, 112, 96, -39, 90, 127, -18, -119, -33, 74, -23, -13, 68, 37, 127, 122, -128, -54, 111, -13, -5, -108, -128, 78, -17, 86, 127, 127, -128, -116, -128, 127, 127, -123, -108, 127, -55, -48, 127, -3, 55, -81, -34, -128, 64, 127, -79, -74, -78, 127, -27, -128, -5, 127, -27, -98, -50, 127, 102, -68, -128, 97, 127, 24, -128, -128, 127, 112, 73, -8, 6, -128, 22, 78, -8, -128, 15, 127, -28, -128, -38, 127, -45, -128, 123, 76, 1, -24, -27, 127, -128, 106, 28, 112, -2, -128, 2, 86, -81, 44, 127, 63, -128, -3, 127, 27, -54, -34, -7, -128, -11, -39, -39, 55, -128, -128, 70, 127, -128, -38, 127, 127, 0, -128, -52, 127, -71, -54, -96, 1, 96, 127, 1, -97, -109, 111, 103, 74, -92, -128, 127, -43, -12, 0, -38, 117, 127, -128, -75, 127, 44, -128, 127, -11, -128, 55, -3, 127, 2, -32, -128, 127, 65, 31, -52, -36, 38, 109, 5, -128, -90, -45, 0, 127, -49, 47, -18, 24, 8, -128, 47, 127, -58, -63, 58, -17, -119, 85, 102, -75, -86, 26, -55, 85, 127, -128, -128, 127, 127, -128, -68, 65, -128, 70, 74, 29, -128, -24, 127, -28, 68, -87, -128, 127, 127, -128, -66, 127, 76, -128, -128, 127, 127, -128, -44, 127, -128, -81, 47, 127, 76, -128, -128, 39, 127, 97, -57, -2, -128, 54, 127, 119, -128, 48, -128, 124, 118, 127, -128, -111, -74, 127, 66, -128, -128, 127, 60, -39, -26, 49, 96, 15, 36, -128, -28, -128, 127, 127, -128, -38, -15, 91, 6, -53, -3, 127, 122, -128, -128, -76, 68, 86, 111, 127, -106, -128, -128, 66, 127, 73, 5, 11, -128, 49, -128, 64, -26, 1, -128, -11, 127, 65, -119, 85, -50, 53, -81, -45, -128, 34, 127, 102, -63, -117, 78, -128, 44, -37, -69, -12, 127, 86, -128, 23, 127, 39, -107, -128, 75, 59, -17, 17, 63, 79, -70, 60, 127, -11, -128, -48, 127, 127, -24, -128, 16, 127, -44, -45, 39, 11, -34, -113, 127, 85, 127, -18, -128, -74, 81, 112, 73, -90, 86, -128, -78, -58, 107, -8, 7, 10, -39, 102, -12, 69, 127, 114, -128, -1, 7, -101, 101, -21, 87, 90, 26, 59, -90, -29, 32, -68, 80, 16, -128, 63, -58, -81, 13, 2, -128, 95, -54, 22, -64, -27, 31, -18, -128, 127, 127, -90, 54, -31, -128, 17, 60, 127, 10, -108, -108, 127, -6, -96, -128, 127, 127, -8, -128, 117, 53, 127, -112, -52, 127, -47, -128, 38, 48, 23, 127, 54, -128, -52, -65, -23, -52, 127, 27, -128, 127, 127, -128, 66, 57, -45, -128, -49, 127, 127, -118, -128, 127, -98, 127, -43, -15, -12, 47, -103, -112, 127, 121, -128, 0, 127, 116, -128, -16, 127, -128, -57, -10, 124, 58, -69, -128, 101, 122, 26, 50, -38, -128, 127, -38, 2, 73, 65, -8, -128, 121, 127, 71, 106, -128, 37, -48, -128, 121, 65, 34, -124, 50, 38, 53, 69, 127, -128, -49, -128, 117, -128, 86, -27, 91, -32, -97, 117, -2, -128, -124, 7, 53, 55, 127, 13, -128, -5, 127, -70, -128, 60, 18, 8, 88, -88, -36, -7, -98, 127, 90, 16, -32, -34, 74, 127, -59, -128, -37, -11, 114, 60, 127, -86, -128, 2, 43, -39, 103, -45, 52, 127, 92, -128, -109, 78, 27, -92, -93, 127, 113, -128, 48, 127, 78, -128, 16, 33, -127, 124, 76, 55, -128, 44, 127, 91, -128, 66, -36, 49, 45, -97, -54, 116, -57, 0, -128, 127, 127, -128, -18, 127, 22, 54, 12, -128, -22, 127, 29, -128, -52, -33, -27, 127, -49, -128, 127, 127, -64, -128, 127, -108, 39, 127, -128, -73, -15, 127, -113, -24, -52, 122, -128, -80, -48, 88, 69, -13, -109, -47, -128, 106, 127, 114, -59, -98, -6, -57, 127, -3, 7, 127, -1, -128, -71, 66, 75, -70, 2, -5, 44, -128, -29, -47, -128, 71, 44, -29, 124, 42, -36, 127, -128, -128, 127, -76, 80, -45, -128, 127, -113, -42, 101, -117, 10, 108, -128, 31, 27, 69, 53, -128, 76, 127, -23, -128, 90, 27, -128, 106, 18, -101, -6, 127, 52, -128, -2, 127, -28, -128, -93, 127, 127, -128, -36, -114, 81, 50, -23, -93, 79, -66, -74, -121, -34, -88, 127, 127, -64, -128, 127, 24, -128, -39, 127, 74, 65, -124, 87, -1, -128, -45, 127, 127, -63, -93, -60, 24, -70, 10, 127, -12, -100, 55, 127, -68, -128, -103, 127, -8, 12, 101, -128, -33, 53, -128, 6, -49, -52, -128, 127, 127, -123, 75, -8, -121, 10, -11, 53, 91, 6, 21, -26, -128, 55, -128, 127, 12, 10, -21, 1, -32, 49, -118, 127, -7, -21, -107, 86, 127, -118, 21, -101, -85, 85, 127, -128, -31, 42, 118, 10, 44, -101, -74, 70, -128, 73, 127, -128, 11, -60, -128, 127, 113, -109, 2, -1, 10, 55, -47, -3, 127, -128, -1, 66, 88, -68, 45, -111, 118, -114, -128, 75, 127, -128, -43, -10, 24, 96, 12, -128, -128, 123, 127, 108, -112, -128, -128, 71, 124, -128, 0, 127, 57, -7, -124, -95, 21, 1, 127, 15, -21, -128, -48, 127, -32, -111, 0, 127, -128, 32, -128, -50, 127, 69, -128, -102, 81, 127, -128, -114, 127, -59, -128, -2, 127, 31, -128, 58, 127, -58, 27, -11, -128, -97, 127, 127, -128, -7, -65, -12, -128, 121, 36, 127, 69, -128, -28, 21, -102, -74, 127, 127, -60, -60, -32, 127, -128, 65, -34, 5, 127, -21, -88, -48, -90, 32, 91, 0, 106, -128, -128, -57, 23, 106, 38, -128, 127, -64, -36, 127, 32, -128, -128, 123, 127, 96, -50, -100, 2, 127, 127, -88, -128, 75, 74, -76, 15, 127, -52, -88, -54, 127, 17, -96, 34, 23, -47, -23, -128, 6, 127, -98, 48, -87, -128, -38, 127, 90, -39, 119, -128, -13, -78, 127, 28, -85, -128, 109, 102, -128, 74, 127, 3, 10, -121, -39, 85, 64, -38, -95, 70, -128, -71, 127, -8, -75, 103, -26, -128, 79, 127, -21, -76, 0, 127, -128, 24, -23, -123, -65, 34, 45, 107, 42, 127, -24, -128, -64, 36, 109, -53, -128, 78, -42, -39, 127, 11, -69, 55, 95, -128, -111, 127, -12, -112, 127, 127, 45, -128, -91, -128, 127, 114, -52, 37, 79, -66, 103, -127, -128, 79, 64, 73, -75, -128, 127, 0, -128, -118, 127, -55, -10, 57, 121, -128, 127, -98, -79, -37, 22, 63, 23, 37, 119, -55, -90, 13, 114, 21, -128, -15, 127, 27, 73, -116, -86, -55, 15, 13, 3, -128, 127, 22, -118, -8, 127, -45, -128, 127, -26, 74, 32, 127, -128, 1, -38, -43, -65, 59, -23, 108, 127, -32, -128, 87, 127, -128, -128, -36, 127, -128, 5, 38, 69, -128, 127, -10, -74, 55, 103, -12, -47, -128, -31, 127, 65, -128, -58, 127, -85, -33, -128, 7, 127, 127, -128, -128, 28, 96, -128, -74, 127, 6, -8, -128, -5, 127, -43, -107, 127, -80, -59, -63, -17, 49, -90, 23, -128, 53, 127, -21, -78, -74, 15, -128, 81, 127, -88, -21, 15, 17, -128, -102, 127, -117, 101, 48, -113, -128, 63, 127, 81, -128, -128, 127, 60, 26, 98, 127, -128, -8, -92, 90, 24, 127, -90, 12, 127, -128, 24, -70, 100, -102, 64, 108, -128, -98, -11, -128, 127, 119, 127, -119, -128, -10, 127, 127, -128, -124, 119, 127, -13, -86, 21, 0, -128, 100, 127, 7, -75, -100, 108, 64, 28, -128, 97, 127, -128, 11, 127, -59, -128, -28, 91, 102, 127, -128, -85, 32, -29, 1, -78, 33, 127, 26, -117, 59, -79, -91, 88, 101, 24, 34, -73, -42, 68, -52, 7, 127, -127, -106, 68, -57, -18, 127, -127, -17, 127, -44, -88, 24, -27, 119, 1, -128, -3, 127, -121, 112, -128, 36, -36, 127, -98, -106, -128, 127, 81, 5, 64, 55, -128, 127, -37, -98, -91, 92, 127, -128, -8, -98, 70, -32, 100, 96, -128, -128, 65, -3, -73, 50, 127, 0, -128, 64, 127, 17, -128, 87, 1, 100, 122, -100, -98, -119, 127, 92, -128, 127, 50, 21, 71, -128, -31, 109, 109, -128, 8, -57, 65, 113, -16, -97, -11, 127, -23, 24, -88, 127, 55, 86, -27, -53, -54, -33, -128, 127, 127, -22, -58, -5, -55, 92, -66, 127, -112, -13, -6, 121, -50, 1, -18, -7, -36, 114, 90, 52, 117, -128, -128, 28, 127, 53, -128, -128, 28, 54, 127, -128, -86, 76, 74, -100, -37, -6, 36, -128, -128, -128, 127, 54, 111, 102, -55, -81, -37, 22, 54, -128, -116, 127, 127, -128, -27, 127, -29, -121, -10, 106, 39, -44, -31, 16, -76, 15, 76, 127, -128, -128, 97, 127, 21, -128, 65, 127, -128, -63, 127, -38, -128, 22, 111, -128, 96, -74, 88, -38, -54, 107, 21, -128, 7, 98, 127, -49, -69, -128, -13, 127, 32, -128, 49, 2, 127, -57, 38, 0, -80, -78, 5, -28, 127, -31, -128, 102, -66, 54, 127, -21, -128, 111, 15, 81, -49, -128, -92, 116, 17, 16, 29, -1, 53, 127, -114, -7, -87, 116, 49, 80, -128, -69, -26, -48, 127, -15, 26, 36, 68, -34, -128, 127, 127, -75, -60, 127, -128, 45, -128, -39, 36, 127, -128, 52, -121, -107, 37, 127, -128, -128, -37, 127, -128, -34, 81, 15, 103, -128, -128, 86, 97, 16, -44, 2, 21, -108, 127, -103, 127, 39, -119, 6, -33, 127, -128, 70, 127, -3, -128, -23, 127, -69, 16, 43, 127, -101, -128, 27, 121, -85, -31, 127, 116, -69, -95, 68, 127, 24, -15, -97, -33, -43, 15, -57, 70, 127, -128, 127, -65, -34, 57, 127, -47, -128, -128, 37, 59, 59, 87, 92, -128, -128, 127, 63, -128, 98, -65, 58, 12, -90, 127, 16, -128, 127, 127, -128, 60, 127, -128, 100, 127, 92, -97, -128, -49, 127, 124, -16, -128, 127, -17, -128, 113, 101, -128, 73, 16, -114, 0, 127, 28, -128, 3, 127, -64, 68, 49, -75, -86, 80, 127, -117, 28, -75, -29, 118, -64, -128, -121, 127, -122, 68, -54, -106, -78, 127, -58, -128, -96, 127, 48, -98, -22, -52, -50, 127, -49, 106, -122, -128, 50, 127, 127, -128, -128, -65, 127, -71, 127, -49, -113, 38, 127, 38, -128, -128, 127, -52, -2, -26, 3, -71, 47, 127, 81, 98, -128, -93, 127, -100, 33, 47, -123, -127, 102, 127, -74, -74, -16, -97, 127, 116, -128, 38, -5, 97, 18, -128, -65, 127, -16, -128, -128, 127, 127, -128, -49, 65, 127, -86, -128, 75, -1, -128, -58, 127, 90, 38, -128, 127, 111, -23, -101, -64, 127, 28, -128, -65, 127, -75, -15, -48, 0, 54, 59, 127, -128, -128, 33, -128, 127, -87, 127, -42, -128, -43, 127, -117, 24, 127, -52, -111, -128, 122, 127, -122, -32, 5, -79, 121, 102, -12, -64, -58, 23, -128, 95, 49, -103, -128, 59, -28, 121, 127, 127, -48, -12, 2, -44, -128, 32, 127, 29, -21, -17, 43, -128, -107, -3, 127, -42, -128, 127, 32, 6, -128, 127, 0, 29, -128, 70, 90, 55, -16, -73, -73, -15, 127, 8, 47, 34, 92, -128, 15, 127, 70, -128, -128, 127, -124, 123, 0, -17, 66, -2, 66, -128, 21, -79, 45, 29, -128, 23, 109, -128, 16, 1, -128, 111, 45, 7, 29, -6, -102, 90, -17, 23, 87, -42, -79, 127, 71, -86, 127, -123, 87, -23, -53, 12, 58, -128, 43, -43, 90, 117, -128, 102, 3, -31, -116, 116, 79, 101, 36, -128, -128, 127, 103, -128, 43, -92, 114, -42, -128, 18, 78, 18, 116, -48, -55, -128, 127, 52, 10, 12, 10, -107, -13, 12, -127, -24, -71, 60, 28, 107, -128, 97, 127, 0, 43, -128, 81, 11, -128, -95, 116, -66, 28, 127, 108, -128, 59, -128, -128, 127, 60, -80, -111, 127, 97, -54, 127, 127, -128, -10, 11, 45, -10, 90, -73, 87, 116, -58, 1, 127, -53, -128, -2, 31, 96, -75, -90, 34, 22, 28, -49, -128, 127, 102, -11, -66, 80, -28, 78, 127, -112, -114, 22, -128, 37, 127, 127, -76, -128, -47, -15, 127, -95, -128, 86, 79, -23, -26, -26, -42, 10, -128, 44, -48, 42, 90, 127, -85, -128, -128, 65, 60, 112, 92, -16, -128, 127, -31, 69, -76, -54, 127, 127, -128, -87, 100, -39, 69, 0, 88, 97, -116, -128, 103, -128, 54, 127, 21, -128, 63, 127, -128, -128, 97, 127, 44, 22, -128, -128, 127, 5, -66, 36, 68, -103, 1, 127, 71, -81, -57, -127, -87, 76, 45, 65, -7, 98, -54, -128, -128, 127, 43, -73, 64, 127, -27, -128, -32, 127, -50, -128, 108, 90, -128, 127, -1, -88, -59, 127, -10, -28, 34, -86, 32, -97, -128, -118, 32, 127, 103, -116, -8, -54, 127, -36, -68, -128, 127, -16, 38, 127, -128, -39, 127, -58, -128, 74, 127, -64, 33, -8, -15, -42, 92, 127, -123, 10, 127, -34, -128, 127, 33, -60, 58, -2, 29, -53, -69, -128, 127, 86, 37, -102, 49, 27, -128, 75, -3, -107, -55, -21, 112, -128, 88, 127, -128, -117, 127, -34, -128, 127, 7, 13, -60, 96, -79, -87, -128, 127, 127, -50, -128, 86, 114, -43, -128, 17, -87, 127, 73, -128, 73, 76, 76, -16, -31, 8, -114, -95, -5, 127, -123, -128, 16, -54, 98, 127, -45, -5, 76, 26, -128, -112, 0, 127, 118, -128, 113, 31, 109, -128, 23, 127, -7, -128, -47, 6, 95, 114, -33, -128, -128, -34, 127, 54, -12, 127, -128, -128, -7, 127, -128, 127, 54, -10, -128, 127, 55, 121, -128, 127, -43, -102, -128, 127, -68, 127, -119, 12, 103, 52, -68, -3, -28, -128, -128, 96, 127, -81, 92, 57, -55, -128, 1, 127, 127, -80, -128, -128, 103, 127, -12, -128, 59, 7, 127, -39, 127, 10, -101, -45, 127, 127, -128, 47, 127, -98, -128, 103, 127, 119, -128, -79, 88, -71, -128, 8, -7, -15, 27, 33, -49, -128, 127, -31, -128, 75, 0, -29, 127, 65, -128, -26, 127, 127, -128, -116, -69, 119, 127, -66, -128, 127, 113, -27, -117, 6, 127, -5, -117, -92, 127, -69, -122 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
