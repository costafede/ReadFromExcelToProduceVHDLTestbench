-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            2, 9, -2, -15, -16, -4, 13, 14, 18, -7, 7, -12, -20, -6     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -61, -123, -69, -88, 28, -31, -70, -68, -84, 83, 105, 74, -76, 10, -108, 26, 73, 21, 24, -1, 40, -62, -74, -85, -75, -126, -69, 4, 59, 51, -72, 83, 45, -102, -86, -8, -46, -78, 70, 96, -100, -67, -11, 30, -74, 50, -126, -109, 29, -4, 111, -29, -46, 74, -117, -26, 86, -107, -90, -41, 71, -75, 112, 84, 14, 98, -27, 12, -86, -96, -49, 127, 64, -15, -105, -109, 127, 103, -103, -63, -64, 74, -44, -5, 58, -79, -104, 6, 12, 57, 32, 1, 55, 58, 77, 6, 33, 31, -13, 113, 71, -6, -104, -37, -119, -74, 1, 111, 80, 57, -38, 12, 103, 98, -5, -80, 36, 84, 4, 49, -69, 29, -31, -88, -108, 16, 63, 20, 75, -43, 105, -15, 126, -112, 78, 123, 0, 127, -40, 37, 91, 12, -127, -61, -17, 11, 12, -111, -94, -75, -32, -60, 6, 45, -56, 25, -28, -58, 56, 69, -47, 86, -127, -72, 86, 19, -75, -90, -107, 104, 112, 51, 39, 5, 37, 19, -49, 13, 37, -16, 55, -48, 23, 13, -40, -5, -62, 58, 98, 98, -49, -117, -29, 52, -1, -31, -76, 4, -6, -77, -51, -24, -23, 90, 2, 99, -83, -44, 98, -41, -116, 0, -90, -61, -98, -31, -88, -106, -3, 71, -15, -24, 68, -128, 12, -35, 8, 105, 101, -58, 90, -58, -96, -47, 32, 126, -10, 69, -36, -97, 125, 2, 68, -90, -3, 0, -45, 27, 101, 98, -88, -126, -49, -105, 119, 56, 116, -66, -97, -50, 88, -97, 32, 7, 126, 38, -22, 79, 6, 30, -31, -77, 72, 4, -77, 76, 81, 79, 85, -65, 2, -45, -85, 87, 85, 7, -103, -81, -72, 116, 114, 65, -98, 76, -49, 99, 25, -110, 79, 70, -45, 3, -78, -70, -7, 115, 106, 51, 7, 75, -107, -34, 96, 32, -85, 101, 93, 22, 11, -37, -110, 9, -101, -101, 81, 95, -61, 125, -50, 73, -63, 84, -84, -101, 111, 54, 86, -32, -88, -64, 55, -60, -63, -78, -118, 24, -76, -40, 120, -50, 12, -50, 30, 1, 11, 62, -87, -89, -14, -33, -17, 113, -98, 75, -31, 122, 88, -20, 3, -19, 79, -9, 124, -27, -3, -83, 104, -51, -30, 121, 112, 26, 98, -31, 59, 26, 72, 89, -76, 13, 38, -6, 96, -24, 25, 41, 24, 80, 42, -42, -15, -9, -44, -16, -103, 74, -51, -53, 62, 22, 68, -92, 126, -120, 39, 92, 35, 20, -13, 107, 55, 78, 17, 115, 116, 82, 49, -126, -85, 7, 44, 2, 113, -18, -39, -115, -76, -119, -5, 51, -33, 13, 79, -43, 124, -73, 22, -36, -50, -33, -111, -104, -76, 48, 1, -62, 90, -85, 87, -93, -103, 49, 50, 88, 63, -2, -41, 109, 84, -115, -58, -84, -109, 110, -58, -24, -56, 95, 20, -40, 120, -71, 15, -46, -108, 81, 72, -51, 85, 43, -84, 88, 84, 54, -53, -50, 56, -74, 73, 120, -52, 56, -55, -23, -40, -88, -88, -4, -98, 15, 120, 88, 108, 95, -67, -113, 3, 36, 127, -92, 87, 8, 65, 123, -98, -33, -104, -30, 95, 59, 61, 42, -4, -20, -46, -16, -62, -83, 53, -82, 58, -28, -86, -11, 38, 25, -67, -96, -73, 85, -97, 73, 31, 19, -34, 100, -33, -100, -107, 11, 17, 30, 119, 77, -56, -96, -85, 93, -70, 13, -37, 6, 110, -111, 127, -90, 65, 48, -1, -50, 64, 111, -56, 83, 87, 124, 21, -84, -26, -97, -30, 12, 94, -40, -56, 105, -16, 31, 26, -40, -85, -6, -100, -34, 94, 93, 59, -49, 11, 83, 95, -8, -49, -47, -105, 94, -111, 19, -56, 112, -64, -20, -64, 90, -33, 66, 127, 19, -97, -18, -37, 32, 63, -52, -87, -62, -107, 53, 83, -50, -61, -111, 126, -42, -16, -100, -119, -128, 77, 34, -74, 40, -118, 62, 70, 26, 104, 57, -30, 124, -37, -121, -30, -47, 34, -20, -97, 61, -113, -32, 32, -38, 126, -43, -7, -110, 68, 38, -41, -21, -75, 106, 65, -74, -39, -60, 48, 7, 110, -58, -11, -72, -13, 35, 52, -111, 48, 11, -12, -78, 82, 120, -43, 126, 15, 7, 65, 30, -11, 97, -122, 31, -63, 86, -66, -68, 23, 108, 100, -29, 36, -63, 14, 38, -70, -24, 99, -50, 30, -71, 70, -121, -51, 32, 82, -47, 107, -58, 121, -101, 100, -56, 95, -45, 42, 22, -40, -100, 105, 104, 127, -90, -75, -84, -67, 91, -116, -120, 82, -1, 7, -10, -110, -64, -92, 38, 19, -87, -16, -6, -2, -16, -63, 19, -48, -9, 11, 125, 121, -71, -127, 83, -102, -59, -121, -54, -91, -83, -35, 55, 110, -12, 16, 110, -101, 4, -34, 14, 22, 68, -109, 96, 15, 82, -85, 2, -47, 33, 91, -35, 120, -87, -115, 9, 16, 43, 14, 77, -75, 7, -109, -122, 123, 74, 28, -22, -86, -113, 125, -52, -23, -104, -126, -36, -11, 117, -80, -61, -91, 21, 39, 78, 17, 18, -18, 108, 66, -58, 109, -21, 40, -116, -20, 114, -13, 48, -104, 82, 89, -121, 31, 41, 119, -3, -41, 34, -75, -83, -64, -102, 32, -75, -24, 97, -35, -61, -4, 53, 57, 109, 59, 118, -90, 6, -85, 119, 21, -89, 79, -127, -18, -6, 127, -128, -25, -101, 33, -19, 97, -53, 118, -34, -59, 83, 37, -60, -39, -109, -41, 99, -45, -111, 69, 38, 70, -102, 43, 119, -105, 26, -8, -79, 113, 87, 72, -67, -26, 6, 3, -16, -43, -82, -113, -118, -39, -99, 109, -17, -104, 84, -58, -33, 119, 110, -22, 95, -124, 26, 100, -106, 123, 31, -49, -103, 54, -72, -114, 35, 106, 9, 121, -58, -51, 65, -55, -100, -127, -90, -106, -47, -66, 95, 88, -90, 89, 117, 98, 97, -28, -84, -61, 121, 52, -83, -123, -41, -34, 111, 43, -126, -54, -1, 85, 59, 94, -25, -92, 30, -88, -6, -22, -55, 115, 72, 92, -46, -9, -64, -110, -42, 80, 92, -76, -70, 22, 58, 47, -127, 63, 90, -43, -80, 51, 69, -8, 119, 98, -34, 62, 125, -22, 20, -64, -87, 48, 79, -27, 106, 79, 92, 56, -1, -7, 21, 110, 28, 76, 40, -16, -102, -89, -104, 59, 44, 52, -72, -111, 75, 0, -43, -122, -48, 66, 39, -59, -79, -124, -66, -86, -57, 69, 127, -74, 5, 45, -106, -63, -94, 109, -44, -69, -49, -6, -13, 82, 10, 43, -100, -82, -122, 124, -12, -22, -107, -24, 26, -19, -42, -106, -48, 73, 92, 33, -68, 84, 40, -8, -10, -53, 126, -44, -18, 101, 99, -88, -111, -37, 125, -124, 84, -84, -31, -117, -11, -36, 52, -121, 78, 35, -74, 126, -81, -96, -81, 100, 47, -110, -21, 58, 112, -107, 119, -124, -9, 27, 21, 83, 98, -126, 90, -22, 122, 74, 41, -30, -29, 12, 88, -3, -110, -18, 91, 30, 112, -105, -89, -33, -52, -126, -1, -27, -58, 70, 9, -126, 126, 74, 62, -1, -13, 45, -118, -28, -96, 62, 91, -8, -87, 119, 74, -127, -76, -80, 39, -12, 113, 90, -80, -125, -72, 72, -52, -67, -61, 14, 95, 84, -6, 64, 28, -41, 8, -99, -9, -123, -24, -15, 91, -77, -101, -50, 88, 60, -19, -54, 116, 99, -108, 120, -44, -56, -82, -45, 40, -107, 82, -67, 63, 93, -77, 1, 84, -98, 4, -50, 27, -24, 40, 11, 61, 10, 27, -2, 84, -120, -123, 108, -31, 115, 35, -118, 106, 104, 68, 85, 30, -1, -28, 72, -37, 14, 7, 52, 89, -5, -31, -84, -69, 14, -46, 50, -118, 62, 86, -59, 43, 2, -8, -47, -111, -38, -110, -47, 48, 111, -79, -50, -16, -121, -32, 34, 98, -70, -120, -69, -52, 7, 32, 112, -90, 76, -72, 7, -50, -43, -43, 82, -58, 51, 85, -18, 8, 71, 96, 103, -69, 50, 70, 45, 103, -27, -128, 32, -6, -43, -20, 10, 77, 75, 7, 84, 27, 13, 25, 35, 89, -57, 113, -44, 12, -28, -86, -61, 68, -60, -24, 37, 94, 41, 48, 96, -118, -119, -18, -42, -75, -105, 60, -109, 84, 102, -82, 45, -2, 26, 15, 40, -13, 64, 20, 66, -90, 69, 61, 2, -24, -66, -11, -59, 76, 28, 60, 92, 20, 57, 94, -102, 76, 58, 50, 126, 122, -110, -94, 78, 55, 117, 124, -17, -8, -56, 67, -70, 91, -111, 103, -81, 31, 100, 12, 52, 94, -110, 31, 5, -62, 120, -47, -76, -106, -109, -19, 123, -14, -88, 126, -10, -20, 56, 88, -97, 87, -30, 56, -87, -53, -113, 10, -29, 107, 115, 114, -91, -48, -117, -21, 117, 13, -42, 3, 108, 108, 119, 75, 83, -52, 6, -21, -116, 49, 34, 74, -48, 120, 113, 87, 88, 126, 36, -40, 98, -51, 63, 44, 68, 22, -124, 117, 29, -18, 104, -49, 103, -74, 9, -69, 59, 56, 19, 5, 75, -62, 29, -21, 39, -104, -19, 86, -2, -53, -86, -60, 125, -11, -94, 116, -87, -86, -112, -101, 45, -88, -31, -43, -41, 72, 20, 73, 33, -26, 25, -25, 63, 51, -26, -35, 19, 96, 109, 50, 127, -88, 88, 14, 124, -34, -54, 105, -56, -9, 88, -1, 41, 65, 9, 93, -121, 76, 54, -68, -85, 10, -70, 87, -62, 34, 68, 35, 27, 32, -91, 114, -100, -32, 21, 99, 106, 6, 61, -32, 67, -28, 6, 27, 18, -22, -26, -122, -86, -26, -125, 81, -123, -26, 39, -39, -48, 110, -64, 26, 124, -57, 28, -65, 111, 62, -19, -24, -56, 35, -123, -27, 50, -74, -6, 58, -18, -72, -126, -125, -2, 116, -89, 12, 71, -58, -26, 110, -50, -10, 77, -126, -39, 39, -125, 19, 111, -67, 74, -72, 102, -48, 75, -53, -52, 76, 18, 80, -3, 113, 13, -29, -35, -3, -58, 73, -27, -74, 38, -74, -71, -62, -59, 68, 58, -116, 26, -76, 53, -104, -113, 16, -95, -44, 72, -27, -40, 38, -23, -24, 40, -58, 120, -95, -115, 53, 82, 51, 42, 98, -61, -46, -42, 92, 68, 116, -23, 60, -123, 20, -117, 24, -64, -22, -82, -31, -74, -112, 29, -85, 79, -97, -66, -91, 34, -47, 0, -79, -36, -39, -4, 122, -90, 23, -110, -105, 93, 125, -104, 33, 22, 59, -110, 22, 118, -50, 92, -13, 77, -29, 29, -37, -71, 64, 49, 60, 123, -93, 20, 43, 109, 88, 112, 108, 50, 74, -48, -82, 19, 37, -78, 120, 34, -22, 85, -89, -32, 114, -59, 117, 122, 84, -21, -126, -92, 0, -67, -85, 86, -41, 11, -59, -77, 27, -127, -15, 47, -61, -107, 14, 0, -54, -73, 89, -107, -35, 78, -53, -39, 96, -1, 122, 2, 23, 84, 10, 28, -59, -96, 105, -6, 64, 71, -29, 73, 40, 113, 1, 13, 43, -25, 114, 11, -116, 119, 93, -13, 77, 110, -122, 2, -31, -92, 35, -59, -47, 38, -96, 1, 13, -70, 0, -122, 41, 114, -16, 49, 29, -117, -101, 82, -39, 105, -121, 52, 55, 97, 38, 98, 97, -24, 108, 12, 127, 47, -2, -58, -33, 26, 19, 69, 42, 101, -21, 63, -3, 94, -112, -122, -49, -90, 70, 52, -76, 78, 75, 79, 98, -8, 37, -13, 89, -27, -21, 111, -93, 36, -115, -105, 91, -45, -77, 113, -53, 47, -9, 103, 112, -26, -58, 71, 113, 95, -10, -90, -21, 11, -90, 104, -23, 44, -51, -82, -37, -71, -72, 65, -101, -16, -20, -44, -28, -92, -34, 116, -28, 47, 37, 31, 9, 106, 70, -89, -97, -37, 20, -9, -14, 107, 119, 88, -108, 75, -55, -113, -94, -6, 77, 24, 60, 16, 69, 53, 86, -72, -72, 12, 90, 93, 114, -52, 114, 63, 22, 100, -76, -117, -122, 58, -48, 103, -72, -14, 95, -41, -35, -90, 49, 22, -43, -104, 19, -54, -14, -60, -7, 35, 26, 82, -51, -121, -33, 121, 46, -50, -5, 13, 19, -54, -72, 104, -89, -43, -10, 72, 53, 41, 71, 3, -83, -11, -56, -123, -70, -112, 110, 107, 89, -39, -107, -5, -12, 66, 5, -28, 76, 30, 94, 43, -40, 78, 6, -107, 22, -76, -33, 62, 95, -55, 49, 115, -80, 38, -119, 127, -28, -84, -76, -75, 95, -119, -125, 45, 20, 118, 60, -54, -54, -65, -13, -47, 105, -117, 17, 106, 3, 38, 21, 102, -81, -69, 28, 7, 6, -128, -12, -44, -102, -114, 32, -17, 108, 81, 37, -127, 12, -24, -118, -64, 11, -1, -33, 125, 4, -105, -78, -69, -107, 85, -21, 9, 115, -30, -19, -73, -90, 18, -11, 122, 23, 54, 90, 41, 53, -78, -12, -32, -106, -89, -105, 51, 42, 30, -86, -87, 78, -121, 43, 52, 66, 119, -63, 64, 0, -101, 95, 64, -36, 91, 18, -36, -74, 19, 43, -61, 0, -113, 124, 77, -17, -119, -26, -80, -82, -3, 87, 51, -49, 60, 95, 10, 75, 24, -32, 50, -28, -4, 75, -113, -85, -126, -50, 104, 11, 94, -28, 112, 53, -63, 71, 28, 42, -37, 78, -62, 71, -31, -55, 52, -18, 90, -22, 18, 111, 66, -36, 6, -51, 64, -109, -25, 68, -65, 6, 56, -51, 97, -127, -59, 87, -59, -87, 23, -82, 38, -96, 48, -58, 126, 41, 11, 126, -51, -86, -29, -33, -26, 51, 64, 73, 6, -14, -69, 77, 39, 92, 111, 7, 81, 108, 1, 118, 5, -31, 95, 59, 98, -93, -42, 24, 59, 88, -21, 49, 77, 92, -117, 71, -88, 86, 80, -40, -54, 14, -119, 98, -24, -43, 62, -62, 45, 33, 14, 83, -19, 85, 15, 90, 119, -1, -22, 85, -89, 107, -51, -86, 65, -128, -48, -113, 54, 119, 113, 42, -1, 65, 52, -84, 0, 11, 99, -77, 66, -28, 95, 23, -118, -44, -50, -29, -121, 8, 122, 69, -37, 107, -67, 77, -1, 71, -17, 86, -4, -74, -51, -106, -16, -96, -52, 87, -97, -82, -57, 127, -49, 34, -86, 86, 43, 114, 50, 41, 79, 93, -106, 0, 1, -46, 85, 14, -114, 125, -8, -23, -28, -20, 74, -42, 67, 65, -116, -63, -61, 115, -126, 32, 57, 17, -19, -9, 81, -65, -44, -127, 73, 115, -112, -8, 90, -7, 81, 93, -42, -52, -101, 120, 28, 92, -74, -61, -126, 34, 58, -62, 74, 87, -105, 6, 105, -44, 44, -7, 64, -71, 47, -14, 77, 52, -39, -87, -8, 29, -70, -33, 90, -34, 82, 34, 1, 65, -126, -109, -57, -7, 56, -40, -72, 17, -33, -17, -127, -84, -27, -14, 61, 27, 97, 55, 38, -74, -101, 14, 108, 4, 73, 13, 44, -82, 4, 34, -33, 44, 94, 110, -24, -41, 119, 7, -75, 21, -12, -13, -57, -89, -86, 39, -26, 108, -11, -49, 11, 74, 36, -110, -128, 49, 30, -58, 20, -91, 4, 30, 65, -20, -77, 51, 41, -16, -107, 14, 9, -113, -42, 56, -12, -65, 32, -3, 26, -4, 70, 73, 75, -99, 73, -123, -77, -92, 5, -120, 96, 49, 113, 18, 46, 80, -91, -58, 81, 21, 81, 113, 15, 26, -30, -32, -77, 96, -19, 127, -58, 62, 94, 73, -5, 21, -30, 17, -12, 33, 100, -21, 72, 126, 49, 2, -111, -85, 38, -12, -23, 52, -85, 45, -38, 46, -15, 101, 11, -12, 100, -44, -59, 88, -18, 86, 51, -94, 71, 104, 90, 59, 71, -93, -28, 23, -16, -128, 3, -49, -123, -120, 26, -58, -128, -46, -94, 105, -99, -27, 13, 25, -33, 95, -58, 112, -100, -9, -36, 64, -61, -31, -56, 76, -17, -32, 19, 82, 127, -37, 117, 30, 53, -109, 64, -65, 46, 71, -75, 91, 76, -71, 5, -32, -116, -49, 121, 73, 109, 104, -78, 120, 96, 75, -12, 124, -124, -111, 118, 77, 118, -77, -36, 103, -19, 125, -119, 88, 11, 93, -113, -70, 116, -5, -116, -73, -80, 118, 29, -86, -97, 72, -101, -89, -103, 114, -105, -43, 3, -99, -11, 81, -40, 109, 23, 23, -108, -45, -116, -32, 31, -119, 116, -64, 20, 56, 67, -88, 72, 115, -7, 100, -31, -58, 105, -25, 14, -115, 25, 94, 81, -125, 121, -46, -5, 81, 67, -81, 13, -29, -37, 20, 119, -27, -20, -30, 46, -126, -85, 69, 91, 117, -37, -31, 51, 68, -98, 79, -121, -44, -110, 50, 88, -82, -25, 62, 49, -50, -44, 122, 36, 121, -45, -108, 102, -35, -3, -128, -89, 82, 28, 11, -9, -19, 115, 58, 56, 98, -9, 58, -24, -12, 20, 69, 69, 41, 89, 1, 22, 1, -87, 114, 12, -37, 116, -59, -78, 3, 66, 19, -61, -50, 51, -40, 34, 113, 5, -12, -94, -111, -91, -105, -122, -126, -75, 71, 102, 110, -39, 23, 8, -41, -105, 3, 58, -49, -53, -77, 9, 23, 45, -30, 11, -1, 42, -84, 87, 106, 126, -111, -123, 109, 38, -104, 12, 63, -52, 91, -41, 118, 22, -107, -120, 95, 104, -107, -65, 31, 59, -91, 108, 61, 94, 110, 74, -22, -127, -20, -81, 80, 77, -70, -66, 114, 10, 32, -82, -122, 85, -77, -42, -25, 121, -36, -56, 27, 117, -42, -57, 59, 117, -110, -15, -58, -69, -68, 125, -12, 105, -24, -72, -93, -55, -9, -75, -97, -114, 119, 29, 12, 34, 90, -98, -87, -37, 127, 42, -70, -126, -71, 49, 36, 21, -126, -126, -35, -125, -102, -52, -24, -103, -86, -25, 104, -52, -58, -112, -64, 111, 37, -88, -77, -77, 28, -109, 42, 114, 17, -7, 81, -9, -96, 94, -115, 6, -92, -9, 39, -62, -24, -3, -89, 70, -74, -48, 63, 5, 62, 39, 52, -72, 0, -6, 110, 57, -67, 70, 82, -41, 68, 120, 99, -32, -48, 78, 90, -2, -112, -76, 116, -92, 7, -81, -113, -47, 86, -7, -19, -15, 124, -33, 109, 59, -24, 38, -100, -94, -21, -37, 65, -104, -103, -59, 48, 94, 30, 18, 14, 92, 98, 115, -66, -20, 78, 78, 46, -23, -28, -18, 12, -126, -79, 30, -11, -101, 109, -101, 82, 26, 82, -57, -17, 71, 110, 4, -72, 109, -4, -78, -101, 59, -123, 103, -46, -71, -45, -15, 117, 126, -53, 4, 98, 10, -2, 45, -62, -55, 114, 34, -118, -90, -109, 114, 121, -38, 15, 61, -124, 122, 37, 81, -102, -71, -12, -53, 82, -115, 113, -8, 69, 21, 89, -47, -105, -75, -50, -51, -103, 14, -4, -38, -29, 11, -97, 101, 116, -26, -85, 45, 75, -122, -114, 10, 105, -12, -81, 35, 25, 106, 127, 77, -75, 98, 121, 24, 45, -50, 29, -87, -61, -65, -52, -103, 57, -75, 124, -87, -45, -92, -126, 7, -114, -64, 24, -107, 109, -69, -19, 28, -6, -42, 108, 100, -38, -48, -126, 120, 33, -88, 88, -7, -51, 99, -69, -118, 127, 1, -80, -58, 90, 11, 9, 95, -92, -85, -2, 61, 115, -14, 116, 31, 33, 22, 87, 34, -52, -21, 44, 75, -29, 28, -31, 121, -64, 18, 90, -100, 104, -90, 105, 32, -3, -71, -45, 21, -12, 5, -101, 53, -109, 47, 124, 124, 64, 13, -121, 80, 23, -117, -83, 26, 88, 70, 111, -121, -101, 45, -63, 87, -125, 14, 74, 56, -57, -27, -116, -107, -78, -24, 101, -3, -62, 69, 72, 67, -28, 26, -74, -113, 89, 45, -40, 4, 127, -68, 56, 0, 15, 92, 115, -88, 102, -94, 115, 88, 123, 17, 123, 123, 113, -124, 28, -104, 92, -67, 61, -128, 17, -86, 25, 17, 70, -38, 11, -12, 61, 87, -75, -88, -34, -102, 113, -72, -38, 33, -80, -103, -33, 122, -1, 101, 28, -110, 53, -101, 48, 70, 26, -86, -7, -78, 4, 96, -68, 105, -49, 89, -115, 126, 3, -30, -19, -19, 94, 73, -69, -2, -16, -122, 120, 69, -68, 19, 21, 46, 69, 50, 105, 76, -107, -127, -83, 104, 9, 79, -1, 0, -83, 104, 35, 117, 37, -114, -66, 117, -94, 68, 95, -88, -123, -119, -101, -79, -52, 0, -125, 3, 62, 18, -50, 27, 58, -61, -91, -25, -31, -73, -26, 100, -93, 29, -21, -67, 1, 77, 73, 112, 116, -113, -104, -15, -114, -41, -118, -52, -98, 7, -88, -1, -99, -64, -15, 126, -97, -76, 106, 66, 23, 86, 30, 54, 72, -62, -61, 65, 55, 26, 109, -5, -122, -92, -52, -43, 106, -8, -67, 15, 91, 90, -72, -92, 117, 49, -72, 3, 29, 27, -78, 22, 33, 90, 23, 49, 63, -62, 0, 11, 105, -90, 124, 20, -45, -82, 43, 65, -31, -65, -65, 122, -32, 33, 11, 22, 96, -120, 39, 72, 83, 120, 33, 92, -73, -115, 62, 105, -108, 11, -7, 19, -87, 10, 102, 17, -87, 6, 18, 122, -72, -112, 45, -50, 14, -124, 113, -81, 31, 12, 37, -113, 88, -46, -27, -103, 88, -14, 66, 48, -96, 49, 72, -37, -66, -115, 114, 82, -36, -78, -63, 124, 73, -4, 117, -6, 23, -58, -56, 54, 37, 60, 35, -108, 73, 46, 42, -89, 69, -18, 82, 96, -40, 123, -43, -118, -35, -109, 62, 126, 121, 7, 47, 38, 98, 114, -106, 4, -125, -14, 72, 119, 64, -49, -49, 39, -101, -106, 21, 54, 68, -58, 30, -35, 86, 105, 19, 72, 82, 69, -52, -106, -104, 123, 11, -119, -63, -74, -33, -109, 124, -78, -128, -99, -21, 60, 76, 13, 59, 74, -19, 81, -93, -2, -37, 118, -57, -15, 51, 28, -68, -110, 4, -59, 49, 79, 78, 82, 112, 54, 42, -50, -77, -85, 24, -10, -95, 80, -118, -111, 7, 92, -121, 12, -52, -7, 82, -54, 33, -117, -83, 2, -120, 102, 99, -18, 68, -15, -77, -47, 63, 26, 36, -66, -77, 82, -53, 103, 58, 92, -18, -84, -67, 94, 110, 115, 53, -4, 5, -58, 28, -92, 97, 109, -102, 78, -34, -111, -2, 86, 29, -64, -64, 116, 82, -58, 11, 34, -74, 88, -2, -86, 83, -128, -102, 97, -64, 27, -109, -89, -45, 64, 47, -62, 2, 70, -85, -17, -59, 88, 65, -3, -26, -5, 19, -116, -11, -65, -15, -95, 119, 97, 0, -125, -84, 56, 104, -30, -111, 114, -122, 58, -42, 8, 53, 0, 88, 51, -119, 55, 115, 109, 28, 9, 124, 125, -77, -113, -43, 88, -2, 15, 12, 80, -81, 36, 11, -107, 117, 89, -126, -80, 18, 103, -3, 16, -79, 51, -124, 13, -1, -84, -3, -36, -123, 115, -34, -60, 67, -76, 35, 39, 37, 37, 95, 25, 119, 119, -67, 28, 52, 7, 55, -62, 17, -90, 112, 49, -30, 84, -71, -74, -9, -30, -57, 109, 82, 74, -114, -91, -30, -14, -30, 38, 39, -112, -101, 9, 10, 78, -49, 51, 126, 121, 55, -28, -81, 36, -78, 53, 14, -54, -110, -127, 47, -3, 10, 57, 121, -15, 16, -93, 64, -75, 68, -31, 29, -44, -117, -96, -33, 36, -98, 7, 39, -88, 75, 49, 73, -125, -69, -67, -73, 60, -30, 98, 65, 29, -113, -24, 12, -24, 90, 89, -84, 117, 113, 70, 124, -71, 65, -99, -71, 0, 32, 27, 20, 53, 25, 125, -19, -105, -61, 60, -82, 77, -93, -98, 89, 24, 39, -121, -101, -44, -18, 48, 27, -116, -116, 43, 67, 57, 79, 48, 32, 32, -44, -61, 2, 68, -71, -110, 9, -89, -68, -115, 15, -4, -86, 99, -72, -99, -71, 88, -16, 126, 70, -127, 43, -29, 114, 106, 12, -82, 103, 38, 9, -85, 119, 9, -64, 58, 64, 20, 99, -89, 123, 41, -121, 64, -64, 57, 108, -69, 24, -29, 14, 74, 34, -96, 21, -17, -12, -84, -51, 35, -107, -90, -12, 20, -81, -120, 117, 68, 91, 7, 60, 89, -32, -111, 16, -8, 51, 29, -110, -52, -121, 39, 95, -29, 9, -45, -82, 64, -34, 3, 41, -94, -69, -72, 76, -120, -54, -28, 90, 24, 100, -52, 27, 5, -36, -97, 6, 47, -68, 62, -19, 68, -69, -75, 108, -61, -56, 57, -82, -35, 27, -54, 109, 118, -82, 41, -68, -127, 54, -68, 87, -43, 46, -7, -7, -74, 106, -124, -28, 20, -88, 0, -54, -59, -60, 7, -4, -107, -109, -125, 21, 34, -26, 82, -116, -91, -74, -76, 41, 117, 23, -20, 85, -121, -69, -74, 31, -42, -45, 2, -101, 12, -58, -24, -104, 117, -27, 112, -54, -21, 92, -110, 41, 40, -3, -20, 111, -26, 57, 52, 43, -98, -83, 95, -16, 95, 9, -48, -77, -125, 39, -104, 26, -43, 53, -94, -35, -32, 82, 107, 20, 80, -99, 91, -92, -114, -100, 43, 9, 9, 5, 46, 60, -58, -50, -58, 3, 37, -10, -16, -13, 79, 90, 91, -70, -124, 31, 116, 115, 111, -50, 80, -29, 89, 39, 8, -72, 54, -59, 37, -128, -2, 40, -95, 61, 41, -17, -112, 64, -113, -54, -13, -109, -50, 0, -77, -98, -60, -100, 10, -5, -53, 103, 15, -128, -93, 64, 32, 52, -11, 57, 69, 11, -36, -48, -82, -104, 32, 44, -31, 24, 56, 2, -118, 86, 13, -123, 119, 100, 33, 77, 117, 91, 78, -84, 126, -82, 2, -38, -17, -8, -76, -89, -35, -91, 104, -38, 8, 112, 57, 46, -80, -15, -45, 113, -28, 3, -88, -20, -68, -64, -77, -44, 28, 77, 34, 57, 28, -78, 71, 91, 102, 88, -125, 8, -71, -81, 91, 104, -102, -59, 96, 112, -24, -114, 92, -2, 0, -116, -86, 104, 49, -64, -48, 19, 22, -56, -8, 40, 125, 38, 80, -1, -101, 97, -119, 76, 96, 60, -50, -37, -57, 86, 106, -85, -76, 16, -97, 29, -13, 61, 22, -32, -120, -51, 20, 88, -13, 109, 7, 47, 106, -82, 64, -18, 67, -102, 44, 78, 113, 33, 22, -121, 109, 86, -42, -128, -5, -23, -54, 106, 97, -11, -33, 45, 13, -48, 92, -111, -43, 11, -9, -65, 84, -8, 116, 52, -66, 14, 48, -114, 103, -43, -7, -97, 83, -71, -21, -33, -53, 100, 18, 76, 124, -84, -109, -99, 66, -37, -80, -112, -125, -115, 46, 92, -35, 119, -29, 100, 83, 20, 123, -22, 0, 81, 115, -82, -45, 65, 105, -53, -31, -94, -44, 49, -40, -125, -62, 37, -33, -51, 17, 33, -108, -28, 103, -70, -14, 25, -40, 80, 100, -31, -105, -116, -13, 54, -23, 88, 93, 1, 7, -14, 61, 28, 39, -93, -39, 85, 122, -84, -101, 53, -5, 22, -27, -84, 64, -6, -116, -46, -100, 124, -87, -88, 13, -81, 60, -71, 30, 56, 85, -50, 67, 36, 0, -30, -48, 13, -30, -47, 27, 4, -25, -37, -105, -115, -12, 108, -121, -26, -53, 28, 69, -65, -72, 54, 2, 6, -122, 72, 64, -93, 127, 107, -51, -85, -79, 102, -102, -33, -55, 110, 101, 49, 84, 112, 19, -95, 70, -128, 66, -2, -39, 50, -3, -120, 99, 125, -30, 12, 119, 7, -78, 14, -66, -48, -41, 21, -2, -95, 82, 116, -48, -29, -108, -122, -21, 77, -16, -8, 45, -37, -30, -102, 27, -46, -9, -72, -36, -126, 107, 39, 45, 37, 94, -29, -122, 106, 65, 109, -112, 58, -4, 2, 60, -68, -122, -45, 7, 14, -80, 58, -108, -68, -36, -39, 124, -107, 61, -126, 71, -94, 108, -121, -52, -30, -77, 126, 61, -54, -60, -54, -81, 96, 61, -53, -115, -122, 94, 126, -8, 72, 60, 117, -119, -77, 16, 76, -38, -79, 22, 111, 119, 3, -62, 60, -76, 21, -85, 121, -103, 23, 26, -54, 7, -4, -30, -45, 127, -42, -90, 113, 22, -105, 82, -118, 105, -43, 102, 89, -1, -4, 11, 89, -27, 117, 77, 70, -123, -94, -88, 62, -108, -14, 119, 115, -5, -22, 14, -85, 31, 3, 111, -32, 120, -37, -127, 14, -16, -44, 120, 8, -21, -2, -108, 90, -124, -41, -93, -79, -82, -124, -92, 56, -87, -109, 32, 79, -54, 112, 59, -41, -97, -128, 20, 118, -54, -72, 8, -63, 64, 29, 120, -34, 110, -74, -4, 39, 91, -78, 42, -9, 74, -95, 64, -93, -9, -104, -10, 64, 28, 77, 28, 62, -15, -15, -59, 18, 16, -127, -119, 77, 102, -45, 110, -89, -102, -83, 103, -85, -52, 42, 90, 48, -89, -68, 54, -3, -108, 53, -121, 105, 124, 94, 37, -98, -84, -53, 71, 26, 114, -85, -69, 124, 23, -105, -31, 25, -67, -113, 15, 52, -45, 63, 58, 45, 84, -102, -90, -26, -19, 3, -24, -119, -25, 86, 36, 80, 113, -84, -64, -125, -81, 6, -111, -8, 7, -23, -40, 15, -53, -106, -82, 114, -83, -27, -15, 60, -75, 41, -117, -78, 12, -115, 44, 95, 41, -118, 79, -23, 1, -54, -52, -92, -45, -28, -10, -82, 60, -83, 43, 16, -80, -68, -66, 73, 103, -65, 116, 17, -95, 8, 91, 51, -36, -19, -38, -86, 33, 96, 109, -116, 9, -85, -35, -70, -38, -24, 98, -101, -15, 63, 100, -127, -128, -51, 62, 16, -40, -13, 55, 24, 72, 112, -118, 116, 101, -69, 65, 86, -24, -37, -36, 52, 118, 28, -37, -10, 51, 38, -104, -51, 61, 115, 104, 51, 0, -70, 48, -108, 64, -73, 31, -39, 89, -102, -74, 54, -15, 61, -50, 38, 57, -10, -54, 124, 101, 92, -52, -5, 101, 26, -90, -94, -16, 12, -121, 52, -118, 125, 115, -37, 33, 92, -49, 8, 13, 109, -82, 92, 48, 84, 2, -1, 101, 72, 0, -92, -115, 85, -116, 11, 56, 27, 19, 124, 57, -64, -117, 69, -73, 23, 121, -113, 53, 37, -87, 118, -97, 43, -113, -41, -2, -37, 116, 64, -80, 93, -101, 29, 16, -3, -68, -3, 90, 113, -56, -74, -102, 45, 113, 98, -111, -88, -78, 63, -51, 83, -22, 72, -121, -109, 33, -30, 95, 20, -66, -30, 108, 89, 43, 52, -95, -111, -118, 87, -1, -19, 107, 74, 108, 70, -6, 10, 107, 49, 124, -36, 28, -67, -89, 76, -123, 60, 53, -23, -104, -125, 77, -16, 19, -49, -69, -56, -8, 78, 70, 5, -60, -30, 101, 90, 108, 32, -108, 123, -72, 121, -109, -35, -7, 14, -126, 99, 26, -67, -73, 5, -18, 123, 71, -73, 73, -84, -90, -56, 73, -106, 96, -89, 80, -122, 64, -115, 13, 52, -100, -49, 37, 28, 22, -27, -4, 119, 57, -102, -105, 69, 101, 55, 39, -60, -35, -25, -111, -69, -121, -41, 88, -35, -83, 98, -13, -40, -46, -46, 111, 43, -2, 85, 59, -101, 62, 105, -74, -1, 96, 6, -124, -98, 30, 114, 65, 67, 122, 114, 11, -64, -98, 73, 76, 97, -24, -12, 69, 125, 50, 111, 6, 44, -75, -9, 73, -12, 41, -95, -124, 45, -93, -23, 27, 47, 86, -6, 78, -73, -30, -3, -27, -119, -96, -53, 41, 67, 86, -72, 75, -103, 117, -22, -95, -71, -2, -40, 65, 67, 67, -18, -83, 70, 123, -8, -83, 25, 90, -95, -94, -37, -110, -85, -110, 94, 28, -47, 45, -69, 98, -33, 9, 53, -3, 84, -31, -29, -92, 38, 49, 88, -121, 78, 66, -91, 107, -125, -106, 97, -37, 63, 42, 44, -21, -27, 103, -76, -61, 95, -45, -108, -25, 7, -18, -30, 17, -86, -36, 13, -112, -21, -98, -112, -49, 35, 37, 82, -16, 93, 123, 84, -90, -125, -124, 24, 76, -35, 99, 108, -24, -59, 121, -97, 0, -41, 101, 104, -100, -19, -45, -79, 123, 25, 39, -120, -91, 121, -62, 46, -61, -57, -32, -96, -28, -125, 20, -91, -94, 74, -64, -107, -76, -108, 118, 60, -101, -36, 36, 40, 73, 50, -92, 68, -22, 15, 124, -13, 32, -113, 82, -16, -72, -21, 87, -4, 91, 127, 38, -84, -116, -111, 62, -77, 62, -79, -110, 40, -48, 0, 20, 106, 40, 5, 97, 127, 53, -17, 96, -7, 70, 27, 65, 28, 37, -122, -58, 13, 72, 118, 58, 106, -31, -97, 122, 44, 57, -93, 54, -35, -19, 70, 100, -76, -18, 33, 15, 73, 53, -109, 71, -110, -26, 30, 38, 57, -39, -44, 68, 17, 39, 117, 118, 1, 84, 37, 120, 40, -3, 96, 2, 6, 122, 7, -115, 122, 76, 82, -77, -18, 94, 127, 67, -28, -89, -126, -121, 40, 61, 21, 39, -72, 12, 99, -39, -81, 98, 70, -20, -86, 96, -88, -57, -96, -51, -38, 107, -17, 38, -60, -57, -44, -80, 45, -88, -88, 17, -119, 61, 79, -56, -108, -80, 18, 82, 61, -124, -37, -124, -75, 73, -30, 51, 106, 124, -120, 44, -88, 97, -20, 117, 75, -93, 91, -94, 80, 3, -92, 75, -1, 82, -31, 1, 93, 69, -4, 76, 47, -109, 90, 87, 52, -128, -93, -86, -36, 41, -56, 30, 23, -44, 12, 20, 120, 11, -60, 75, -95, 64, -90, 16, 73, 14, 12, 21, 126, 100, -119, 83, 56, 81, 6, 42, 72, -97, 78, 75, -50, -58, 29, 44, -51, -98, -52, 39, -58, -24, -71, -3, -21, -79, -109, 55, 26, 124, 108, -100, 11, -111, -45, 109, 73, 8, -44, -63, -24, 55, -64, -119, -55, 90, 122, -122, 125, -6, -86, -67, -67, -23, -20, -1, 122, 91, 108, 122, -73, -53, -69, 99, -59, 42, -1, 13, -57, 59, -95, 11, 91, 8, 48, -45, 30, 73, 10, -37, 37, -63, -32, 3, -52, -43, -88, 85, -114, -86, 36, -90, -127, 35, -49, -51, -56, -41, 120, -18, -62, -53, -69, 55, 72, -106, 18, 104, 127, -44, 27, 30, -1, -99, 72, 83, 91, 27, 15, -119, 77, -128, -105, 95, -67, 31, -69, -47, 1, -19, -28, -23, 90, 120, -103, -95, -90, -120, -22, 13, -6, 61, -47, 115, -84, -64, 39, -86, 118, 115, 77, 111, -71, -26, -83, 63, 35, 8, 81, -98, -81, -91, -23, 23, -123, -87, 76, -11, -122, -9, 42, 9, -22, 23, -86, 26, 86, 52, 2, 28, 108, -87, 25, -121, 23, -89, -99, -101, -82, 101, -92, -78, -15, -107, -59, 109, 98, -123, -37, 86, 83, 124, 56, 90, -77, -34, 83, -23, -54, -124, -56, -38, -102, 90, 127, 6, 118, 73, 102, -85, 44, -23, -38, 121, 127, 106, 92, 101, -61, 40, -87, 113, 71, -56, -104, 19, -105, 32, -57, -70, 83, -114, 58, -85, -112, 16, 38, 123, -75, 7, 115, -44, -89, 118, -96, -54, -97, -100, 104, -11, -122, 121, -120, 53, 57, -102, -49, -11, 22, -4, -19, -34, -38, 109, -60, 57, -92, -76, -70, -116, -89, 127, 30, -65, -11, -97, -111, -97, 25, 13, -41, 63, 1, 62, 20, -117, -3, 75, -108, -19, 103, 57, -50, -99, 5, -54, 24, -37, 63, -125, 13, -62, -80, -82, 96, -18, -115, -80, 57, -46, 23, 124, 52, 41, 89, 60, 74, -97, -76, 108, 94, -27, -42, -10, -98, 45, -118, -27, -17, -11, 102, -22, -124, 124, -83, -106, 14, 104, 104, -21, -110, -111, -57, 78, 34, 45, -71, -87, 75, -100, 104, 82, 84, -4, 127, 96, 45, 31, 51, -87, 67, -91, 20, -59, 15, 85, 56, -79, -90, -49, 109, -123, -65, -124, 117, 107, -35, -13, -34, 58, -42, -17, 122, 17, 16, -7, 19, 11, 123, 115, 5, -54, 49, -99, 31, 117, 119, -8, 55, 76, -53, -112, 91, -104, 112, 25, 82, -128, -74, -61, -41, 12, 75, -13, 49, -59, 113, 22, 125, -15, 119, -39, 108, -19, -126, 126, -29, -105, 77, -75, -80, 54, -7, 58, -62, -84, 25, -69, 58, 1, 100, 30, -46, 4, -34, 112, 111, 8, 9, 61, -61, -15, -64, 15, 33, 120, -25, 81, -36, 126, -52, -39, 112, 22, 88, 102, 107, 52, -96, 62, 124, -97, 79, -96, 95, -68, 1, 112, -83, 98, -11, 63, -49, -32, 72, -75, -115, -109, -45, 126, 73, 28, -102, 30, 89, 32, 91, -81, -86, 34, 29, 111, 19, -107, 109, 90, -66, 126, 68, 43, 38, 42, 95, 79, 90, 90, -13, -120, 119, 13, 35, -61, -11, -5, 36, -99, -98, -33, -99, -55, -62, 61, -59, -45, 86, -67, -29, 6, 28, 124, 14, -44, 6, -46, 41, 116, 109, 99, 49, -120, -72, -14, 31, -78, -10, 35, -94, 106, 69, -126, 14, -28, 26, 36, -62, -119, 66, -68, -92, -48, -9, -50, -24, -116, -47, 121, 3, -81, -69, -62, 63, 67, -36, 117, -41, 126, 37, 78, -10, 55, -36, -106, -40, -54, -69, -124, 1, 44, 112, 3, -59, -126, 73, -43, -121, 82, 62, 125, -37, -8, 14, 118, 43, -29, -56, -117, 79, 56, 54, 83, 10, -14, 100, -8, -98, -8, 116, 91, 101, -33, 42, 127, -88, -87, -106, 65, -34, 61, -91, 6, -106, -109, -21, -50, -106, -37, 94, -10, 38, -93, -66, 49, 50, 124, 103, 52, 37, -114, -73, 24, -96, -7, -121, 103, 62, -55, 54, -77, 75, 61, -18, -63, 80, -63, -32, 16, 58, -48, -57, -49, 2, 46, 28, 11, -75, 122, 20, -55, 67, 7, 116, 119, -43, 113, 119, 72, 95, -87, -34, 42, -39, 63, 23, -18, 27, -38, -78, 43, 99, -89, -68, -16, -104, 27, 109, 118, 106, 71, 70, 30, -19, -124, -78, -79, -76, -55, 2, -78, 36, -12, -101, 83, 17, -44, -110, 73, 61, -34, -127, 78, -40, 83, 18, 49, -36, -85, -110, -33, 27, 101, 89, 60, -110, -121, 8, 2, 41, -19, 123, 124, 114, -39, 18, 88, 53, -29, -69, -32, 8, -5, 19, -74, 48, 11, 126, 71, -116, -23, -72, 87, 22, 48, -4, -102, -109, 123, -49, -76, 89, -108, 51, -78, 70, 25, 39, -109, 65, -104, -69, 88, 0, -50, 90, 15, 84, -99, 49, -106, -20, -117, 100, 100, -49, 50, -119, 108, -36, 31, 49, -105, 24, -48, -68, 123, 83, -28, 114, -44, -77, -13, 119, 17, -32, -82, 35, -124, -11, 93, -27, 111, 121, 23, -5, -15, 56, -74, 34, 120, -66, -38, 44, -124, 18, -100, -83, -107, 56, 89, 101, 2, 87, 16, 53, 53, -89, 37, -81, -14, -114, 120, 16, -121, 9, -34, -123, 52, 53, -105, -30, 32, -114, -42, -19, 121, 59, -94, 123, 58, -106, 67, -34, -30, 69, 52, -19, -75, 85, -95, -66, -96, 75, -79, -23, -15, 57, -20, -65, -65, -60, 113, -88, -66, 12, 123, 68, -31, 4, -23, 82, 102, 112, 65, 84, 109, 101, -75, -95, -28, 127, 56, -112, 2, -113, 89, -100, 70, 58, -76, -41, 68, -78, 56, -82, -29, 15, 12, 78, 101, 2, -57, -88, 5, 116, -63, -58, 126, -106, -127, 53, -91, -107, 37, -125, -112, -111, 48, 103, 48, 48, -90, -2, -8, -21, -87, -14, 13, -50, -90, -95, -126, -28, -28, -47, 43, -113, 108, -49, 76, -43, 94, 21, 104, 25, 60, -104, -23, 50, 36, 116, 45, -2, -92, -78, 127, -25, 65, 36, -13, -112, 32, -20, 59, 47, -33, 35, 28, 54, 81, -102, -10, 64, -14, 38, -27, -36, 40, -41, -32, -78, -6, 119, -97, -90, 97, 60, -96, -7, 114, -121, -8, -89, 85, 81, -104, -71, -85, -57, 18, -62, -25, -69, -116, -104, -73, -34, -11, -45, -56, -33, 68, -10, 63, 24, -40, 120, -68, -57, -45, -15, -63, -58, -69, -8, -107, 24, 63, -79, 47, 30, -101, -36, 83, 88, -35, 61, 29, -49, 111, 39, 51, 75, -59, -113, 111, -88, -81, 53, 24, 35, -94, -71, -72, 12, 48, -104, -67, -113, 17, -18, 14, 26, -115, -117, -10, -63, -78, 82, -89, -4, 76, 104, -16, 39, -51, -86, 37, -6, 117, -88, -56, -61, 110, -25, 6, 0, -124, 124, -40, -84, -52, -110, 63, 18, 47, -58, 95, -119, 118, 62, 91, -53, -107, -13, 56, 8, 110, -123, -16, 54, -84, -36, -37, 9, -57, 84, -23, 40, -25, -26, 37, -91, -120, -99, -46, -22, -21, 108, 45, -84, 119, 36, 89, -62, 1, 116, -91, -102, -22, -39, 4, 10, -48, 37, 86, 100, 13, 25, 95, -62, -99, 18, -119, 6, -68, 4, -88, 40, 106, -44, -35, -105, 21, -55, 7, -119, -70, 108, -43, 110, 75, -65, -70, 127, -97, 115, -69, 124, 107, -105, -33, -60, -45, 102, 7, 119, -11, -2, 102, 65, -16, 8, 112, 61, -2, -1, 64, 56, 91, 36, 70, 123, -48, 76, 12, -113, 43, -6, 27, -16, 56, 122, -16, -27, 116, 54, -12, -124, -26, 112, 17, 105, -58, 40, -41, -105, -128, -80, 27, 111, -28, -79, -109, -92, -31, -73, 81, 11, -30, 63, 111, -94, -4, -64, -48, 78, 36, 45, 64, 52, 119, -74, -16, -117, -85, -55, 113, 49, -21, 37, 57, 96, -30, -50, 9, -40, 65, -103, -94, -42, 48, -2, -67, 52, -21, -105, 64, 12, -40, 22, -122, -61, 33, 87, 99, -101, 94, -4, 22, -2, 2, -20, 59, -88, 34, -51, 6, -94, -114, -100, -21, 75, -86, 91, -60, -112, -113, -45, -29, -94, -38, 45, 113, -13, -30, 38, 1, 31, -84, -53, 42, -101, 78, -4, -2, 98, -105, 60, -50, -73, 69, 117, -51, 116, 76, -70, 59, 90, -115, -1, 20, -65, -38, -10, -128, 31, -16, -20, 41, -17, 58, 88, 119, 3, -119, -106, 83, -109, 127, 92, 24, -24, 110, 42, -114, 15, -54, -77, 43, 72, -55, 126, -64, 5, 15, 104, 61, -62, 115, 127, -93, -83, -116, 79, -127, 40, 7, 69, 79, 60, -59, -83, 14, -127, 68, 30, -64, 45, -40, -22, 34, 14, -44, -7, 107, -89, 100, 13, 72, -20, -123, 49, 102, -69, 116, -34, -110, -77, 105, 89, 101, -98, -16, 43, -94, 57, -75, 31, -77, 8, -70, 65, 72, -29, -37, 99, 29, 5, 4, 65, 112, 34, 46, 122, 94, -94, -56, 72, 75, -29, -24, 94, -57, 36, -78, 93, -21, 45, 84, -31, -40, -86, -117, -101, -64, -10, 14, -122, 103, 11, 70, 99, -75, 87, -126, -41, -17, -55, -15, -76, 91, 82, -60, -49, -42, 61, -46, 115, -57, -52, -51, 62, 45, -10, -28, -58, -78, -7, 88, -41, 101, -37, 16, 61, 54, -9, 103, -101, -36, 127, 126, 105, -52, 4, -119, 62, -73, -92, 55, 81, -58, 13, -119, 102, -33, 75, -26, -108, -18, 7, 74, -69, 102, 18, -96, 103, -102, 66, 30, -24, -55, 121, -115, -50, 43, -76, -79, -89, 18, 123, -72, -64, -119, 38, -71, 110, -102, 58, 108, -73, -40, -72, -74, -17, -34, -7, 82, -52, -89, -89, 109, 124, -52, 60, -7, 49, -17, 60, 107, 40, 9, 46, 57, -118, -112, 52, 89, -108, 96, -48, -15, 83, -92, -82, -31, -49, 106, 60, 114, -71, -83, 102, 46, 13, 82, 78, 15, 13, -122, -66, -88, -103, 9, 95, -21, -86, 85, -77, 83, -123, -36, 116, 60, -57, -118, -68, -37, -52, -70, -110, -112, 12, -95, -55, 97, -75, 105, -124, 103, 96, -43, 63, 38, -110, 15, -39, -33, 40, 10, -116, -81, 20, -68, 73, 23, -32, 83, 122, -56, 30, -108, 38, -103, -7, 34, 97, 53, -83, -4, -43, 50, 92, 104, 17, 106, -26, 52, -115, 81, 79, 87, 105, 59, 62, 110, 30, -104, 42, 124, -18, -86, 56, 125, -16, -52, -78, -128, 6, 16, 44, -74, -47, 20, -22, -1, 49, -53, -120, 63, 47, -12, 40, -107, -98, 90, -74, 20, -24, 91, -41, 88, 109, 77, -76, -48, 43, -35, 61, -68, 124, 18, -71, -118, 44, 111, 19, 40, -41, 117, 40, 8, -43, -104, 120, 26, -34, 103, 112, 42, -60, 86, 88, 14, -4, -84, 118, 40, -24, -66, -2, -47, -23, -44, 111, 86, 75, 111, -39, 32, 70, -62, 2, -4, 17, -59, 35, -79, -64, 41, 99, 124, 61, -102, -71, -76, 29, 90, -30, 59, 18, -39, -89, -67, -79, -116, -16, -76, 74, -51, 97, -70, -98, -10, 50, 95, 69, -128, -80, 94, 28, -78, -47, -18, -73, 124, 117, -96, -48, 100, 59, 46, 30, -11, -87, 63, -48, 125, -97, -46, -38, -38, -79, -111, -115, 25, 125, 60, -20, -39, -106, 84, 65, 47, 127, -13, -23, 6, 72, 108, 96, 25, -128, -98, 42, 30, -82, -25, -95, 55, 88, -6, 15, -80, 42, 25, -87, 81, 63, -85, 5, 56, -44, 4, -74, -116, 114, -36, -101, -39, -66, 63, -126, 23, 13, -45, 96, -2, -114, 50, -90, 98, -24, 71, -19, -110, -33, -32, -60, 125, -102, 123, -20, -79, 118, -10, 1, -109, -119, 109, 43, -16, -56, -10, -69, -38, -71, -34, -126, -111, -53, -43, 26, 1, -69, 115, -40, -108, -11, 63, 14, -24, -100, 84, 29, -120, 37, 35, -38, -67, 124, 49, 76, 31, 78, 57, -44, 73, 0, -94, -28, 9, -86, -91, 74, 79, -120, -108, -102, -69, 64, 3, -104, 92, -70, -59, -109, 76, -32, -87, -30, 67, -31, 86, -105, 5, -21, -112, 104, 74, -111, 5, 121, 3, -4, -13, 30, 7, -12, -65, 4, -107, -104, -98, 107, 55, -69, -96, 49, 83, -12, 69, 45, 112, 1, -49, -48, -39, -13, -77, 57, -85, 81, -12, -36, 97, -124, 85, 90, 98, -128, -23, 95, 107, 46, 28, 123, -98, -72, -64, -40, 7, -50, 41, -122, -99, 87, 126, -125, -4, 2, 66, 14, 56, 19, 53, -31, 55, -98, 13, 100, -69, 85, 0, 14, 116, -50, -13, 72, 11, 43, 90, -90, 84, -115, -49, -83, -89, -1, 111, 86, 73, 117, 53, 92, 77, 46, -51, -74, -125, 4, -38, 93, 56, -47, -80, -5, 77, 91, -81, -119, 59, 56, -41, -26, -108, 55, -58, 57, 20, 119, -32, -95, -118, -48, -102, -97, 45, 65, -110, 20, 80, 107, 47, -77, 16, 18, -70, -102, 23, -19, -99, -32, 115, 90, -72, -84, 24, 73, 43, -98, 41, 77, -1, 52, 66, 42, 0, 85, -40, -108, 16, -5, -1, 17, -65, 65, 97, 95, -30, -20, -13, 38, -65, -29, -39, 61, -45, 43, 2, 97, -62, 112, -64, 118, 107, 16, -79, 1, 41, 39, 20, 7, 103, -44, 115, -43, 36, -118, 38, -66, 32, -73, -38, -18, 69, -23, 28, -38, 91, 67, -32, -95, 48, -7, 18, 93, 40, -14, -13, -108, -21, 53, 57, -23, -123, -44, 73, 60, -13, -83, 47, 51, -96, 89, 50, -106, -40, -86, -98, 116, 107, -56, 35, -7, 91, 24, 10, -25, -29, 57, 55, 105, 90, 32, 72, -70, -83, 13, -59, 120, 121, 66, -10, -64, 79, 79, 28, -44, -108, -28, -30, -31, 98, -48, -21, -26, -35, 37, 76, -98, -111, 36, -11, -14, 78, -38, 93, 77, 92, -120, -24, -101, -123, 29, 44, 77, -57, -43, -26, -97, -81, -54, -67, -31, 85, 9, -18, -74, -58, -73, -77, -127, 89, 8, -99, -66, -86, -21, -85, -100, 5, -109, 13, -50, -9, 99, -27, 125, 58, 71, 66, -20, 109, -103, -85, 67, -7, -110, -46, 18, -44, -88, -115, -104, -12, -11, 85, 6, -7, -2, 78, -118, -102, -47, 22, -85, -39, 117, 10, 12, -97, 71, 123, 111, 4, -91, -30, -14, 50, 14, 12, -83, 8, -69, -115, 14, 119, -23, -128, 97, 6, -40, -6, -59, -126, 70, 82, 119, -38, -64, 20, 31, -42, 73, -44, -96, 98, 60, -85, -39, -24, -33, 26, -43, -54, 111, 122, 35, -86, 58, 123, -98, 56, 12, -98, 127, 115, -115, 72, 7, -121, 50, -46, -25, -30, 30, 76, 117, 48, -60, 74, 2, -97, -71, -60, -47, 41, 46, 97, 71, -67, -102, 101, 112, 71, 53, -2, 60, 91, -18, -79, 36, 31, -17, 39, -48, -91, -15, -91, -90, -107, 87, 126, 45, 13, -112, -72, -78, -40, 43, 8, -77, -81, 11, -89, 99, 23, -106, 77, 89, 120, -122, 1, 104, 75, 1, -6, 70, 39, -83, 79, 42, -62, -86, -47, 120, -67, 115, -22, 83, -124, 53, 91, 31, -62, -74, -4, -10, -90, 0, -76, 15, -35, 87, 11, 74, -67, -16, 127, -80, -57, -69, -99, 5, 15, -123, -45, 40, 105, 10, -13, 114, 117, 24, 37, 2, 111, 107, 102, -52, 51, -23, 34, 6, -90, -54, -96, -16, 104, -66, -22, 70, -125, 104, 62, 94, -5, 0, 70, -71, 104, -122, -66, -101, 50, -114, -54, 23, 86, 124, 45, -28, 44, -60, -87, 60, -61, -44, 43, -80, -60, 49, 11, -59, -21, -6, 79, 24, 29, -82, -32, -35, 87, 36, -82, -86, 4, 77, 82, -93, 35, -13, 71, -63, -35, 53, 36, -80, -125, -8, -84, -126, -81, 45, -100, 30, 58, 67, 72, -105, -54, 126, 54, 56, 4, 69, -16, -14, 4, -126, -68, -58, -25, -23, 65, 34, 79, 123, -75, -111, 7, -106, 57, 124, -26, -62, 124, -126, 10, -69, 13, -18, -22, 73, 66, -99, -86, 54, -9, 50, 118, 50, 114, 123, -32, 68, 2, 36, 38, 60, 79, 75, 75, -17, 115, -57, -65, 93, 109, -80, -75, 127, 86, 67, -20, -91, 72, -82, 24, -95, 105, 109, 25, -19, 111, 87, 82, 90, 117, 49, 58, 29, -59, 100, 5, -63, -122, -115, 1, 74, 17, -23, -118, -4, -93, -12, -18, 13, 116, -91, 14, -3, 100, 2, -90, -20, 79, 32, 35, 10, 110, 63, -94, 77, 63, 127, -20, 122, 70, -96, 43, 105, -3, -115, 116, -78, 120, -123, 109, -126, -111, 13, -49, -35, -70, 19, -13, 70, -49, -17, 61, -112, 42, 24, 4, 21, -28, 26, -77, -31, -104, 73, -1, -58, -49, 30, 125, -87, -69, -109, -83, 112, 48, 10, 64, 79, -62, -25, -5, -37, 0, 11, -25, -40, 47, 11, -24, -115, 48, 82, -112, 16, -48, -42, 18, 9, -74, -53, -20, -107, -43, 85, -58, 29, -85, 20, -121, -78, -90, -92, 47, 21, 34, -113, -68, -59, 103, 5, 30, -50, 61, -89, -39, 5, 118, 86, -43, 97, 9, -47, -41, -124, 81, -16, 79, 53, 43, 9, 113, -81, -55, -28, 66, 31, -82, 105, -2, 117, 21, -70, -113, 20, 11, 17, 88, 88, 37, -71, -122, 109, 15, -57, 99, 122, -65, -109, 18, -109, 90, -1, -94, -69, -37, 25, -113, 125, 11, -6, -125, 29, -124, -83, -30, -56, -89, 10, -10, 37, 112, 80, 1, -11, 4, 35, 80, 68, -82, -7, 87, 21, 57, -17, 71, 18, 103, -118, -109, -19, 5, 13, -119, -46, -40, 38, 1, -101, -37, 22, 19, 94, -29, -16, -68, 23, 76, -119, -46, -34, 1, 113, -26, -13, -79, -35, 19, -25, 81, -69, -123, -49, -7, -59, -111, -43, 49, -47, -88, 67, -100, 43, -86, -59, -5, 33, 92, 22, 9, -92, -46, -113, -12, 51, 61, 115, -41, 19, 15, 70, -12, -104, -35, 66, 79, -67, 24, 54, 72, -93, -16, -34, 57, 89, -120, -88, -60, 80, 36, 78, -89, 5, 51, 9, -50, -3, -18, -17, 8, -66, 23, 60, 126, -49, -53, -33, -89, -17, -53, 37, 94, -81, 2, 0, 25, 69, 75, -121, -18, 68, 88, 7, 37, -36, -107, 39, 102, 47, -103, -122, 15, 34, -58, -110, -103, -49, 94, -69, 48, -9, 26, 4, 127, 35, -53, -113, 114, -21, 15, 101, 69, 45, -127, -53, 122, -10, 38, -17, -79, 106, -80, 4, -52, -86, 45, -52, -10, 89, -37, 98, -70, 123, -57, -56, 116, 0, -66, -27, -69, 89, -128, 25, -106, -51, 52, -68, -92, 48, -128, 35, 37, 118, 124, -94, 85, 24, -29, 78, 69, 64, 33, 78, 77, 18, -11, 74, -35, -73, 10, 42, -13, -35, -6, 27, -30, 116, -45, 12, -8, -117, 19, 125, 32, 111, -35, -35, -111, 17, 13, -103, -93, 52, 38, 28, 105, 99, -68, -13, -115, -94, 76, -76, 2, -64, 81, 80, 86, 48, -6, -78, 13, -79, 44, -31, 59, 85, 21, 54, 117, 58, 31, -119, -43, -76, 72, -121, -55, -90, -18, -112, 37, -29, 75, 43, 55, -128, -74, 54, 116, 121, 98, 25, 49, 5, 42, -47, -1, 32, 14, -75, 17, 72, -19, -111, -79, 44, 110, -4, 85, 99, 41, 85, -112, -40, 73, -106, -123, -44, -64, -54, -22, -83, -27, 98, -33, -127, -118, 34, 31, -104, 7, -78, -50, 107, 9, -64, 23, 126, 83, 72, -77, 67, -52, 46, 68, 64, -60, -32, -14, -83, -29, -43, -71, 97, 122, -96, 86, 88, -20, 90, 33, -47, -23, 95, -123, -1, -42, 84, -64, 126, 108, 37, 72, -32, 9, 29, -82, 124, 124, -80, -73, -35, 34, 28, -36, -70, -45, -99, 69, 110, -33, -101, -105, -109, 34, 100, 114, 72, 1, 21, -52, 51, 17, 38, 24, 55, -76, -51, 39, -104, 88, 107, 10, 22, 72, 60, 42, -88, 48, -120, -2, -92, 2, -98, 58, 116, 29, -14, -88, 55, 49, 79, -9, -70, 120, 123, 1, 19, -94, -125, -117, -6, -113, 57, -109, -18, -62, 123, -108, -118, -12, -21, -26, 63, 84, -15, -7, -83, -18, -37, -127, -29, -58, 29, -25, -20, 38, 83, -83, 99, 17, 4, 115, 19, -47, 93, -36, -76, -61, 98, 51, -22, 50, 41, 37, 83, -126, -59, 90, 54, -25, 91, 106, 107, -74, -72, -123, -18, 88, -47, -99, -121, 26, -86, -106, -110, -14, -117, -66, 102, 82, 36, -12, -14, 51, -80, 41, 89, -83, 8, 52, -55, 100, -116, -6, 70, -92, -44, -39, -62, 122, -112, 91, 100, -20, 124, -84, -22, 59, 125, -58, 108, -32, -9, -68, -81, 102, -109, -63, 84, 47, 99, -78, -14, 84, 1, 36, -114, -29, 13, -2, -4, 4, -128, 72, 2, 119, 81, 120, 1, -90, 46, 53, 115, -38, -54, 69, -111, -47, 112, -111, 104, 26, 47, 62, 92, -8, 92, -47, 9, 2, -2, -13, -32, 76, 88, 15, 74, -51, -106, 12, -64, -33, 52, 35, -66, 120, -63, 79, 56, -105, 100, 27, -118, -42, -66, 23, -46, -100, 100, 14, -19, 121, 53, -83, 31, 6, -119, -84, -43, -128, 55, 55, 93, -56, -31, 59, 71, 37, -39, 117, 13, 78, 76, -113, -101, 19, 105, -35, 79, -85, 63, 127, 127, -121, 93, -122, -66, -49, -27, -4, 85, -26, 1, -14, 1, 73, -63, 55, -82, -87, 94, -96, -37, 47, -58, 33, -17, 10, 19, -76, 106, 111, 36, 103, 2, -65, -97, -70, -29, -60, -22, -115, 71, 78, 114, 124, -14, -54, -74, 39, 22, -110, 22, -48, 65, -78, -88, 120, 67, 72, -42, 9, -83, 13, 44, -81, 110, 98, 81, 28, -74, -41, 101, -17, 36, -93, 40, -94, 74, 98, -73, -103, -32, -123, -39, -49, 71, 26, 40, 54, -7, 104, 100, -117, 43, 15, -100, -41, -95, 15, 52, 44, -72, 46, -125, 56, 106, -82, -34, 37, 79, -117, 1, -93, -76, 75, -56, -119, -19, -99, -126, 70, -72, -43, -85, -17, -37, 14, -119, 110, 43, -14, -59, 90, 68, 111, -40, 45, 80, 99, 93, 75, 70, -74, 8, 12, -101, -65, 36, 74, -103, -41, -3, -74, 32, 62, -10, 81, 86, -54, -8, -106, -92, 109, -108, -31, -116, -17, -85, 74, 10, -9, -103, -86, -5, 110, 68, -63, -29, -85, 0, 106, 119, -107, -14, 20, 80, 109, 69, 106, 127, 52, -55, -12, 31, -106, -70, 0, -79, -10, -38, -105, -63, -94, -127, 82, -35, -11, 71, -86, -78, 81, -79, 68, 32, 61, 1, -107, -93, 26, -38, 127, 87, -82, -119, 94, 27, -86, 38, 49, -8, 62, -78, 76, 38, 71, -15, 55, 71, 18, -69, 14, -15, 127, 81, -117, 68, 73, 38, -18, 29, -40, -17, -68, 73, 12, -42, 27, -44, 4, -126, -14, -92, -60, 19, 2, -33, 22, 2, -81, 72, 17, -45, 78, -113, 60, 56, 87, -119, -64, 60, 80, 95, -89, -42, 99, -32, -29, 0, -7, 40, 48, -66, -78, -118, -112, -95, -62, 78, 96, -65, 61, -48, -91, -108, 18, -79, -65, 41, -26, 93, 112, 121, -20, 5, -21, -71, -125, -25, 19, 115, 9, 112, -125, -54, 62, -117, 38, -113, -25, 89, -50, -97, 70, 100, 109, -118, -57, 59, 21, 59, -125, -115, -7, 54, -100, 98, 82, -90, 94, 47, 2, 125, 24, 55, 34, -102, -51, 75, -94, -46, -27, -44, -43, -41, -121, -17, -32, -10, 68, 75, -8, -53, -36, -107, -13, -78, -36, -56, 1, 53, -100, -89, 39, 89, -1, -60, 115, -127, -75, -124, 65, 94, 47, -28, -121, -21, 92, 109, -64, 91, 99, -22, -22, 122, -91, -34, 114, 100, -113, 6, 120, 79, -10, -84, 102, 1, 52, 69, 114, 17, -28, -107, 126, 114, -77, 99, -82, 41, -22, 124, 7, 51, 14, -45, -85, -103, 95, -27, -77, 55, 17, 103, -114, -103, 115, 52, 67, -10, -83, -114, 11, 9, -17, 96, 50, 105, 5, -38, 100, -37, 85, 71, -79, 54, 92, -103, -102, -18, 3, 16, -105, -95, 115, -119, -99, -20, -85, 67, -58, 74, 46, -112, 74, 115, 1, -32, -70, -120, 85, -68, 20, -71, -42, -30, 114, -88, -117, -40, 103, -10, 72, -7, -3, 13, 97, 3, -50, -66, 57, -64, 40, 14, -62, -95, 108, -5, -106, -73, -48, -34, 65, -38, -45, 100, -42, -26, 44, 120, -89, 78, -101, 75, -46, -108, -81, -39, -31, 62, -15, 68, -94, -126, 84, 16, 28, 82, 81, 61, 37, 39, -80, -49, -104, -70, 75, -48, -104, 68, -47, 125, -17, 83, 23, 73, 59, 106, 52, -111, 124, -91, 75, -41, -67, -120, 116, 107, -1, -55, 45, -16, -102, 2, 42, 114, 13, 60, -2, -56, -65, 40, -29, 29, -70, 7, 104, -112, -47, 41, -22, -4, -79, -4, -49, 81, -7, 122, 44, 20, -98, 53, 104, 14, -14, 73, -128, -96, 98, -117, -125, -118, -24, -88, 19, 106, 77, 32, -116, 66, -86, 35, 125, 39, 35, 85, -1, -84, -87, 101, -84, 70, -27, 49, -30, -21, -74, 2, 93, 8, -116, 38, -86, 62, 60, 48, 93, -117, -123, 65, 8, -17, 43, 93, 62, -84, -7, 54, 106, -121, 84, -24, -101, -86, -74, 121, -17, -6, -75, 63, -8, 97, 101, -19, -5, 8, 90, -2, -4, -124, 58, 2, -48, 66, 4, -100, -13, 81, 43, -101, -50, 23, 64, -75, -85, 6, 11, 9, 117, -44, -74, -62, 47, -89, -117, 45, 84, -66, 16, 11, 31, 49, 40, -65, -55, 38, -45, -110, 3, -44, -93, 71, 5, -126, 62, 108, 6, -61, -50, 42, 122, 26, -4, -18, 88, -104, -38, -48, -19, 3, 90, 32, 119, 58, 33, 31, -76, 1, 15, 121, 27, -91, -28, -57, 76, 14, 30, 92, 112, 46, -113, -121, 116, -79, -26, -55, 58, 126, -113, 94, 68, -98, 83, 2, 37, 72, -73, -87, -22, 50, 89, -25, 61, 24, 95, 73, -14, 49, 124, -23, -17, 85, -55, -88, 58, -70, -88, 86, 70, 113, -93, -27, -75, 98, -69, 38, 16, 106, 22, -84, 47, -21, -101, 47, -125, -13, 82, 45, -11, 9, -116, -55, -96, 29, 24, -17, 88, 117, -74, 45, 15, 61, -73, 123, -88, 119, -43, 16, -87, 9, -22, 10, 102, -105, -106, 46, -37, -20, -30, 87, 109, -112, 51, -38, -117, -37, 92, -34, -75, -104, -20, 42, 70, -120, -95, -45, -69, 87, 5, -3, -95, -86, 84, -5, -14, 75, -74, 58, -10, -92, 57, 21, -30, -7, 87, -76, 12, -90, -90, -6, -25, -3, -113, 100, 24, -23, 92, -109, -100, 125, 31, -52, -50, -41, 57, -91, 119, -105, -10, -99, -84, 3, -97, 41, -36, 100, 21, 2, 24, 88, 99, -8, 123, -62, 63, -115, 95, 122, 10, -13, 0, -22, -4, -106, -109, -75, -28, -92, 95, 116, 10, -118, -20, -37, -80, 106, 116, -37, -43, 57, -81, -72, 8, -94, -47, 95, -1, 70, -119, -50, -90, 44, 44, 21, 127, -65, -66, 59, 1, 111, -127, -89, 96, -99, -92, 14, -99, 17, 31, -113, 109, -101, 111, -38, 55, -72, 50, 18, -82, -25, -6, -110, 26, -124, 34, 63, -98, 27, 14, 17, 30, 120, -64, 114, -66, 126, 38, 4, 50, 39, -109, 77, 88, -111, 86, -125, 62, -54, 107, -115, -112, -65, -103, -20, 82, -45, -3, 123, 4, -36, 24, 88, -33, -83, -34, -81, 88, 121, 110, -125, 38, 125, -58, 77, -40, -4, -21, -67, 78, -114, 66, -77, -70, 1, -57, 117, 126, -83, 103, -75, -84, 77, -80, 34, -36, -43, -58, 64, -86, 80, -30, -105, 69, -11, -80, -25, 5, -70, 48, -38, -41, -59, 77, -118, -88, 9, 111, -76, -49, 42, 36, -84, -128, 5, -37, 37, 118, -100, -79, -77, -5, -44, -10, -69, 106, -71, 126, -79, -74, -48, -23, -76, 37, -23, 61, 74, 31, 64, -21, 15, -86, 30, -24, 62, 36, -99, 40, -119, -128, 62, 1, 51, -23, -43, 25, 108, -23, 126, -32, 90, 59, 49, 118, 96, -93, 86, -114, -5, -26, 71, 7, 36, 5, -35, -14, -78, -20, -124, 84, 41, -125, -126, -63, 127, 106, -45, 74, 24, -49, -77, 57, -79, 126, 57, 92, -110, 123, -84, 41, -38, 42, -117, 67, 115, 23, -61, -23, -121, 103, 29, -48, 34, 36, 94, -70, -10, 52, -48, -53, 70, 11, 6, -99, 65, 123, -35, 41, -109, -95, 17, -40, -117, 119, 113, 95, 5, 45, -32, 83, 79, 116, 41, -26, -102, -127, 122, -9, -16, -119, 21, -56, 72, 19, -34, -93, -58, -88, -106, 41, -34, -1, -77, -101, 24, 17, 40, -48, -62, -46, 14, -56, -92, 80, 26, -85, -86, 78, -56, -38, -86, 50, 11, -59, 53, 42, -73, 122, 7, 86, -27, -61, -71, -110, 92, 55, 79, 8, 101, -8, -26, 40, -32, 50, -49, 23, 106, -49, -26, 11, -45, 126, 35, -93, 59, -115, 53, -123, -8, 37, -26, -21, -12, -122, 90, 104, -24, -75, 17, -93, -119, -10, 106, 66, -41, 51, 19, -11, 95, -35, -27, -40, 82, -48, -26, 36, -80, -80, -53, -27, -59, 15, 85, -48, 10, 0, 2, 111, -107, 127, 11, 40, -32, -120, -115, 28, 92, 21, -53, -11, 14, 49, 39, 114, -50, -43, 122, -68, 27, 23, 19, -53, 34, 87, 13, -83, -50, -42, -63, 35, -79, 91, -122, -82, 4, 16, 94, 92, -8, -105, 28, 32, 112, -121, -75, -73, -16, -127, 19, -85, -31, -3, -32, 123, 39, -125, 101, 61, 25, -124, -83, 94, -36, -107, 106, -119, -5, 1, 118, -53, 84, -29, 113, 39, 40, 5, -121, -121, 57, 119, -55, -125, 46, 2, 124, -60, 92, -71, -82, 34, -109, -93, -68, 90, -53, -72, 76, 104, -109, 9, 108, -18, 59, 20, -127, 90, -17, 90, -127, -31, -107, 61, -32, 47, 42, -38, 23, 88, -12, 124, -66, -12, 123, -14, 26, -37, 84, 45, -64, 118, -81, 90, 62, 91, -39, -8, 12, -109, 24, -39, -24, 83, -59, -45, 94, 15, -117, -45, -125, -121, 57, 87, 87, 125, -43, -52, -18, -49, -97, 119, -36, -120, -102, 93, 95, -100, 70, -7, 102, 102, 57, 75, 28, 35, -127, 36, 12, -37, 43, 20, -122, -9, 90, -61, -125, -7, -42, -36, 53, 21, 85, 78, -111, 45, -125, 2, 63, -16, 111, -68, 26, -9, -4, -45, -96, 5, -119, 109, 12, 34, -15, 115, 19, 25, 125, -56, 17, -62, -94, 52, -126, 2, -47, 14, -58, -91, 126, 27, -44, 26, -80, -91, 26, 36, -70, 33, -44, 89, -60, -90, -106, -11, -63, -117, 68, -14, 98, 34, 5, -125, -19, -123, 50, -99, 92, 48, -115, -73, 99, -5, -6, -82, 60, -99, 93, -45, -1, 47, -66, 109, -101, 89, 63, -97, -56, 49, -119, 108, 95, 119, 3, -81, 74, -61, 98, 43, -115, 67, 111, 44, -105, -58, 74, -47, 120, -34, 48, -79, 17, 68, -4, -93, -13, -17, 10, -120, -121, 21, 46, 66, -97, 44, 35, -106, 105, 33, -73, 75, 120, 74, -50, -56, -43, -84, -82, 122, -48, 44, 101, -97, 81, 72, -46, -95, 15, 66, -80, 83, 123, 11, 120, 14, -4, -26, -37, -56, -53, 30, 63, -7, -81, 103, -58, -74, 77, -87, 96, 18, -119, -60, 12, 4, -32, 34, 4, -57, -17, 109, -15, -127, -112, 6, -54, 70, 15, 67, -103, 101, -80, 41, -86, -91, 67, 3, -6, 61, -116, -44, 88, 99, -91, -68, 90, 87, -16, -58, -47, -125, 15, -60, 26, -94, 111, 73, -31, -77, -77, -89, 11, 55, 16, 100, -25, -94, -22, -17, -61, 50, -56, 78, -18, 19, 61, -56, 1, -44, -17, -75, 125, -73, 87, -87, -102, -27, -7, -107, 40, 113, -57, -102, -31, 127, 30, -22, -102, -12, 30, 107, 24, -21, 61, 86, 94, -84, 103, 90, 39, 109, 14, 65, 90, 79, 97, -109, 39, 56, -1, 17, 96, 51, -44, -21, -90, -6, 79, -43, -64, -2, -11, -8, 58, -22, 111, -66, -128, -66, -40, 28, -42, -12, -39, 58, 119, 114, 111, -114, 16, -46, 86, -128, -87, 124, -4, 78, 46, -81, 75, -74, -78, 66, -8, -94, 66, 68, 81, 48, -106, 58, -58, -49, 92, 112, 24, -121, -55, 84, -10, -120, -116, 84, 59, -42, -85, -111, 60, 13, 50, -4, -115, 8, -108, 78, -32, 107, -79, 27, -77, 126, 33, -16, -61, -83, 60, -29, -53, -54, -20, -80, -83, 33, -70, -40, 9, -96, -30, -95, 115, 117, -36, 88, 63, -125, -50, -72, 46, 62, 69, 42, -15, -34, -77, 124, -84, 123, -91, 103, -67, 61, -117, 8, -128, 84, -114, 24, 126, -72, -9, 23, -84, 107, 47, 60, -32, -63, -19, 25, -94, -56, 80, 66, -91, 9, -57, 81, -110, -58, 4, -94, -105, 0, -74, -116, -102, 26, -116, -65, -80, -16, 8, 127, 86, -80, 60, -128, -110, -126, 15, -73, -67, 109, 8, -126, -103, 37, 95, -39, -85, -56, -73, 105, -24, 76, 91, -45, -38, -102, 61, -87, -36, 39, -10, -82, 96, -87, -109, -50, 108, -107, -94, 67, -126, 102, 114, 36, -26, -60, -87, 46, -52, -60, -79, -79, 81, -7, 70, 90, -109, -105, -6, 100, 49, -75, -22, -117, 75, 66, 49, -106, 30, -103, -52, 87, 7, -82, -101, 99, -122, 36, 36, 70, 40, -93, -56, 6, 35, -4, -27, -120, -118, -44, 82, 95, -107, -112, -109, -114, 99, 94, -95, -30, -55, -17, -37, -97, -97, 101, 3, -31, 6, 45, -33, -94, -90, 110, 102, -84, 116, -113, 88, 19, -110, 125, -68, 58, -53, 118, 68, -58, -13, -123, 9, -82, -90, -117, 101, -73, -36, 34, -128, 104, -4, 108, -82, 110, -43, -114, -94, -93, -109, -29, -104, 50, 125, -128, -15, 19, 39, -123, -69, 94, -98, 90, 84, 11, 37, 74, 108, 113, -55, 51, 42, -117, -3, -6, -126, 51, 47, -31, 120, 11, 53, -28, -106, -108, -9, -107, 34, 114, -51, 124, -11, -16, -14, -42, 123, 42, 84, 41, -4, -85, -50, 33, 47, 2, 31, -13, -27, -92, -118, 96, 73, -120, 99, -31, 37, 109, -41, 30, -99, -126, 0, 68, 102, -95, 52, -9, -127, 98, -6, -15, 74, -26, -11, 31, 70, -81, 60, -20, 8, -27, 121, -112, -71, 114, 68, -117, 69, 108, 69, 7, -108, -45, -73, 116, 18, -30, 69, -98, -117, -57, -119, -33, 82, -20, 35, 37, 81, -99, -111, 97, 22, 45, -24, -55, 121, -32, -100, -79, -54, -126, -47, 113, -6, 1, -102, 111, -82, -19, -127, 99, -61, -52, 28, -1, 35, 9, 11, 90, 86, -124, -12, -84, 109, 42, 52, 1, 13, 64, -116, -57, 102, -79, 66, 44, 62, 117, -45, -128, -98, 102, 57, -125, -59, -85, 105, -121, -91, 92, 1, 95, -74, -57, 121, 53, -78, -56, -104, 8, -121, 68, 68, -52, 96, 101, 36, -108, 52, -125, -82, 96, -32, -91, 14, -24, 76, 45, -13, 29, 110, -60, 91, 68, 72, 57, 18, -84, -66, -124, 40, -5, 89, 8, 15, -45, -68, -61, -23, -62, 38, 100, -81, -58, 51, 9, 83, -89, -70, -2, 16, 88, -33, -120, -89, 118, -102, -127, -121, 102, 43, -53, -27, -54, -84, -40, -10, 70, -39, 60, 34, 16, -113, 10, -76, -88, 47, 115, 46, -53, -41, -84, -32, -58, -32, 90, -112, -66, -112, 84, 54, -124, -58, 82, -73, 38, -25, 5, 42, 66, 126, -93, -115, 107, -25, -37, -10, 6, 111, 73, 88, -38, 121, 21, -110, -78, -76, 44, -62, -46, -64, 31, -58, 49, -53, 115, 75, -85, -14, -125, -73, 31, 84, 103, -106, 20, 24, 47, 39, 10, -52, -49, -63, -46, -31, 14, -35, -112, 70, 8, -60, 6, 127, 102, -5, -102, -68, 39, 114, -54, 104, 115, 40, -55, 38, -76, 13, 26, -82, -68, -43, -85, -72, -45, -28, -14, 49, 20, -90, 51, -78, -62, 127, 122, 55, 90, -70, 30, 95, 32, -85, 18, -128, -113, -81, -110, -86, -30, 125, -127, -33, -65, 121, 22, -64, -82, -10, -66, -18, 80, 1, 107, 26, 57, -59, -112, -112, -15, 107, -109, -88, 73, 111, 126, 68, 44, 26, 123, -39, -113, -42, 1, 29, 43, 123, -79, -118, -93, -116, 77, 20, 35, 97, 63, -108, 79, -116, -57, -49, 49, -8, -55, -74, 70, 96, -85, 4, -112, 35, -79, 68, 95, -60, -102, -3, 69, 13, -62, -38, -13, 106, 2, 78, -119, -74, 6, 39, -54, -127, -10, -118, 4, -103, 22, 87, 68, -87, 45, 88, 110, -62, 111, -57, -48, -63, -27, -117, -4, -49, 20, 11, -126, -88, 68, -121, 82, 109, 3, -103, 36, 48, -44, 18, -15, 77, 31, 104, 57, -28, -83, 27, 11, -117, 98, -103, 30, -34, -56, -60, -113, 4, -97, -14, 109, 125, -121, 110, 21, 102, 118, 43, 22, 72, -64, -87, 33, 106, -11, -33, 32, -99, -88, -15, -95, -111, 34, -55, -89, -4, -76, 18, -77, -60, -25, 110, -70, 9, -81, 5, -35, 8, 2, 73, 75, -6, -67, 43, -109, 56, 45, 45, 62, -83, 125, 87, -111, 70, -115, -75, 107, 28, -112, 32, 95, 124, 35, 10, 107, -43, 97, -58, -45, -51, -23, -101, -35, -120, -26, 114, -35, 44, -23, -44, -83, 12, 107, 26, -28, 49, -90, 34, 7, -17, 117, -102, -90, 32, -31, 18, -100, -113, -88, -60, 58, 64, 38, 12, 119, 41, -56, 79, 21, 41, -72, -2, -119, 27, -10, 21, -11, 75, 105, 12, -68, -33, 46, -31, -49, 118, 47, -69, 5, -116, -116, -25, 68, 99, 82, 95, 95, 57, -125, -35, 93, 37, 104, -62, -59, -46, -105, 54, -120, -40, 124, -92, 126, -110, 2, -2, -90, 0, 124, 33, 33, 22, 66, -60, 44, -36, -7, 90, 125, -92, -71, 91, -20, 93, 34, -36, 41, -120, 19, 20, -112, 88, 100, -125, 122, -58, 4, 19, 52, 45, 89, -110, -118, 114, 55, -118, -36, 76, -85, -69, -73, 76, -19, -91, -36, 29, 0, -109, 82, 100, -37, 89, 82, 14, -115, 59, -52, -15, 64, -123, -33, 126, 102, 58, 12, -24, -17, 38, 99, -126, 68, 56, 95, -66, -61, -102, 107, 70, -108, 126, -75, -11, 94, 78, 3, -67, 81, 44, 109, 122, 35, 19, -91, 14, 63, 19, -115, 94, -91, 72, 53, 120, -2, -34, 1, 54, 119, -87, 116, 77, 93, -21, -24, -108, 99, -33, 85, -74, -121, 79, 75, -98, -23, 78, 101, 108, 41, -42, -46, 70, -59, -108, 16, 122, 80, -1, -104, -88, -5, -6, -17, 124, -126, -2, 95, 6, 68, 103, -57, -90, -41, -81, -51, -9, 39, -52, 19, 73, -97, 126, 9, -71, -25, 32, 34, -76, 72, 7, -89, -18, 61, -109, 63, -32, 92, 48, -122, 79, -54, 18, -38, 48, -3, 120, 40, -118, 44, 99, 67, 0, 30, -4, 126, 94, 82, 32, 38, 22, -115, 75, 83, 116, -111, 61, 54, 90, 78, 54, 29, 98, 25, 96, -124, 120, -36, -4, -96, -64, 88, -2, 40, 19, 115, -125, -21, 64, -125, 74, -91, 64, -107, 52, -30, 42, -123, -101, -4, -69, 32, -95, 108, 45, -97, -4, -115, -62, 56, -11, 4, -63, 60, 63, -123, 121, 115, 89, -30, 126, -99, -93, -45, -38, -98, -118, -35, 0, 66, 32, 60, -99, -2, 94, -127, -21, 91, -114, -15, -10, 13, -2, 22, -102, 113, 73, 127, 123, -54, -102, 81, -102, -88, 43, -78, -9, 38, 50, 86, 17, 56, -92, 33, -75, 127, -87, 48, 91, 108, -53, 114, 126, 65, -120, -41, -52, -85, 97, 85, -65, -43, -18, 12, 42, 113, 92, -58, -126, 30, 80, 58, -38, 76, 38, 42, 90, -45, -71, 35, 70, -83, -85, 42, 101, -12, -77, -107, 0, -93, -105, -120, 98, 1, -49, -127, -110, -85, 58, -3, -115, 44, -76, 52, 39, 78, -9, 101, 5, -92, -60, -30, -75, 9, -6, 28, -106, -14, -106, 59, 52, -27, 2, 68, -25, -100, 17, -50, -40, 112, -29, -88, -125, 102, -119, -4, 30, 116, -58, 110, 84, -85, 90, -102, 86, -21, 124, 38, -13, -103, 119, -60, 14, 27, 53, -43, -86, 80, 56, -128, 78, -100, 39, 77, 39, 127, -116, 81, -7, 50, 8, -52, 30, 126, 92, 72, -87, -95, 126, 122, 18, 119, -127, -45, -37, -2, 38, -35, -122, 25, 76, -25, 70, -115, -30, -8, 58, 66, -70, -26, 86, -75, -10, -40, -106, -82, -24, -126, -66, 42, 66, -14, -17, 47, 42, -117, 114, 97, -83, -35, -84, -57, -19, -116, 7, 101, 118, 125, -53, 108, -102, 81, 83, -58, -71, 68, 59, -58, -58, -120, 119, -107, -111, -11, 79, 76, 57, -36, 7, -118, -19, 28, -65, -15, 81, -68, -48, 66, -15, 87, -102, 85, -30, -126, 86, 125, 20, 4, -41, 14, 58, 10, -5, -103, 100, 54, -13, -53, -95, 18, 124, 12, -47, 47, 22, -67, -74, -112, 77, -99, 98, -108, -123, -30, 110, -97, 40, 84, 113, 34, -59, 48, -99, -87, 88, -110, 57, -10, -43, -122, 4, 123, -2, 87, 67, -115, -52, 51, -77, -113, -24, -114, -53, 111, 29, -107, 87, -57, 90, -112, -94, 76, 77, 69, 94, 82, -60, 87, -37, 84, 59, -24, 8, -84, -106, 43, 118, -61, -32, 7, -114, -127, 118, 117, -53, 12, -62, -48, 6, -6, 58, -81, -17, -16, 78, -59, 97, 29, -73, -124, -96, -116, -52, 121, 80, 74, -116, -15, 30, -27, -101, -7, -59, -25, -62, 90, -21, 67, 37, -85, 116, 32, 10, -125, -74, 10, -75, -18, -34, 74, -112, -15, 4, -121, 124, 111, 105, 111, -75, 72, -56, 59, -64, -24, -34, 68, 50, -58, 51, 28, 54, -122, -10, 33, -62, 2, 114, -54, -101, 68, 0, 44, 29, 21, 70, 58, 111, -91, 21, -107, 52, -108, -110, 37, 62, -70, -78, 126, 26, -120, -24, -67, 85, 38, -28, 78, -24, 13, 38, 40, 71, 49, -28, 14, -47, 111, 66, 70, -84, 39, 94, -108, 52, 24, 44, -7, 71, -55, 5, 121, 127, -13, 26, 10, -120, -85, 71, -13, -11, 119, -79, 52, 120, -9, 30, -94, -29, -8, 115, -128, 85, -9, -93, 9, 2, -12, 68, -58, 25, -66, 40, 58, 51, 39, 94, -43, -125, 116, -57, -128, -22, -3, -31, 21, 119, -97, -112, 85, -85, -30, -91, 60, 76, 24, -65, 118, 77, -84, -75, 58, -52, 10, -91, -122, 74, -106, -41, 119, 73, 114, 51, -42, 87, 85, -97, 24, 111, 47, 101, 102, -112, 54, -117, 4, 30, -63, 77, 21, 17, 27, -24, -127, -113, 56, -47, -128, -31, 23, -87, 50, -11, 112, -89, -5, 80, -104, -54, 17, 36, 43, -94, 110, -10, -36, -70, 120, 107, -4, -36, -6, 43, -29, -95, 113, 84, -30, -86, 118, 46, 20, -57, -48, 41, -15, 13, -62, 81, -105, 63, -12, -47, 70, -57, 30, 65, -128, 113, 34, 66, -127, 91, 124, -71, -111, -100, 90, 1, 44, -34, 38, -98, 110, -3, -122, -115, 98, -14, -61, 1, 113, 11, 11, 1, -10, -126, -95, -61, 39, -19, -42, -20, 33, 61, 127, -80, -24, -83, 56, 1, -58, 93, 88, -118, 33, 122, -58, -10, -94, -28, -4, -114, 68, 0, 51, -45, -52, -27, -117, 38, -47, -116, 37, 67, -79, 51, -59, 21, 41, -10, 126, -108, 122, 16, -107, 5, -119, 92, -19, 70, -107, -14, -55, -106, 45, -9, 35, -11, 108, 99, -91, -2, -72, 122, 5, -55, 98, -110, -32, 13, -83, 37, 113, 100, 54, 48, -123, 4, -124, 96, 41, 3, 121, -63, 86, 102, -100, -5, 65, 42, 104, 72, 58, -42, -126, 95, 41, -93, -55, 93, -66, 4, -49, 79, 117, 60, -110, 66, -66, 93, -30, 10, -23, -94, -69, -114, -62, 89, -77, 126, 110, 82, 12, 72, 84, 42, 59, 75, 58, -100, -123, -46, -70, 33, -2, 10, -16, 31, 12, 102, 43, -100, 114, 99, -74, -42, 68, 105, -68, 106, -104, -118, 25, 126, 11, -63, -30, 85, 64, -111, 45, -32, -85, 81, 8, -124, 38, 43, 98, -52, -37, -60, 122, 105, -110, 35, -127, 116, 55, 11, 7, -61, -100, -34, -11, 78, -111, 61, 123, 25, 84, 13, 109, -37, -111, 120, 57, -31, 77, -58, -58, 23, -46, -128, -18, 13, 63, 39, -83, -22, -61, -22, -124, -39, 107, -64, 126, 50, -28, -23, 22, -13, 109, 30, -8, -6, -14, -17, 1, 52, -122, -68, -126, -28, -24, 11, 12, 85, -105, -123, -44, 122, -31, -50, 85, 45, 93, -35, -114, 41, -49, 116, 118, 80, 49, -55, -44, 25, 27, 42, 6, -26, 75, -45, -96, -52, 110, -58, -37, -108, 8, -66, 122, -53, 82, -100, 69, 64, -35, 80, -53, 35, 54, -64, -96, 49, -56, 47, 8, -122, -42, 40, -95, 89, -126, 78, 116, -3, 11, -75, -37, 28, 117, -91, 54, 50, 36, -84, -3, -87, 119, -45, 116, 8, 6, -103, 8, 96, 101, 61, 56, 115, -114, -97, -69, -124, 23, -55, -25, 104, 102, -1, 37, -126, 74, 39, -8, 107, -74, -64, 75, 68, -83, -77, 63, -24, -40, 32, -86, 114, 82, 75, -114, -90, -112, -74, -112, 43, -75, -59, -31, 77, 10, 48, 31, -108, 71, 99, -125, -123, -12, 13, 5, -65, -42, -11, -29, -39, 127, -77, -27, -111, 3, -114, -51, 119, 72, 78, -102, -41, -26, -38, 91, 1, 5, 55, 108, 62, 87, -112, 76, -21, 115, -12, -62, 114, -36, -58, -26, -15, 56, 53, 119, -32, 108, 67, 42, -24, 126, 34, -35, -26, -104, 52, -102, 1, 1, 79, 26, -128, -81, -128, 57, 57, -31, -34, 120, 84, 50, 48, 55, -14, 88, 80, -82, -108, 121, -10, 108, -44, -12, -89, -7, 5, -23, -50, 68, 22, 80, -56, -114, 2, 12, -47, 13, -95, 38, -63, 90, -126, -1, -61, -62, -50, -38, -50, 104, -92, -46, -17, 127, -128, -51, 89, -51, 107, -68, 3, -50, 49, -91, -127, 37, -45, -29, 77, 19, 78, -73, 22, -118, 7, -3, -100, -106, -104, -53, 117, -122, -56, -117, 63, -77, -41, -63, -55, 58, -109, -29, 39, -73, -45, -92, 41, 10, -22, -122, 0, 22, 28, 36, -79, -40, 114, 37, 72, 67, -85, 34, 79, 47, 113, 19, 102, -127, -37, -55, -31, 14, -3, -76, 101, -57, 31, -8, 81, 60, -70, -113, 27, 16, -6, 108, -2, 113, -89, 125, 85, -89, -76, -76, -26, 72, -109, 79, -21, 46, -52, -121, 68, -67, -70, -94, 77, 118, 40, 117, -88, -77, 96, 88, 55, -112, 37, -1, -34, -106, 44, -100, -29, -114, -33, 113, -98, -115, -33, -57, 122, 9, 28, 55, 120, 89, 74, -22, -37, -88, 43, -69, -102, 35, 101, 7, -84, -71, -24, 35, -116, -69, -35, -44, 85, -110, -101, -70, 85, 10, 115, -86, -87, 2, 109, 36, -29, 37, 120, -98, -19, -87, 42, 64, -12, -79, -82, -89, -95, -72, 40, -106, -48, 60, 61, 90, 120, 65, -112, -92, -84, -16, -121, 48, -4, -5, -52, 106, -32, -76, 61, -41, 66, 99, -38, -108, 58, 79, 80, -45, 99, 35, -84, 89, 9, -119, -93, -43, -58, -3, -48, -23, -47, 69, -53, -101, -15, 80, -12, 125, 93, -113, -96, 110, 87, -86, 117, 92, 44, -45, 29, 115, 14, -64, 105, -94, -79, -51, 25, 68, 10, -128, 48, -7, -56, 93, 100, -38, -85, -53, 110, -8, -52, 117, 76, 89, -39, -78, 46, 86, 102, -34, 43, 51, 18, -126, 75, 2, 36, -27, -44, -67, -32, 96, -105, 111, -15, -112, -96, -102, 9, -6, -26, -43, -80, 103, -121, -113, 127, -118, -26, -53, 43, -27, 90, 24, 89, 90, 7, -128, 121, 29, -4, 118, -76, -21, 68, 122, -76, -64, -26, -78, -21, -118, 3, 46, 104, -104, -105, -77, -124, 100, 75, 83, -61, -125, 70, -33, 109, 64, 43, 22, 27, -124, 1, -90, -109, 19, -72, 48, -125, -126, 57, -63, 97, -28, 100, -92, -17, 79, -54, 92, 64, -16, 32, -72, 104, 36, -22, -67, 83, -58, -98, -112, 46, 69, 105, -101, 118, 10, -59, 77, 73, 26, 122, -81, -62, -40, -86, 103, 68, 25, -64, -24, 9, -3, 80, 44, -102, 67, 118, -25, 53, -96, 51, -71, 124, 32, 75, -91, -72, 84, 73, -96, -23, -125, 116, 69, 59, 107, 15, -64, -108, 85, -103, 6, -122, 53, -110, -24, -39, -104, -9, -56, 84, -127, -77, -17, 19, 27, -7, 103, -44, -37, 3, -72, -3, -80, 21, -111, 103, 112, -85, -125, -33, 106, 68, -28, -30, -29, -31, -3, 17, -11, 101, -85, 90, -104, 59, -111, 21, 97, -93, 105, 62, -90, -72, -108, 43, 123, -3, 12, -2, -107, -36, 126, -77, 67, -36, 16, -68, -41, 124, -67, 74, -46, -49, -117, -125, 65, -40, -22, 104, -99, -18, 57, -10, -17, 25, 65, -10, -14, 28, 23, -109, 117, 44, 104, 54, 116, 125, -13, -54, -121, 96, 99, -28, -102, 27, -126, 38, -44, 35, 54, -26, -115, 3, -81, -52, 112, -43, -39, 72, -84, 3, 20, 37, 92, -78, 7, 73, -93, -74, -9, 111, -65, 68, 4, 78, 67, -58, -104, -114, 15, -58, -94, -84, -74, 75, 45, 116, -103, 115, 85, 60, -102, -72, 78, 96, 55, -12, -10, -103, 72, -97, 101, -60, 111, 44, 14, -24, 104, -43, 61, -96, -55, 11, 85, -72, -82, 127, -81, 60, -30, -55, 52, -55, 36, -40, 0, 103, -92, 25, 89, -125, 23, -127, 45, 31, 73, -85, -125, -99, 83, -1, -64, -49, 24, -94, -52, -79, 102, 66, -126, -6, 94, -20, -48, -70, -95, -32, 28, -120, -18, -7, -91, -95, 71, -88, 119, -28, 60, 4, 18, -49, -105, -104, -94, 33, 56, 87, 30, 27, 72, -2, 84, -102, 58, 96, 34, -6, -21, 103, 81, -95, -123, 76, 90, 59, -106, 122, -116, -102, -44, -5, -79, 52, -107, 113, 114, 43, 71, 56, -128, 82, 127, -41, -92, 79, 77, -34, 124, 16, -99, -47, 80, 26, 97, 83, -87, 107, 39, 85, -120, -42, 103, -108, 4, 122, -102, -63, 85, -68, 46, 123, 27, 79, -17, 34, -122, -68, -2, -62, -115, 96, 99, -56, 83, 93, -119, -64, 30, -92, -53, 34, -41, 87, 45, -49, -26, -121, 121, 79, -14, -43, 71, 61, 56, -11, -93, 43, 121, 6, -72, -107, 114, -48, -33, -81, -8, -81, 8, -72, 18, 69, 14, 34, 8, -78, -101, 53, 77, -100, 113, -21, -68, -54, -14, 102, -65, 46, -92, -44, 61, -110, -123, 103, 38, -98, 107, 11, 65, 0, 10, -97, -125, -71, -110, -90, -14, -1, 6, 88, -17, -57, 40, 26, -26, -2, 34, 108, 6, -113, 44, -49, 54, 18, 61, -92, 125, -125, 117, -73, 61, 69, -21, 66, -41, 22, -87, -128, -104, 39, 72, -114, -42, 95, -93, 107, -100, 0, 77, 62, -102, -13, -67, 94, -19, -12, -123, -44, 24, 69, 37, 97, 72, 0, -95, 58, 116, 53, 66, -75, 55, -100, -7, 20, 123, -9, 113, -32, -13, 75, -63, 48, 55, 30, 39, 14, 17, -113, -57, -15, -10, 46, 123, -50, 71, -39, -84, -79, 74, -72, 52, 5, 75, -86, 96, -55, -49, 3, -3, 123, 28, -92, 84, -6, 3, -92, 13, 8, 120, 30, 94, 84, 123, -97, 13, -107, -5, -71, -57, 105, -125, 108, 98, 127, -79, 40, 111, -66, 22, -34, -89, -116, 15, -57, -26, 114, -80, -84, 99, -46, 101, 72, 53, 57, 96, -109, -64, 35, -30, -18, -86, 45, 126, -23, 115, -21, 14, -3, 71, 100, 80, 113, -9, 32, -53, 41, -123, 92, -113, 28, 116, 15, -94, 62, -113, -119, -93, 67, -50, 4, 59, -112, 41, 63, -116, 1, 63, 45, -41, -12, 18, 115, -72, 54, 33, -48, -74, 6, -74, -21, -97, 71, 103, -121, -67, -19, -15, 99, -91, 103, -74, 14, 110, -104, -58, 36, 10, -79, 37, -21, 5, 63, -3, 62, 6, -103, -14, 73, -128, 105, 17, 127, -45, 114, -36, -15, 102, -83, -94, 65, -97, 95, -55, -26, -68, 6, -34, -49, -126, -96, -40, 126, -107, 116, 76, 108, -111, 57, -115, -113, 70, 24, 124, 11, -71, -89, -3, -82, 56, -102, 122, -108, -75, -92, -58, 37, 31, 69, 101, 86, 71, 82, -38, 48, 71, -60, -72, 119, -18, -88, 106, -96, 89, -78, -90, -39, 14, 54, -94, 35, -128, -118, 15, 88, 19, 64, -64, -20, -61, 105, -65, -3, -96, 61, 87, -77, 22, 2, -96, -84, -52, -60, -33, 54, -98, 82, 18, -81, -54, 64, -114, -57, -42, 125, 79, 114, -92, -85, -28, -2, 5, -81, -126, -122, 5, -17, 83, 1, 43, -15, 64, 42, -99, 83, 37, -118, -41, -127, 85, -55, -43, 113, 6, 82, -29, 123, -18, -92, -119, -73, 121, 11, -111, -80, -72, -120, -28, -89, -94, 56, 1, 56, -101, 24, -107, 25, -128, -61, 18, -4, 55, 103, -43, -83, -105, 121, 76, 96, -5, -81, 46, -100, 67, 16, 59, -19, 60, -53, 112, -105, 110, 75, -119, 77, 36, -45, 64, -66, -100, -12, -73, -87, -121, 47, -92, 102, -16, -122, -21, 79, -43, 18, -18, -111, 106, -8, 34, 53, -112, -8, -85, -85, -5, -33, 83, 78, -56, 55, -8, -120, 60, -18, 91, 127, -126, 94, -90, -45, -17, -36, -68, -79, -77, -2, 5, 89, -55, -46, -61, -75, -20, 33, -23, -111, 2, 76, -125, 27, 44, -5, 3, 29, -86, 68, 1, 1, 38, -93, -125, -14, 47, 58, 24, 7, 121, -2, 115, -98, -17, -125, 107, 41, 31, -119, -74, -20, -65, 36, 73, 1, 93, -76, -76, 65, 7, 125, -65, 68, -7, -2, -62, 35, -48, 97, 15, 98, 109, -27, -127, 74, -37, -97, 22, 39, -108, -33, -124, 55, 64, 120, 89, 21, -95, -56, 33, -111, -9, -37, -92, -21, 90, 117, -124, 15, 110, 109, 24, 18, 115, -32, -127, 21, -87, -91, 100, 66, 105, -114, -63, 111, -20, -97, -99, 77, 80, -25, -46, 18, -119, -110, 59, -55, 55, -17, -104, 66, -84, 68, -68, 102, -82, -94, 32, 125, -37, 109, 77, 59, -128, -34, -45, 122, -38, -105, -101, -77, -2, -106, 17, -5, 19, -98, -40, -13, 18, 53, 105, -28, -31, -106, 50, 125, -67, -120, -111, 120, 81, 57, -85, 72, 53, 97, 65, 105, 85, -21, -42, 10, 61, -8, 46, -62, 78, 93, -125, -100, -41, 83, 2, 60, 6, 82, -75, 76, 51, -9, -95, -58, 8, 2, 52, -69, -59, -50, 67, 5, -25, 23, 23, 51, 70, -110, -47, 12, -83, 41, -3, 24, -78, 101, 13, 93, -89, -102, 36, -66, -2, 47, 7, -19, 78, 20, -47, -97, 72, 34, 102, 17, -78, 54, -80, 30, -120, 2, -5, 70, 44, 43, 0, 87, 13, -21, -11, 114, 127, -82, -121, -94, -106, -26, -110, 125, -123, -126, -67, 18, 53, 112, -63, -82, 106, 57, 57, -5, -75, 106, -40, 51, -9, -52, -15, 90, 30, -52, 55, 105, 114, -80, 119, 120, -78, -1, -74, 105, -81, 67, 101, 54, 106, -123, -77, 41, 18, 56, -81, 107, -121, -38, 61, -76, -48, 66, 110, 85, 72, 101, -71, -124, 110, 10, 84, 45, 122, 57, -9, 19, -32, 107, -61, 1, 95, 102, -95, 24, -115, -69, 53, 4, 80, 96, -31, -9, -69, 93, 42, -14, -125, -69, -95, 44, 40, -10, -25, -26, 86, 99, -86, 67, -114, -66, 23, 60, -58, -111, 112, 5, -54, 110, 87, 9, 20, 95, 23, -79, 47, 90, -88, -99, -84, -51, -7, -37, 8, -48, 99, 49, 57, 81, -7, -13, -45, -9, 74, -47, -83, -123, -23, -5, 108, 88, -49, 89, 109, 54, -119, -40, 38, -44, -82, -12, -50, 89, -39, -106, 102, -37, -6, 120, -88, -28, -30, -112, -115, 16, -96, 27, 39, -75, -128, 98, -77, -93, -41, 113, 38, -92, 79, -14, 95, 82, 25, 109, 72, -119, -125, -52, -21, -66, 59, -63, -95, -4, 87, 75, -20, 122, 105, 65, 116, 30, -30, 78, 94, 14, -25, -93, 113, -60, 17, -96, -104, 1, 92, 66, 27, 8, 113, 113, 17, -25, -95, 101, 99, -41, 38, 65, -15, 108, 54, -95, 114, 99, -16, 56, -113, 94, -108, 54, 28, 70, 92, 86, 82, -16, -92, -89, -1, 48, -47, 14, -49, 64, 80, 79, -11, 26, -95, -61, -31, 41, -99, -64, -99, -114, 78, 51, 9, -52, 42, 2, -54, 107, 32, -108, -48, -60, 35, 38, 6, -43, 75, -38, -54, 35, 12, -72, -6, 110, -83, 118, 45, -50, -2, 122, 127, 127, -53, 1, 121, -63, 123, -34, 21, -62, -11, -81, -96, -5, -70, 125, -50, -4, 114, 37, 126, -50, 95, -60, 75, -61, -10, 50, -123, -24, -100, 61, -20, 63, 68, 73, -71, -118, 30, -34, -38, -83, -48, -55, -125, -96, 86, -57, -44, -118, -115, -32, -95, -55, -82, -115, 4, 95, -54, 54, -16, -69, -102, 59, 79, 116, -72, 6, -78, -52, -35, -54, 6, -50, -12, -25, -42, -78, 119, -15, -70, -35, 74, 58, -41, -115, 49, 74, -29, 72, 119, -25, -58, 45, -52, 109, 86, 41, -49, -97, -115, 75, -76, -56, -20, 113, 22, -60, 121, -19, -29, 105, -14, -28, 48, -38, 36, 19, -14, 110, 45, 47, 33, 57, 86, -74, -21, -34, -10, -23, -112, 74, -115, 13, -102, -14, -127, 8, -65, 42, 81, 109, -35, 106, -9, 105, 74, -115, 52, 62, 17, -46, -45, -71, 20, 76, 52, -110, -123, 61, -21, -13, -76, 14, 1, -128, 109, 58, -64, -111, -71, 70, -115, 43, -38, -79, 49, 125, -49, -55, 121, -90, 59, 48, -9, -127, -37, 61, 49, 31, 79, 115, -86, -62, -71, -112, 32, 65, -68, -107, 39, 60, -86, -113, -51, -34, 115, 19, 83, 90, -87, -24, -81, -119, 115, 21, -91, -123, -102, -38, -115, -69, 2, 86, 6, 109, 25, 93, 38, 120, 50, 39, -119, 30, -45, -8, -125, -74, 8, -119, 11, 15, -41, -55, 49, -42, 15, -119, 111, -4, -84, -70, -123, 59, -2, -51, -102, -12, 39, -116, 29, -6, 121, -38, -59, -52, -50, 80, -13, -52, 52, -34, -81, -127, 38, 78, -97, 13, -55, -58, -85, -80, -24, 19, 50, 75, 73, 22, -49, -78, 84, -103, -48, -56, -88, 90, -95, 6, 67, -47, -7, 17, 118, -98, 119, 30, 109, 88, -101, -25, -110, 45, 39, -76, 43, 26, 46, 55, 48, -106, 95, 29, 11, -108, -15, 104, 101, -1, 122, -101, -115, -37, -128, 47, -41, -78, 112, 122, -83, -58, -76, -85, 98, 88, 31, 92, -118, 61, 12, 119, 9, 34, -15, -76, -119, 123, 36, -72, 122, 97, -58, 97, -40, 90, 12, 23, -2, 47, 88, -81, -8, -11, 44, 23, 89, 77, -52, 120, -75, 125, -100, -67, -108, -65, 79, 104, -95, -30, -113, 20, -19, -35, -25, -72, 65, -8, 111, -113, 32, 32, -84, -112, -56, -96, -11, -42, 59, -36, 127, -18, 6, 30, -128, 123, -85, -50, 33, -86, -35, -25, -77, 28, 90, 84, -69, -64, 35, 65, -90, -7, 71, 8, -105, -120, -86, 0, -69, -78, 46, -11, 79, 70, 49, 20, -1, -47, -73, 124, -121, -123, 95, 123, 101, -62, -11, 118, 29, -16, -76, -53, -17, -46, 29, 82, 56, 87, 96, -47, -21, -34, -67, 95, -12, 49, 23, 10, 113, 98, 6, 13, 22, -93, -74, 30, 118, -94, -2, 38, -60, -28, -3, 83, -25, 70, -121, 41, 100, 118, -95, 6, 35, 72, -98, -30, 13, 5, -40, -59, -23, 5, 27, 123, 60, -67, -94, 13, -71, 96, 30, -127, 46, 77, 124, -122, 3, 26, 120, -6, 37, 119, 59, -110, -11, -50, 120, -120, -5, -101, 36, 32, -1, 7, -81, 11, -122, -91, 47, 84, -40, 127, -87, 107, -4, -35, 108, -61, 10, 124, 18, -11, 29, 56, -124, -127, -42, -57, -110, -16, 20, 5, -28, -123, 67, -12, 97, -30, 124, 125, -60, -18, -117, 52, 73, 102, 64, 97, -85, 126, -31, 13, 32, 114, -44, 67, 4, 72, 67, 92, -52, 62, 23, -63, -84, 115, 68, 44, -113, -5, -64, -87, 56, -90, -15, -86, 5, -9, -2, -110, -19, 22, -4, 89, 43, 104, -73, -48, 126, -94, 77, 37, -59, -77, -66, 113, 97, 56, -127, 67, 36, -106, 15, 37, 77, 115, 124, 98, 70, 7, 0, -34, 93, -25, -64, -41, 18, 105, -127, 75, 56, 44, 9, 49, 83, -8, -22, 127, 69, -48, -108, -123, -101, 25, -17, 27, 74, 71, -39, -92, 108, 92, 12, -15, 41, 55, 38, -51, 122, 23, -21, -112, -68, 101, -36, -7, -127, -62, 127, 89, -37, 95, -105, -46, 26, 23, -108, -72, -95, -46, -96, -41, -28, -76, 22, 62, -70, -72, 90, -70, -52, 93, -55, 123, -53, -57, -28, 109, -117, 89, -62, 120, 59, 29, -6, -18, -116, 101, 8, 35, -89, -41, 33, -68, 19, 16, 114, -88, -57, -101, 18, 64, 117, -74, -10, -60, 107, 96, -72, -14, -7, 46, -38, -67, -109, -51, 118, -103, 14, 69, -59, 36, -87, 110, -109, 14, 62, 33, -97, 16, 21, -80, -79, -56, -128, 77, 99, -4, 105, -20, 95, -12, 88, 95, -117, -51, 23, 117, 85, -70, -78, 113, 104, -9, 10, -25, 108, -27, 23, -13, -63, 56, 24, -28, 11, -127, -54, -59, -100, -41, -46, 118, 1, 73, -9, 15, 61, 2, 37, 76, -120, 127, 121, 48, -34, 104, -79, -71, 118, -97, -8, 70, -100, -96, 0, -7, -17, 89, -123, 34, -118, -70, -103, 2, 39, -77, 90, 38, -24, 79, -13, 117, 91, -91, -53, -17, -5, -47, -7, -112, 60, -105, -87, 66, -7, 3, 63, 11, 38, -7, 86, 12, 71, -83, -55, -4, -104, -116, 38, -47, -127, -59, 0, 92, 24, 68, -91, -111, 84, 37, -92, -123, -92, 71, -116, -94, -70, 101, 95, -113, -81, -116, -48, 76, 41, 20, -100, 18, -125, 87, 120, 15, 50, -13, -73, 68, -125, -109, -100, -91, -82, -13, 86, -119, 77, -31, -97, 71, -96, 84, 126, -37, -22, 69, -59, 80, 122, -48, 51, -76, 59, 82, 37, -52, -84, 8, -10, -45, -128, -23, 75, -93, -47, 34, 3, 31, -34, 0, 32, -128, -25, 32, 61, -19, 42, 50, -41, 94, -93, 126, -22, 54, -55, 59, 79, -113, 89, -53, -85, 105, -25, 7, -76, -110, 101, 105, -125, 67, -128, -60, -111, 100, 53, -68, 111, -54, 113, 2, -28, -34, -96, 62, -46, 87, 78, 117, 76, -57, 7, 4, 80, -53, 123, 97, -114, 14, 97, -80, 56, 37, 48, -99, -22, 18, 109, 61, 104, -13, -44, 33, -32, -67, 105, 103, 43, -80, -49, -97, 72, 24, -79, -121, -63, -105, -13, 36, 107, -71, -99, -74, 101, 48, -60, 28, 4, -51, 3, -65, -97, 72, 11, -34, 30, -108, -68, 85, 17, -86, -65, 81, -42, -66, 52, 42, 99, -6, 39, -96, 49, -79, -2, -17, 29, -116, 72, -93, -14, 41, -76, 63, 87, 55, 16, -106, -57, -2, 12, 40, 47, -117, 58, 99, -118, -111, 92, -82, -49, 116, 115, -85, 110, -82, 40, 4, 57, 74, -93, -40, -56, -114, -96, 60, -14, 126, -13, -31, 51, -12, -107, 96, 55, 108, 96, -35, 77, 127, -63, -71, 96, 23, -107, -12, -52, -19, -67, -5, 105, 121, 60, -126, -95, -16, 70, 45, 54, -107, 7, -10, -124, 12, -121, -110, -95, 38, 31, -8, 48, 31, -75, -26, -123, -40, -33, 12, -127, -75, 80, 121, -20, -42, -70, -120, -72, -87, -36, 62, 87, 100, 82, 10, -96, -22, 102, 0, 63, 6, 81, -5, 89, -106, -47, -31, 82, -32, -72, -103, 76, 102, 59, 28, -47, 63, 118, 92, -30, -61, -74, 77, -43, -112, 41, -37, -50, -43, 111, 20, -98, 103, 15, -101, -54, 124, -126, -95, 67, -77, 14, 110, 22, -104, -65, -81, 117, -65, -34, -119, 49, 9, 62, 9, 19, 90, 24, -106, -13, -49, -93, -9, 84, -70, -116, 110, 53, 0, -40, 3, 42, -33, -52, 119, -71, 70, -78, -50, 25, -34, 110, 107, -103, 20, 32, -56, 90, -77, 11, 74, -18, -76, -17, -122, -114, 9, -96, 4, -118, 121, 37, -51, 71, 52, 75, 31, 30, -101, -90, 112, -37, 102, 59, -20, 41, 97, -50, -82, 13, -11, -95, 19, 67, 47, 118, 86, 103, 56, -8, -12, 71, 47, -23, -43, 100, -75, 107, 101, -98, 80, -38, 12, -124, 77, 26, 105, -40, -101, -124, 46, 96, -121, 90, -36, 113, 117, 125, 109, 107, 100, 66, 17, 31, 47, 83, -32, -51, 89, 70, -62, 33, -32, -7, 12, 31, 19, 6, 115, 100, -91, 37, -20, -38, -101, -51, -113, 69, -80, -35, 122, -66, 116, 90, -73, -61, -59, -62, 86, -67, -65, 37, 72, 109, -41, 65, -20, 12, -87, -41, -82, -36, -99, -43, -121, 19, 64, -101, 0, 59, 42, 77, -111, -60, 17, -52, 85, 78, -120, -52, -52, -35, -97, 112, -88, -106, 87, -7, -20, 52, 71, 27, 105, 89, 27, -26, -39, 30, -89, -55, 109, -30, -38, 119, 44, -16, 34, -26, -94, -13, -112, 116, 13, 29, 107, -98, -88, -1, -70, 92, 104, -89, -86, 56, -22, 122, 62, -5, 119, 67, -49, 115, 4, -109, 45, -27, -97, 5, -73, -117, 126, 120, 43, -59, -108, -11, -86, 38, -36, 25, -67, 11, 126, 65, -64, 48, -114, 1, 95, -81, 46, -45, -1, -124, 67, 55, -112, -46, -28, -62, 51, -94, 32, -6, -73, 95, 119, -120, -42, -90, 61, -117, -91, 61, 106, -128, 90, -72, -25, -41, 51, 59, 74, 111, 30, 127, 51, 35, 62, -10, -68, -117, -114, -121, -95, 47, 46, -71, -46, 93, -101, -93, 36, -55, -102, -99, -102, -120, 2, 75, -107, 45, -98, 10, 83, -104, -32, 39, 65, -17, 42, -114, 100, -112, 8, 89, 39, -57, 67, 79, -94, -69, -1, -77, -30, 16, 112, 55, -74, 126, 76, 85, -58, -4, 22, -72, 58, -42, -95, 8, -6, -105, -89, 32, 104, -109, 110, 8, -45, 96, 64, -100, -36, -86, -115, -37, 119, 2, -19, -106, 98, -89, -55, 62, 82, -44, 18, 69, 103, -100, 100, 39, -63, -97, -56, -118, -65, -29, 33, -113, -35, -104, -37, -99, -59, -83, 32, 88, 51, -89, -20, 75, 124, -119, 5, 124, 72, -76, -74, -91, 106, -58, -43, -97, -127, 75, -19, -47, -81, 77, -9, -125, -21, 80, -102, -120, 96, -81, -83, 72, 64, 19, 67, -51, -57, 106, -97, 112, 91, 62, 28, -5, 98, -63, -54, -115, 104, 111, 21, -54, -102, 26, 60, 95, 56, -43, 97, -4, 121, 76, 111, 111, 48, 29, -16, 108, 27, -48, -23, -111, -44, 11, -96, 45, -53, 36, -73, 1, 90, 5, 73, 44, -42, -126, 2, -31, -81, 12, -62, 64, 98, 85, -51, -26, 62, -13, -58, -37, -70, -7, -89, 10, -109, 91, 70, 116, 68, 17, 90, 99, -56, -17, 54, -42, -100, 85, 35, -10, 120, -117, 6, 32, 122, 126, -98, 22, 89, -81, 23, 58, 104, -126, 38, -59, 111, -52, 116, -116, 99, 35, -77, -10, -61, 102, -71, -39, 89, 85, 120, -70, 123, -99, -26, 68, 53, -68, 63, 9, 85, -45, 16, -17, -127, 122, -13, -4, -27, -54, 9, 67, -110, -9, 88, 62, -88, -16, 80, -20, 119, 110, -9, 49, 20, -31, -31, -12, 127, 30, 14, 18, -126, -50, -97, -92, 22, 52, -97, -101, 84, -49, 84, -37, -90, 45, -8, -42, -105, -80, -118, 5, 97, 39, 121, -34, 80, 24, 63, 23, 64, -50, 67, -117, -70, 76, 72, 17, -127, -114, 63, 116, -39, -43, -95, -113, -101, -85, 90, -10, 103, -44, -8, -9, 124, 71, 73, -60, 77, -83, 0, 104, 116, 81, -46, 8, 86, 44, -105, 15, 53, -63, -12, 14, 64, 111, -29, -43, -76, -78, -54, 97, 30, 90, -32, -6, 120, 119, -92, 22, 62, -95, 46, -55, 81, -16, -27, 53, 60, 86, -53, 107, -123, 33, -122, -123, -77, -98, 76, 5, -63, -109, -119, -106, -121, 120, -86, -9, 122, 51, -14, -32, -67, -39, -94, -6, -124, 87, 81, 42, -94, -36, 78, 109, 6, -121, -89, 109, -29, 8, 77, 104, 104, -13, -83, 89, -7, 4, 52, 17, -128, 76, -71, 48, -43, -100, 93, -43, -22, 76, -109, 100, -13, 64, -8, 92, -21, -109, -71, -124, -105, 19, 74, -117, -93, -97, -125, 96, -95, -122, -8, 118, 73, -47, 64, 59, -36, 40, 83, 50, -51, -16, -31, 49, 70, 33, -112, 85, 29, 26, -2, 7, -67, -122, 34, 88, -12, -65, -100, -1, -118, -112, -3, -37, -51, 35, 66, -11, -34, 19, 93, 47, -94, 61, 64, -92, 84, -75, 25, 90, -126, 60, -86, 60, 71, -42, -92, 73, 114, 66, -69, -17, -46, -67, -69, -45, 104, 72, -34, 33, -54, 104, -2, 62, 105, -76, 60, 114, 108, 45, -102, 22, 20, 34, -22, 79, 27, -82, 54, -52, 77, -119, -118, 88, -1, -85, 59, 24, 84, 52, 116, 6, -85, 68, -78, 112, -41, 34, 22, -62, -18, -103, -125, -73, -55, -15, -28, -3, -23, 52, 118, -114, 14, 69, 41, 12, -59, 78, -64, 86, 107, -118, 71, 75, -37, -57, -31, -107, -60, -17, -108, 31, 78, 91, -53, 112, -52, 86, -127, -81, 85, 81, -80, 62, 13, 7, -20, 38, -11, 75, -117, 7, -102, 94, 60, 8, -70, 1, -70, -93, 96, -35, 87, -26, -81, -14, -54, -67, -95, -32, 10, -124, 55, -19, 117, 79, 78, -107, 114, 4, -38, -107, -54, 85, 53, 97, 22, 5, -58, -95, 2, -40, -92, -124, -3, -128, 125, 55, -119, -110, -94, -90, -53, -116, -24, -2, 39, -35, 69, 5, 126, 85, 8, -38, -24, -84, 7, -109, -117, -16, -8, -51, 91, 18, 28, -16, 97, -109, -72, -15, 74, 76, 64, 36, 52, -122, -117, 49, -108, -102, 34, -66, -117, -41, -75, -36, 3, -99, -117, 79, -96, 65, 23, -95, -6, -42, 28, 13, 29, -95, -1, -20, 78, -91, -116, -66, -8, 82, 103, 105, -119, -59, 116, -98, 88, -1, -23, -51, -123, 99, 5, 33, 79, 50, -83, -84, -109, 123, -78, 29, 109, 34, 102, -62, 115, -34, 16, 32, 13, 40, 114, 23, -27, 96, -27, 22, 103, -68, -38, 49, -41, -81, -60, -43, 9, 25, 12, 75, 41, -75, -126, -30, -81, 8, -10, 77, 88, -116, -52, -57, -72, -105, 5, -84, 13, 3, -96, -100, -32, -4, 22, 44, -52, 48, -6, 30, 19, 75, -94, -94, -104, -46, -36, -87, -66, 59, -125, -34, 76, 34, 56, 67, 76, -64, 101, -75, 116, 20, 126, -88, -124, 43, 45, -3, -88, -6, 115, 75, -61, 56, -96, -44, -31, -60, 113, 84, -6, -127, -93, -81, -77, -52, 29, -35, 30, -40, -106, -6, 101, -115, -42, -21, 98, 126, 69, 47, 12, 72, -34, -89, 16, 88, -80, 58, -58, 31, -37, 122, 7, 98, 72, 104, -117, -66, 108, -4, 78, 49, 18, 51, -106, 117, -103, 110, -79, 93, 2, -99, -85, 93, 29, -109, -111, 56, 91, -48, 119, 58, -55, -58, 110, 46, 127, -66, 106, -9, 69, 0, -95, -35, 52, -79, 13, -14, 77, -13, -30, -30, 127, -107, 57, -52, 58, 67, -32, -57, 76, -46, -66, 92, -104, -99, 63, 53, -58, -50, -118, 54, -48, 27, 124, 36, -84, -111, -112, -22, -56, 120, -113, -102, -4, -44, -26, 49, 116, -107, 118, -26, -67, -87, -66, -68, 106, 88, -37, -57, -116, -76, 69, 28, 113, -107, -7, 103, 29, 94, 58, -94, 115, 25, 93, 3, 87, -20, -58, 79, 125, 110, -46, -72, 68, -99, 49, 40, 33, -108, 56, -81, 112, 29, -104, 7, -70, -34, -22, -60, -46, -2, 96, -125, 50, 110, -12, 8, 48, 112, 17, 109, -82, -66, -108, -124, -49, 73, 3, -14, -103, 110, 73, 39, 85, -45, -40, -7, -105, -116, 112, -49, -78, 63, 93, -49, 127, 33, -40, 71, 81, -119, 11, 26, -93, 71, -7, -26, -6, 71, 104, 116, -105, -43, -99, 61, -14, -98, 35, 102, -97, 89, -113, -48, 75, -110, 97, -11, -100, -104, -61, 40, 49, 34, -39, -97, -21, -28, 10, 127, 26, -61, -46, -20, 37, -108, 72, 10, 5, -49, 21, 2, -124, 21, 54, -111, -10, -42, -67, -93, 59, 33, -24, 107, -67, 108, 18, -72, -106, 71, -21, 73, 56, 78, -36, 70, 19, -99, -69, 9, 64, -17, 16, 43, -55, 89, 55, 117, -112, -29, 119, -105, 51, 15, 65, 28, 91, -74, 77, 94, 41, -90, -52, 117, 74, 74, -115, 62, -10, 28, -47, 82, 37, 114, 40, 35, 83, 106, 95, -65, -43, 101, -28, 95, -60, -69, -4, -25, 47, 9, -79, -100, 76, 74, 104, -72, -77, -65, -9, -10, 89, 64, -37, 48, -96, 16, 91, 14, 76, 42, 20, 124, 1, 98, 29, 84, 81, 43, -46, -88, -10, -50, -95, 48, 90, 59, 55, 70, -42, 18, -71, -40, 105, 121, -20, 26, -55, 118, 81, -113, -25, 37, -22, -10, 0, -64, -42, -22, -36, 120, -114, 70, -5, 92, -50, 35, 105, 117, 85, -47, -20, -57, 9, 52, -96, -100, 90, -117, -89, -73, 15, 6, 60, 89, 54, 127, 115, 112, -93, -58, -7, 64, 111, 116, 115, 101, 32, 125, 36, 63, -84, 68, 101, -124, 104, 20, -47, 57, 66, -32, -112, -77, -63, 2, 123, -75, 92, -8, 42, 83, -59, -15, -70, 41, -113, 33, 104, 42, -9, -65, 78, 92, 124, 64, 48, 94, -27, -63, 10, 82, 45, -105, 59, 99, 38, -63, -7, 99, 93, 38, 94, 95, 74, 59, -74, 67, 106, -70, -13, -39, 93, -22, 32, -96, -61, -123, 89, 85, 120, 118, 31, 95, 44, 53, 72, 40, -76, -111, -71, 53, -7, 62, -97, 77, 68, 11, -125, 25, 55, -63, -50, 109, 121, 122, 15, 26, 62, -100, 122, 127, 40, 86, 79, -50, 5, 31, 98, -35, 10, 6, -63, 43, -124, -77, -53, -105, -98, -70, -7, 26, -27, -64, 23, -9, -78, -7, -89, -80, 48, 12, -24, 37, -69, 112, 88, -47, 24, -14, -45, 79, -99, -74, -120, -73, 94, 24, 33, -17, 87, 61, -70, 54, 114, -32, -41, -86, 36, -109, -42, -107, 118, -47, 102, -88, -104, 56, 24, 21, 8, 76, 33, -84, 107, 74, 95, 85, -22, -76, 18, -82, 73, -14, 18, -52, -90, -67, -75, 46, -17, 60, 119, -5, -97, -37, 29, -82, 118, 122, 51, 37, -97, 63, -124, 26, -104, -4, -39, -111, -77, 81, 89, 91, 33, 73, 110, -70, 122, -102, 17, -109, -89, -4, 85, -12, 52, 40, -91, 101, -100, 61, 77, 7, 84, -11, -100, 21, -98, -36, -128, 60, -87, 26, 42, 32, -116, -69, 124, -79, -86, 99, -101, -51, 108, -88, 37, -119, -114, 39, 55, -57, 94, -105, 54, 109, 114, -16, -78, 12, 12, 37, -3, 97, -72, -76, 66, 24, 98, 66, 119, 35, 31, -116, 14, 104, 106, -35, -71, 6, -91, 85, 127, 126, -120, -27, 12, 56, -34, 77, -60, 70, -57, -15, 5, -48, 65, -76, 101, 99, 96, -65, -68, -87, 85, 15, -34, 106, -51, 44, -111, -111, -16, -119, 88, 95, 76, -112, -49, -19, 7, -39, -66, 121, 113, -25, -108, 86, 89, -21, -82, -126, -21, -27, 8, -37, -123, -64, -49, -30, 92, 78, 43, -116, -95, 81, 75, -114, -24, -72, -73, 107, -44, -49, 121, -22, 91, 100, -103, 117, -105, -16, 30, -72, -127, 122, 28, 76, 30, 62, 33, -27, 69, 79, 16, 9, -117, -23, -44, -123, -106, -115, 89, 50, -124, 104, -59, -26, -91, -124, 53, 31, 103, 14, 20, -103, 80, -79, 7, 122, 119, -126, 73, -71, -105, -10, 107, 67, 14, -111, -77, 100, -88, -16, -114, 118, 65, -32, -50, -68, 37, 118, -96, -103, -59, -2, -104, -128, -103, 104, -103, -100, -111, -59, -3, -13, -81, 17, -36, 14, -74, -40, -121, -15, -43, 28, 86, 53, 35, 53, 92, -108, 67, -77, -91, -79, -77, 29, 64, 30, -86, -28, 124, 19, -53, -54, -67, 94, -8, -18, 41, -87, -16, 114, 92, 70, 126, 37, -19, 60, -119, -36, -50, 27, 5, -82, 78, 97, -5, 13, -96, 84, 47, -21, -26, 125, -72, 29, 99, 97, -35, 11, 69, 77, -13, 10, 3, 54, -89, 43, 30, 117, 103, -20, -23, 67, 14, 65, -38, 72, -60, 73, 60, -23, 92, 19, 17, -63, 101, 42, -121, -121, 11, 46, 94, -20, 82, -42, 3, -90, -111, 39, -56, -17, 80, -71, 96, 6, 92, -99, 25, -20, 61, -25, 44, 107, -54, 114, 41, 34, 70, 45, 117, 127, -45, -4, 105, 3, 74, -1, -85, 24, 55, -4, 79, 101, -29, 10, 69, -113, -45, 104, -65, 51, -81, -48, -45, -78, -105, -18, 73, 11, 118, 73, -28, 18, 100, 28, 41, 47, -56, 64, 14, 100, 42, -89, -34, -17, -31, -42, -99, -85, 54, 29, -19, 15, -60, -122, 66, -29, 22, 34, -6, 5, -17, -42, -26, 80, 125, -60, 8, -92, 73, 121, 17, 60, 22, 93, 18, 40, -54, 19, -42, 103, -93, 41, 25, 37, -60, 57, -88, -99, 3, 55, -128, -16, -27, -120, -101, 47, 63, -14, 115, 39, -91, -69, 1, 100, -3, -58, 102, 103, -126, 126, 40, 11, 110, 115, 33, 47, -51, 27, -83, -127, -60, 16, -80, -46, 71, -54, 3, -96, -109, 69, -8, 53, 127, -5, 41, 33, 66, -75, 21, -48, 91, -108, 116, -9, -93, -34, -76, 64, 5, -101, 53, 88, 68, -61, 0, 84, 95, 25, 83, -1, 54, 88, -47, 100, -71, -87, 64, 65, 52, 66, 55, -24, -98, -38, -104, 76, -78, 55, 127, 117, 39, -87, 33, 82, -106, 41, -96, 3, 78, 112, -43, -28, -9, -122, 15, -82, -112, 117, 79, -64, 113, 97, -4, -39, 91, -99, -47, 11, 33, -43, -118, -107, 63, -8, -100, 86, 67, -47, 25, 74, -35, -94, 77, 52, -89, 76, 115, 26, 47, 77, -127, -108, 9, 126, -84, -58, 91, -55, -128, 83, 66, 75, -74, -119, -105, -25, -7, -69, 62, -125, 106, -112, 41, 4, -103, 50, 76, -98, 26, -84, -25, 39, -1, -84, -95, -46, -107, -92, -42, 100, 45, -109, -51, -68, 24, 14, 85, -60, -41, 93, -95, -105, -60, 54, -46, -116, -79, 50, -55, 114, 90, 67, -50, -121, -14, 88, -32, 59, 14, 108, -62, 59, 106, 3, 34, 35, -28, 49, 21, -51, 46, -10, -47, 35, -90, 58, 40, -18, 70, -80, -30, 97, -77, 77, 126, -34, -12, 43, -33, -116, 107, 47, -74, -80, 25, 65, -23, 58, -88, 54, 97, 69, 65, 22, 25, 18, -89, 125, 69, -17, 17, 101, -33, -41, 82, 23, -18, -104, -23, -14, -73, 17, 59, 92, 23, 80, -109, 33, -29, 84, -88, 23, 110, 96, -82, -28, -21, -1, -55, 39, -42, 111, -13, 63, 12, -107, 38, 78, 65, 91, -73, 110, 127, -57, -63, -59, -62, 108, -65, -105, 71, 4, 115, -116, 92, -100, -106, 103, -2, 60, 31, -25, -94, 81, -118, 75, 99, -18, -36, 70, 93, 63, 38, -109, 74, 94, 83, 61, -9, -107, -6, 14, 82, -65, -72, 8, -36, -100, 116, 81, -72, 68, 35, -11, -60, 108, -116, 54, -48, 124, -120, -12, 19, -126, -105, 84, 47, 73, 115, 39, 105, -22, -44, -86, 85, 89, 57, 39, 13, 82, -52, 94, -106, -93, -86, 68, 71, 10, 95, 85, 112, 107, 91, 64, 52, -101, -34, -26, 126, 49, 43, 122, 37, 55, 25, -128, -46, -100, -51, 44, 47, -58, 92, 17, 99, -88, -111, -51, -66, 41, 93, -9, -104, -119, 45, -36, -124, 110, -84, -10, 100, 116, -15, 20, -2, 18, 75, -74, 107, -89, 12, 125, 18, 92, 58, 23, 47, 70, 9, 60, -34, 21, -12, -105, 11, 99, 95, -27, -105, -99, -91, 66, 3, -88, -64, 94, 7, 61, -89, 16, -59, 60, 11, 37, -37, 82, 17, 15, 46, -14, 31, 33, -99, -94, 14, -91, 118, -108, -34, 13, 61, -20, 55, -97, 59, 66, -3, 8, 55, 67, 7, 119, 104, -121, -102, -13, -113, 17, -52, 25, -44, -123, -30, -67, 86, -80, 27, 121, -101, 6, 84, -11, -25, -113, -92, -80, 22, 26, -46, -21, 54, 13, -45, -18, -95, 47, 106, -81, 118, 35, 74, 88, 87, 17, 36, 39, 55, -33, -68, -50, 103, -103, -24, 123, -78, 114, 71, -36, 79, 35, -72, -62, -57, 18, 91, -43, -122, -46, -77, 27, 105, -6, 99, -42, -3, -94, 31, -65, 41, 27, -66, -127, -91, 10, 3, -65, 17, 68, -3, 85, 5, -1, -73, -97, 99, -62, -105, 17, 25, -81, -46, -110, -102, 86, 27, -34, -50, 124, -85, 52, -62, 51, -27, -24, -79, 19, -88, -44, 58, -111, 104, 116, -6, -29, 72, -94, 52, 84, -5, -71, 10, -119, -91, -11, 60, 74, 53, -27, 39, 106, -114, -91, -46, 67, -103, -127, 53, -78, -114, -103, 96, 90, 59, -86, -21, 41, 91, 67, 73, 58, -39, -80, 2, -38, 10, 11, -107, 58, -107, -50, -32, 126, -123, 95, -18, -37, -75, -28, -73, 37, 8, 64, 21, -37, 14, -32, -9, -28, -48, 14, -91, -30, 117, 47, -44, -87, -37, -21, -49, 99, -14, 37, -30, -87, -96, -32, -115, -83, 15, -42, 127, 101, 9, 57, 31, -29, 19, 52, -42, -89, -92, 70, 118, -42, 33, -90, -68, 104, -90, 94, -105, -38, 48, 57, 90, -31, 84, 67, 19, 78, 33, -18, -114, -69, 101, 113, 24, 5, 102, -26, -100, 117, 27, -113, -80, 73, -40, -60, 69, 120, -78, -23, -114, -9, -68, -123, 76, 39, -116, 41, -120, 119, -24, -2, -13, -28, -6, 70, -95, -122, -17, -117, 66, 19, -67, 99, -80, -69, -6, -20, -15, 43, 33, -32, 112, -25, -31, 84, 15, -96, -80, -60, 81, 26, -40, -58, -19, 20, 65, -57, 46, 46, -114, 73, 88, -96, -67, -19, -70, 54, 76, -107, -29, 97, -121, 113, -57, -69, 24, -67, -19, 55, -40, -29, 28, -112, 53, -89, 116, -21, -34, -50, -118, 65, -27, -89, 43, -102, 77, 117, 104, 102, 61, -101, 18, -74, -67, 31, 116, -89, 116, -62, -36, -38, 84, 111, 110, 90, 104, -104, 70, -92, 17, 54, 82, -70, 64, 82, -122, -38, 23, -15, -36, 36, 81, 122, 26, -7, 104, 108, -42, 12, -41, 32, 33, -104, 68, -95, -109, 32, 119, -20, 99, -70, 70, -45, 10, 80, 72, -14, 111, 44, 46, -74, -36, 119, 56, -38, 90, 75, -116, 99, -125, -54, 81, 41, -102, 60, 15, 67, -31, -94, 122, -17, 121, -8, -23, -42, -118, 111, -110, -118, -73, -47, 120, -79, -81, 64, 9, -62, 76, -59, -6, -60, -113, 19, -44, 2, -97, -80, -48, -84, -32, 38, -107, -75, -112, -98, -28, -3, 123, -112, -5, 79, 72, 97, 80, 65, -105, -18, -61, 44, -16, 75, -67, -2, -83, 13, -38, 122, -4, 73, -11, 76, -15, 27, 59, -82, 116, -48, -12, -111, 81, -27, 124, 106, -73, -110, 9, 74, -119, -95, -91, -42, 69, 61, -89, 80, 29, 95, -84, 83, -124, 112, -90, 43, -92, 68, -48, -94, 93, -13, 72, 6, 88, 112, -93, 58, 68, 2, 41, 47, -41, -13, 48, -6, -70, -48, -17, 6, 26, 113, -6, -113, -18, 0, 48, -19, -53, -79, 11, 33, 49, -104, -72, 42, 37, -55, 73, -17, 48, -16, 26, -79, 50, 33, -48, 108, -126, 118, -18, -2, -122, -68, 24, 32, -103, 36, 79, 65, 45, 103, -23, -43, -41, -57, -25, -34, 13, -86, 120, 89, 105, 63, 125, -53, 56, 40, 123, -8, -87, 59, 123, -19, -7, -108, 86, -49, 75, 110, -6, 3, 6, -13, 91, 80, 34, 41, 18, -2, 31, 89, -93, -103, 9, 72, 81, -34, 14, -64, -79, 43, -75, -84, -20, 55, 9, 80, -102, -17, 87, -45, -66, -15, 108, -47, 39, 85, 118, 76, -105, 76, -124, 73, 82, -126, -86, 29, -7, 108, 122, 51, -35, 83, -49, -115, -71, -113, -56, -38, 95, 110, -102, -125, -53, -8, -117, 102, 117, -7, 60, -35, -38, 105, -79, -110, 42, 91, -72, -37, 62, -76, 45, -98, 47, -88, -12, -70, 42, 17, 33, 92, -78, -81, 21, 57, 126, 5, 13, 27, -19, 22, 21, -56, 31, 21, 73, -122, 57, 71, -67, -110, 28, 27, -71, 126, -81, 121, 24, 79, 66, -101, -29, -94, 89, 54, 45, -64, 103, 110, 83, 59, -103, -106, -94, 8, 71, 44, 91, 66, -91, -57, -117, 9, -3, 109, -20, 64, -45, 32, -84, 48, 11, -44, -20, -75, -113, 87, 109, 113, -108, 118, 23, 55, 13, -44, 39, -91, 74, -54, -88, 74, -46, 2, -68, 43, 5, 97, -103, -25, -15, -81, 61, -24, 113, 14, 118, -90, -72, 34, -57, 57, 44, -31, -7, -11, 37, -119, 46, -45, -16, -84, 30, 33, -111, -99, 119, 81, 109, 114, -56, 117, -77, -120, 118, 114, 3, 107, 80, -128, 23, 69, -69, -50, -128, 10, 116, -49, 90, -2, 18, 126, -78, -27, 64, -38, 44, -124, 57, -124, 123, 8, -87, -97, 23, -25, 101, 123, -50, 85, 25, -68, 77, -111, -110, -42, -65, 104, -101, 12, 100, 127, -95, -26, -23, 98, -62, -91, 10, -43, -62, 32, 123, 89, -128, -128, 12, -88, 121, 64, -64, -66, -83, 105, 54, 21, -88, 60, 14, -27, 83, 19, 25, -70, -95, 95, 56, -45, 127, 61, 114, -100, -34, 81, -38, -29, -65, 104, -23, -107, -19, -51, -15, -5, -91, -78, 39, -79, 29, 61, 5, -69, 31, -37, -96, -13, 32, 123, 72, -62, -22, 40, -128, 119, 11, -120, 118, -10, -15, 63, 76, -9, -8, -116, -108, -3, -100, -16, -74, -3, 87, 125, 7, 40, 98, 55, 85, 83, -99, 99, 16, 1, 39, 6, 110, -104, 112, 77, 80, 109, 53, 124, -31, -50, -24, 125, 111, -58, -80, 43, 5, -73, 107, -58, 27, -18, -67, -58, -108, 81, 21, -108, 52, -90, 24, -25, 10, -107, -109, -56, 60, 35, 97, -106, 121, -68, -21, -72, -104, -47, 11, 68, -15, -88, -47, -117, -61, 27, -110, 86, -126, 59, -99, -34, 126, -11, -97, 49, -107, 62, 4, -86, -104, -54, 50, -7, 66, -25, 41, 92, -5, -5, -73, 35, 57, 126, 51, -52, 24, -29, -10, 24, -90, 72, 2, -50, 27, 64, -33, -110, 100, 109, -121, -90, 15, -125, -45, 100, -92, -52, 37, 49, 86, 86, 125, 27, 49, 110, -122, 102, -100, 59, -17, 90, 94, 43, 37, 64, 56, 86, -104, 110, 5, 55, 6, -76, 117, 46, 62, -106, 123, -77, -2, -54, 105, 96, 86, -10, -21, -75, 25, -80, 34, 119, -77, 68, 34, -69, 59, -51, 23, 118, 95, 73, -114, -7, 64, 23, 17, -101, -63, 23, -119, -110, -51, 21, 122, -90, 122, 94, -6, -61, 15, -28, -106, 99, -78, 61, -11, -47, 120, -53, 116, -14, 125, -54, 36, -63, 101, 12, 19, -111, -96, 58, -69, 73, -39, -47, -56, 34, 30, 1, -62, 76, 52, 89, 45, -54, -108, -63, -86, 83, -54, 79, -50, -50, 76, 9, -4, 71, -39, 5, 4, -32, -71, 4, -93, 95, -63, -116, 7, 52, 50, -57, -31, 24, 127, -56, -25, 60, -115, -65, 124, 67, -60, -96, -51, 59, 90, 103, -48, -81, 22, 124, -41, 126, 40, 12, -19, -96, 101, -45, -33, 108, -27, -57, 126, -67, -62, -16, -122, -31, -70, -105, 115, -102, 103, -11, 9, 7, -17, 6, -27, 79, -22, -97, -103, 83, 35, 81, -124, -108, 115, -36, 69, 102, -102, 88, -104, 86, 93, -128, -29, -87, 18, -39, -114, -35, 10, 125, 63, 99, -25, 50, 41, 85, 11, -39, 61, -88, -123, 124, 123, 2, -33, -37, 85, 20, 37, 126, -73, 88, 12, 86, -39, 105, 23, 60, -98, 31, -128, 34, 77, -106, -94, -64, 37, -33, -61, -32, -3, 24, -115, -5, -56, -100, 125, -66, -103, -12, -6, 27, 73, 93, -4, -90, -128, 85, 98, -115, 85, 69, 102, 94, 18, 105, -13, 72, -51, 47, 86, -126, 106, 78, -51, 66, -113, -99, -112, -79, -13, -14, -107, -95, 8, -116, -3, 104, 118, -77, 23, 5, -92, 126, -75, 99, -55, 14, -45, 42, 93, 62, 6, -28, 10, 123, -127, -31, -78, -22, -110, 85, 17, 93, 58, -94, -96, -15, -31, -55, -2, 14, -59, -5, -107, 67, -41, 22, 47, -38, 74, -58, 50, 17, -54, 61, 49, 13, 127, 55, -110, -87, 21, 125, 121, 78, -89, -53, 91, 120, 70, 32, -35, -99, 110, 28, 101, -40, -53, -4, 127, 16, 56, -111, 42, 41, 28, 77, 32, -89, 16, 82, 51, -23, 29, -64, -86, -115, 99, 42, -61, 47, -103, -74, 123, 66, 58, -111, 62, -7, -34, 40, 44, -96, -122, 97, -15, 123, -43, -46, -59, 92, -74, -86, -111, 7, 56, 17, -90, -49, -7, 70, -48, -48, -16, -74, -78, 37, 36, 45, -52, -117, 71, 107, 119, -77, 127, 21, -24, -48, 98, 42, -55, 124, -122, 49, 58, 25, 106, 73, 59, -108, -61, 113, 63, -95, 85, -23, -78, -15, -83, 85, -123, -21, 109, 94, -36, 53, 120, 56, -66, 29, -82, 8, 62, -57, 126, 26, -35, 91, 60, 47, -49, 109, -123, 6, -128, 74, 75, -15, -32, 88, 18, -125, 42, -9, -115, 9, 31, 29, -46, -44, 0, -89, -4, 13, 103, -43, 115, 84, 28, 41, 37, -77, 21, -110, 117, 6, 38, -78, 45, 34, 37, -27, -93, -28, 69, 111, -19, -110, 31, -32, 124, 42, -65, -53, -94, -34, -47, 2, -116, 104, -117, 11, -120, -56, -42, 47, 36, -67, -78, 55, -60, -34, -39, -50, 16, 84, 36, 97, -118, 1, -42, 42, 42, 59, -92, 46, -126, -24, -126, -73, -82, 54, -39, 49, 52, -109, -36, -10, -108, -76, 5, 93, 25, 67, 118, 77, 119, -42, -91, 75, 99, 28, 51, -105, 70, 113, 0, -125, -37, 2, 18, -21, -15, -37, 33, -4, 0, 73, 28, 89, -17, -124, -52, 56, -101, -5, 29, -69, 29, 19, -67, 51, -121, -35, 55, -34, 31, 32, -13, 107, 65, 71, -34, -1, 12, -48, 49, -127, -54, -48, 73, 101, -48, -43, 123, 22, 103, -123, 49, -40, -66, -108, -74, 57, 107, -101, -82, -47, -108, 48, 118, -37, 70, -5, 0, 17, -49, -86, 43, 94, 55, 80, 114, 6, -30, -46, -39, -91, 38, 50, -51, 81, -59, -77, 76, -87, -44, -36, -41, 22, 127, 38, 107, 121, 21, -71, -95, -78, 82, -26, 16, 33, -83, -125, 63, 30, 96, 57, -53, 81, 47, 49, 78, -111, 14, -70, -34, 65, 118, -32, 89, -107, -106, -46, -78, 58, 123, -1, 99, -30, -24, -58, -107, 123, 87, -122, 34, -112, 2, -115, 18, 84, -111, 116, -8, -36, -52, 51, 7, 96, -61, 21, 9, 45, 54, 75, -34, -87, -116, 14, -43, -41, -99, -23, 8, 124, -16, 114, -6, -128, 65, 55, -64, 55, 91, -102, 58, -88, 30, -7, 47, 46, -8, -19, -84, -84, 126, -19, -38, 41, 100, 109, -43, 25, -69, -111, 85, -97, 38, 26, -23, -84, 16, -56, -123, 75, 124, 117, -79, 105, -7, -58, 0, 53, 114, 2, -25, 20, 53, 113, -75, -3, -108, 117, -15, -49, -90, 0, 32, 33, 53, -49, 105, -72, 74, -86, 122, 103, -111, 79, 81, 111, 60, -46, -9, 50, -15, 0, 10, 46, -45, 55, -51, 94, -87, 53, -48, 52, -100, 57, 30, -28, -63, 71, 96, -87, 12, -92, 123, 42, -88, 38, 17, -69, -36, 114, -99, 26, 16, -16, -56, -112, 64, 117, -101, -29, -33, -105, 101, 19, 80, 51, -14, -114, 67, -86, 34, -99, -73, -88, -62, -37, 127, -114, 99, -104, -92, -80, -66, 22, -126, -8, -54, 27, 59, 55, -66, 104, 125, 45, -79, 92, -100, -123, -40, 73, -60, 120, -42, 3, 109, 15, -101, 29, 108, -66, -34, -45, -116, -93, 41, 1, 77, -16, -18, 85, -1, 20, -59, -106, -7, -60, 69, 122, 31, 16, 7, -15, -56, -12, -91, 98, -42, 113, -82, -98, 65, 106, -22, 78, -67, 93, 81, 115, 78, -67, -128, 110, -102, -76, 22, 27, 106, -11, -113, 51, -6, -91, -127, -112, 44, -2, 38, 87, 11, 116, 121, -80, 20, -84, 41, -12, 30, 111, 50, 94, 53, 111, -96, 115, -19, 19, 39, 46, 13, 98, -67, 48, -43, 66, 71, 104, -47, 10, 108, -57, -17, -19, 117, 108, 114, -17, 25, 56, 42, -120, -123, 54, -59, 22, 11, 54, -10, -70, 32, 107, -57, -116, -34, 76, -28, 3, -64, -29, 119, -59, 65, 39, 101, -72, 28, 23, 3, 47, 15, 75, 9, 84, -21, -96, 98, 110, 74, 43, 107, 23, 66, 28, 13, 84, -67, -41, -117, 109, -111, -118, 64, 33, 11, 51, 67, 21, 11, -109, 124, 22, -36, 83, 56, 16, 31, -111, -22, 106, -108, -81, -106, -88, 120, -24, -4, -69, -54, -77, 59, 111, -67, -26, -50, 71, -56, -112, -5, -105, -30, 44, 123, 12, 2, -86, -60, 104, -88, 109, -127, 103, 100, -31, 92, 59, 63, -93, -78, 43, -97, 0, -52, -11, -13, 59, 18, 78, -112, 37, 19, -3, 79, 69, -31, 74, 22, 92, -57, -113, 114, -119, -80, 31, -92, 18, -106, 29, -36, -8, -36, 31, -5, 39, -68, 90, 90, 114, 98, 87, 117, -18, -95, 39, -71, 94, 75, -6, -80, -123, -18, -126, -91, -47, 3, 71, -15, -87, 112, -83, 33, -22, -75, -66, 105, 84, 0, 80, -127, 93, -26, -42, -82, -84, 20, 62, 7, -10, 97, -33, -99, 2, 100, -86, 49, 108, -6, 113, -26, -89, -70, -85, -100, 47, 99, -108, 11, -26, 111, 79, 45, -10, -41, 102, 13, -6, 93, -79, -15, 54, 11, -125, -1, 93, -92, -115, -83, -70, -64, -104, -16, -12, -34, -74, -99, 97, 36, -59, -108, 62, -35, -37, -42, 14, -64, 42, -16, 110, -15, 86, -111, -95, -49, 7, 123, -38, -33, -126, 79, 114, 107, -1, 89, -112, -15, -87, -69, 60, -101, -89, -115, 97, 89, -9, -121, -119, 48, 16, 4, -27, 101, 112, -74, -49, 104, -6, -122, -36, 89, 51, 65, -72, 115, -78, 92, -24, -64, -34, 126, -1, 114, -53, -114, -108, 90, 33, 59, -9, -115, 125, -3, -68, 88, 11, 46, -100, -17, 85, 59, 109, 88, 55, 68, -41, -1, 72, 85, 13, 7, 14, -84, -121, 101, 55, -49, 55, 100, -50, 75, 70, 42, -126, 82, -125, -37, 10, -56, 62, -21, -3, -123, -100, 39, -38, -49, 12, 56, -11, 91, -114, 14, 74, 110, 124, -82, 60, 14, 3, 88, -126, 45, -91, -35, 111, 100, -51, 81, 41, -76, 18, -50, 114, -7, -127, 98, -33, -53, 22, 96, -101, -13, 28, -42, -100, 21, 104, 28, 100, -18, 26, -37, -36, 13, 102, 75, -87, 47, -76, 122, -57, 73, -86, -77, 58, -35, 24, -10, 59, 22, 6, -47, -122, 45, -66, 68, -121, -94, 38, -12, -69, 9, 14, 59, -98, 66, 36, -70, 39, 116, 72, 99, -106, -5, -60, -36, 103, -122, -44, -87, -35, -119, 115, -74, -70, 40, -15, 79, 89, -26, -67, -9, -88, 104, -128, 46, 97, 86, 24, 101, -75, 30, 84, 43, 78, 32, 99, -5, 90, -62, 31, -125, 0, 113, -126, 92, -71, 85, -83, -51, -108, -8, 35, 0, 56, -13, 26, 102, -34, -82, 93, -66, -57, -10, -18, -89, -110, -119, 117, 121, 32, -71, 68, -101, -99, 8, -39, -115, 120, -123, -38, 119, -73, 112, -11, 100, -32, 112, -3, 10, 20, -9, -121, -6, -105, -41, -84, 6, -93, -29, 35, 6, -3, 117, 95, -71, -126, -24, 89, -110, -72, 45, 82, 91, 11, -74, -107, 101, 2, -63, -23, 119, -84, 26, -98, 7, -127, -25, 11, 56, 32, -62, 62, 31, -31, -112, 60, 57, -45, 16, 3, -71, 63, 121, -122, 95, 112, -90, 31, -33, -91, -31, -97, -73, -52, -22, -87, 5, 0, -96, 123, -112, -76, 45, -74, 15, 74, 106, -109, -128, -91, -54, -30, 92, 67, 94, 52, -111, 7, 26, 94, -48, -47, 53, 83, 23, 13, -97, -89, -44, -56, -115, 122, 6, -88, 3, -87, -71, -96, -78, -121, -118, -118, 81, -20, -82, 29, 24, -33, -73, -38, 76, 58, -36, 31, -37, 38, -63, -121, -13, 58, -42, -117, -107, -20, 119, -19, 50, -59, 95, -46, -38, 104, -43, -58, -111, 67, -56, -42, 7, 50, -89, 33, -96, -93, 35, 114, 119, -110, -75, -128, -128, 35, 114, -102, -22, 88, 26, 98, -122, 57, 12, -40, -101, 48, -61, 113, 16, -84, -36, -63, 104, -33, -44, 66, -124, 3, 86, 110, 104, -121, 40, -73, 3, 6, 98, 110, 50, -114, 29, -56, 111, -50, -43, -26, -72, 108, 99, -46, -14, -59, -16, -106, 98, 61, -111, -108, 1, 40, -13, 123, 106, -124, 59, 81, -94, 116, 107, -97, -8, -22, 89, 101, -16, -32, -102, 29, -71, 91, 0, -8, -79, -55, -68, 60, 114, -126, 21, 113, -110, -17, -121, -83, -18, 23, 46, 86, -54, 117, 10, 55, 77, -71, -67, -116, -104, 117, 15, -105, 8, 15, -108, -85, 115, 76, 53, 60, -109, 38, 19, -50, -112, 7, 8, 107, -110, -27, 9, -98, 126, 108, 72, -122, 44, 22, -73, -117, -20, 26, -85, 49, 83, 70, 72, 114, 85, -28, -6, 122, 49, -63, 38, 79, -83, 4, -86, 105, 21, -113, -70, 54, 60, 37, 101, -67, -48, 35, 37, 29, 110, 121, -18, -73, 80, -56, -29, 85, 85, 52, 17, -126, 32, -118, 73, -77, -23, -83, 27, 98, -97, 95, -63, 75, -92, -66, 18, -120, 109, -49, 73, 113, 52, -17, -12, -127, -31, -93, 77, 85, 57, 112, -88, 46, 102, 26, 84, 35, -120, -119, -105, 53, -14, 83, -110, 43, -94, -64, 75, -48, -30, -102, -39, -58, 80, -76, -82, 120, -93, -102, 85, -121, 12, -84, -10, -11, -49, 93, 104, -8, -17, 28, 39, -32, 100, 99, 80, 72, -44, 20, 37, 7, -22, -28, 109, 88, 52, 66, -80, -69, 30, 40, -11, -88, -101, 97, -39, 33, -23, 89, 29, 37, -60, -71, 12, 72, 31, -41, 121, -82, -48, -1, 76, -18, -39, -23, 60, 30, -118, -99, 43, 127, 50, -51, -65, -82, -128, -76, 63, 22, -43, 66, -14, 112, 10, 81, 10, -93, -30, -36, 70, -10, -25, 8, 24, -82, 72, 115, 38, 11, 69, -102, -75, -23, 34, -72, 24, 97, 66, -123, -16, 43, 80, -41, -63, -58, -76, -64, -100, 68, -68, 79, -78, -39, 16, -19, 102, -56, -121, -39, -121, -7, 27, -83, 103, -79, -17, 87, 24, 51, -108, 55, 39, 64, 54, -110, -12, -87, -22, -39, -116, -116, -17, 123, -26, -34, -18, 111, -14, 74, 17, 95, 68, 14, 78, 61, -12, 19, 36, 24, -87, -78, 11, 15, -13, 41, -21, -29, -38, 31, -44, 95, -77, -86, 120, 104, 68, 61, 1, -71, -75, -35, -14, 32, 75, 27, 65, 3, -26, -23, -2, 106, 83, 38, 59, -37, 32, -53, -99, -26, 39, -90, 10, 53, -67, 75, 127, 89, -43, 96, 113, -86, 22, 116, 16, -9, 90, -97, 88, 96, 8, -69, 97, -19, 74, 73, 12, 68, 84, -23, 98, -26, 126, 34, 83, -78, 20, 120, -10, 93, -126, -102, -84, -121, -34, 62, 19, -33, -70, 10, -46, -6, 36, 18, -7, -44, -69, 123, 21, -67, -7, 24, 38, -53, -17, -14, -22, 76, 124, 107, 114, -74, 62, 13, 93, -59, 19, 25, 17, 119, -76, 103, 6, 8, 94, 120, -30, -61, -66, 28, 82, 7, -98, 59, -122, 39, 60, -91, 10, -4, -2, 127, -88, -114, 64, -113, 60, 2, -31, 40, 80, 3, -102, 114, -95, -95, 77, -43, -72, -75, 39, 82, 60, -69, -74, 99, -69, -103, -66, -71, -96, -14, 37, 16, -10, 114, 61, -97 );
    signal scenario_output : scenario_type :=( 127, 127, 127, 1, -6, 81, 127, 127, -79, -128, -128, 48, 127, 127, 16, -109, -128, -48, 7, -17, 73, 127, 127, 127, 127, 127, 24, -128, -128, -1, 0, -76, 38, 127, 127, 33, 73, -24, -128, -32, 127, 127, -64, -2, 52, 127, 127, 127, -128, -128, -59, 49, 85, 55, 103, 27, -16, 127, 127, -80, -86, -123, -128, -128, -66, -28, 38, 127, 127, 127, -128, -128, -80, 127, 127, -58, -128, -70, 127, 127, -69, -66, -16, 16, 33, 127, 127, -81, -128, -109, -58, -54, -128, -128, -80, -29, -21, -58, -128, -128, -71, 127, 127, 127, 127, 44, -128, -128, -128, 44, 45, -128, -128, -95, 127, 96, -128, -128, -32, 80, 50, 80, 127, 127, 81, -128, -128, -107, -26, -76, -88, -128, 45, -34, -128, -128, -116, -24, -49, -68, -121, 127, 127, 123, -79, -33, 127, 127, 127, 87, 58, 0, -60, -33, 42, 66, 45, -1, -128, -102, 15, 127, 127, 53, -128, 36, 127, 127, -80, -128, -128, -55, 6, -28, -26, 33, 54, -36, -79, -32, 16, 2, 15, 0, 91, 85, -59, -128, -128, 7, 127, 127, -48, -128, 36, 127, 95, 16, 68, 127, 109, -16, -123, -128, -128, 66, 113, 24, -81, 127, 127, 127, 127, 127, 127, 127, 127, 102, -128, -128, 12, 36, 71, 123, 100, -97, -128, -128, -88, 32, 79, 127, 127, -52, -128, -128, -63, 88, 112, 10, -128, -128, 127, 106, 81, -13, -13, -128, -128, 38, 127, 127, 114, -128, -128, -128, 53, 127, 127, -53, -53, 23, -7, -128, -128, -58, 7, -81, -65, 86, 114, 24, -78, 1, 18, -128, -128, -128, 26, 127, 127, 90, -27, -128, -128, 127, 127, 127, -128, -128, -128, 91, 111, 1, -128, -53, 33, 76, -128, -122, 123, 127, 127, 71, -128, -128, -128, -28, -1, 96, 127, -21, -128, -1, 6, -128, -128, 28, 127, 127, 127, 127, 127, 8, -128, -128, -27, -31, -78, 65, -53, 103, 127, 34, -128, -128, 37, 127, 127, 16, -22, 124, 127, 127, 103, 44, 13, -59, -128, 11, 127, -15, -23, -76, -43, 65, 127, 127, 15, -36, -100, -55, 0, 7, -128, -128, -124, 102, 63, -92, -119, -128, -54, 36, 127, -36, -38, -15, -71, -128, -128, -78, -18, -44, -52, -128, -128, -6, 102, 12, -128, -107, -65, -36, -16, -128, -128, -113, 11, 127, 80, 44, 98, 127, 15, -1, 23, 38, -128, -128, 36, -6, 53, -21, -66, -128, -50, 17, -119, -128, -128, -86, -128, -128, -128, -57, 127, 127, 127, -128, -128, -128, -69, 93, 127, 127, 127, 63, -86, -111, -12, -60, -108, -88, 1, 18, 127, 63, 127, 127, 127, 127, -33, -103, -12, 21, -15, -38, 127, 127, 124, -128, -128, -128, -37, 74, -71, -128, 17, 127, 127, 127, -18, -95, 22, 127, -101, -128, -68, -16, -36, 32, 127, 117, 21, -128, -128, -13, -70, -22, 15, -128, -128, 69, 127, 59, -26, -90, -128, -128, 42, 108, 63, 127, 127, 127, 127, 76, -2, -128, -128, -128, -128, 54, 127, 127, -123, -128, -66, 1, -28, -128, -128, -15, 127, 127, 68, -114, -128, -128, -68, -5, 85, 121, 97, 121, 127, 57, -7, -34, 45, 79, 127, -49, -118, 73, 127, 127, -22, -58, -53, -57, -128, 36, -57, -26, 127, 127, 103, -101, -128, -128, -128, 11, 127, 127, -18, -81, 2, 111, -50, -98, -58, -12, 38, -92, -32, -118, 86, -22, -128, -128, -38, -128, -128, -106, 127, 127, 127, 96, -11, -128, -68, 80, 11, -128, -88, 21, 31, 127, 127, 127, 74, -100, -128, -128, 42, 76, -101, -128, -95, 127, 127, 127, 12, 5, 36, 100, -128, -23, 65, 127, -71, -93, -128, -128, -128, 127, 127, 90, -86, -112, -12, 127, 127, 127, -17, -128, -103, 127, 127, -39, -121, 2, 127, 127, 127, -7, -128, -64, 127, 122, -18, -128, -128, -128, -128, -68, -45, -16, 127, 127, 78, -64, 1, 91, 103, 85, 88, 71, -109, -128, -65, 48, 127, 2, -107, -76, 127, 123, -95, -128, -42, 127, 127, -38, -122, -128, -21, 96, 127, 52, -42, -124, 49, 87, -11, -60, 123, -39, -128, -128, -75, -79, -101, -12, -106, -58, -29, 53, 106, 108, -108, 34, 101, 92, -128, -128, -97, 71, 112, 17, -6, 3, 90, -43, -113, 10, 114, -6, 122, 127, 64, -128, -117, -52, -26, -107, 38, -50, 24, -128, 10, -63, 8, 16, 127, -24, -128, -128, 45, 127, 127, 107, -38, 27, 127, 127, -128, -107, 101, 127, 127, 127, -12, -74, 21, 127, 55, -45, 32, 92, 68, 39, 16, -22, -128, -128, -26, 127, 127, 17, 127, 127, 127, 127, 127, 106, -118, -128, -128, -18, -47, -13, 123, 127, -57, -58, -108, 33, 7, -96, -128, 76, 114, 122, -76, -128, -128, -75, 75, 127, 127, -91, -128, -92, -88, 29, 116, 127, 127, -11, -128, -128, 101, 127, 127, -8, -122, 23, 127, 127, 127, -34, -128, -43, 127, 127, 22, -128, -128, -114, -22, 18, -128, -128, -70, 3, -59, -48, 127, 109, -70, -128, -45, 127, -26, -124, -49, 127, -44, -128, -112, 55, 118, 88, 127, 127, 127, 55, 34, 10, -49, -103, 91, 127, -98, -128, -128, -128, -128, 39, 127, 127, -124, -127, -16, 127, 106, 102, 66, -128, 6, 127, 127, -2, -48, -128, -59, -108, 0, 32, 43, -128, -10, 127, 127, 117, -74, -100, 127, 113, -128, -128, 76, 45, -106, -98, 109, 109, -5, -58, -128, -128, 75, 127, 87, -50, 10, 107, 127, 127, 127, 127, 76, -96, -90, 37, 119, -11, -13, -79, -128, -128, 11, 122, 53, -36, -119, -37, -85, -37, 127, 111, 45, 127, 111, -128, -128, -128, 18, 103, 93, -8, 127, 127, 127, 127, 127, 63, -128, -128, -81, 10, -128, -128, -128, 13, 127, 127, -108, -128, 18, 127, 127, 16, -128, -128, 87, 127, 92, -128, -128, -128, 0, 127, 127, 75, 49, 91, -1, -108, -128, -128, 22, 127, 127, 127, 127, -112, -128, -33, 127, 118, -128, -128, 95, 78, -124, -128, 127, 80, -128, -128, -128, -128, -121, -7, -128, -128, 45, 127, 127, 43, -128, -128, -109, -128, -128, -121, -21, 60, -12, -128, -128, -128, -63, 12, 127, 127, 127, -23, -128, -128, 102, 127, 88, -113, 1, 127, 127, -50, -128, 7, 127, 127, 127, 127, 75, -96, -128, -113, 100, 74, 48, 127, 127, -79, -85, 73, 127, 50, -44, -128, -128, -57, 127, 127, 127, -68, -128, -31, 127, 127, 2, -68, 91, 127, 127, -79, -128, -128, 58, 22, -117, -98, 96, 70, -90, -90, -13, -42, -128, 0, 127, 127, -123, -93, 21, 127, 75, 127, 113, 38, -68, 66, 0, -58, -90, 3, 18, 127, 127, -91, -128, 16, 127, -33, -128, -59, 38, 119, 55, 75, -128, -128, -128, 16, 90, -27, -128, -128, -128, 75, 118, 26, -128, -91, 127, 127, -91, -128, -128, 91, 127, 127, 87, 127, 127, 36, -5, -18, -66, 57, 13, -128, -128, 8, 47, 39, 109, 127, 127, -74, -128, -128, 116, -3, -128, 15, 127, 127, -28, -112, -128, -128, 7, 127, 127, -26, -78, 107, 127, -1, -128, -128, -121, -28, -37, 1, 114, 127, 127, 127, 116, 32, -128, 6, 127, 127, -113, -128, -80, 111, -69, -128, -76, 58, 17, 54, 127, 123, 8, 10, 5, 12, -122, -102, -71, 97, 1, -32, 118, 127, -37, -2, -66, -58, -121, -68, -48, -13, -64, 114, 127, 101, -128, -128, -63, 33, 49, -128, -128, -128, -76, 8, 71, -24, -39, -6, 15, -128, -128, -96, 97, 127, 127, 71, -23, -22, 91, -5, -113, -128, 45, 18, -26, 127, 127, 127, 127, 106, -50, -128, -57, 127, 127, 127, 127, -28, -128, -17, 127, 127, 118, -32, -128, -128, -44, 38, 96, 15, 127, 76, 96, -64, -65, -68, -97, -128, 11, -68, -128, -128, -15, 49, -79, -128, -128, -3, 127, 127, -15, -28, 100, -10, -128, -128, -128, -81, -88, -66, -2, -88, -128, -57, -50, -8, -11, 127, 127, 127, 0, -49, 36, 8, -128, -128, -128, -81, 97, 127, 127, 33, 98, 127, 66, 2, -96, -128, -127, 87, 26, -103, -29, -71, -34, -69, -95, -101, 57, 3, -101, -128, 91, 127, 119, 58, -81, -128, -128, -128, -128, -100, -95, 0, 32, -100, -128, -128, -128, 39, 127, 102, -128, -128, -128, -106, 116, 127, -6, -16, -48, 59, -37, 53, -71, -81, -128, -107, -78, 17, 116, 63, -49, -43, -45, 127, 127, 127, 78, -128, -128, 55, 37, -128, -64, 15, -128, -32, 39, -3, -93, 127, 127, 127, 78, -28, -128, -128, -128, 53, 127, 127, 73, -128, -128, 2, 96, -128, -128, -128, -128, -123, 38, 103, 127, 122, 74, -124, -128, -36, -122, -128, -128, -128, -128, -128, 18, 23, -39, -78, -75, -128, -31, 118, 34, -128, -128, -15, -71, -79, 50, 48, 127, -66, -128, -128, -18, -45, -6, 34, 44, -39, 119, 102, -42, -128, 70, 127, 127, -112, -128, 32, 86, 6, 127, 127, 127, 48, 3, 79, 127, 22, -65, -128, -128, -73, -11, 54, 8, -92, -113, -44, 109, 27, -128, -128, -128, -128, 2, 3, -58, -128, -26, 68, 43, -68, -3, -16, -128, -95, -73, -128, -73, 65, 22, -52, -49, 127, 127, 13, -70, -16, -55, -66, -128, -74, 0, 63, 8, 38, 71, 78, -128, -128, -128, -21, 21, -44, 2, -15, 5, -70, 13, 118, 127, 127, 127, 93, 27, 70, 66, 73, -66, 48, -28, -79, -48, -85, -128, 52, 114, -128, -128, -109, 127, 127, 52, 118, 122, 36, -48, 50, -12, -76, 127, 127, 127, 86, -128, -121, 49, 10, -69, 65, -32, -103, 11, 42, 47, 127, 114, 22, 55, -97, -128, 3, 60, -91, -18, -91, 76, 59, 22, -128, -128, -76, -128, -87, 11, 127, 79, 38, -39, -22, 63, 123, 65, 127, 127, 88, -76, -128, 16, 127, 112, -31, 127, 127, 127, 59, 64, -3, -102, 28, 64, -21, 10, 27, -24, -78, 53, 127, 127, -128, -128, -123, -108, 5, 127, 127, -128, -128, -128, -74, 21, 127, 127, 127, 38, 95, 43, 127, 122, 127, 127, 117, 12, -53, 87, 127, 127, 21, -12, 10, 127, 122, 109, -37, -128, -66, 93, 127, 127, 0, -128, -121, 124, 18, -128, 86, 73, -103, -128, -57, -24, -128, 2, -11, 97, 91, 13, -128, -128, -128, -8, 97, -10, -128, -128, -128, -128, -128, -76, 69, 127, 127, -68, -45, -64, -128, -117, 27, 50, 81, -12, -128, -128, -128, -128, 31, 127, 127, 127, 36, 97, 15, -91, -21, 127, 127, 118, 107, 98, 16, -32, 127, 127, -26, 12, 127, 15, 13, 81, 39, -87, 45, -10, -128, -128, -88, -79, -50, -128, -26, 127, 127, 11, -128, -128, -81, -88, -36, -122, -128, -97, -21, 17, -57, -119, -79, 60, 37, -128, -128, -47, -128, 1, 127, 127, 55, 93, 42, 47, 74, 42, 70, 47, 3, 124, 127, 6, -128, -128, -42, 26, 127, 127, 69, -128, -128, 78, 15, -69, -128, -128, -128, -128, -111, -58, -114, -128, -128, -47, 127, 127, 7, -117, -128, -128, -128, -71, -39, -26, -108, 118, 127, 127, 92, -79, -128, -66, 8, -128, -128, -128, -78, 6, 15, -103, -36, 0, -17, -42, 70, 127, 127, 69, -95, 26, 37, -106, -68, 11, -128, -128, -108, 127, 27, -128, -128, -38, 127, 127, 47, 6, -34, -90, -96, 119, 127, 127, 127, 106, 18, 16, 88, 124, 17, 112, 127, 92, -107, -128, -81, -26, -117, -54, -128, -128, 50, 127, 127, -26, -73, -34, -128, -128, -128, 68, 124, 98, 127, 127, 75, -128, -128, -128, -64, -119, -128, -128, 53, 127, 118, -128, -128, -128, -57, -54, -128, -128, -58, 57, 127, 127, 52, -108, -128, 22, 22, -5, -102, 100, 127, 13, -86, -10, 127, 127, 36, 23, 121, 32, -45, -128, -128, 26, 127, 127, -128, -128, -32, 127, 24, -58, 64, 127, 3, -24, 98, 127, -128, -128, -128, -100, -31, 127, 127, 127, 127, 127, 127, -121, -128, -128, 38, 127, 127, -10, -128, -79, -12, -26, -128, -128, -108, -17, 6, -29, 81, 127, 106, 32, -42, -128, -95, -3, -106, -97, 103, 127, -75, -43, 59, 127, 127, -42, 34, 127, 127, -128, -128, -128, 8, 127, 127, 80, 12, -87, 15, 33, -63, -128, -64, -28, -128, 27, 127, 127, -93, -28, 127, 127, 127, 127, 127, 88, -109, -128, -128, -128, 127, 127, 102, 109, 127, 65, -76, -44, -116, -119, 113, 127, 127, 127, -17, -113, -116, -86, -112, 73, 127, 127, 88, -87, -128, -128, -128, -112, -128, -68, 100, 127, 127, 127, 127, 127, -13, -128, -128, 127, 127, 79, 0, -1, -64, -128, -128, -55, 22, 52, 43, 24, -128, -128, -21, -69, 7, 127, 70, -73, -29, 118, 127, -93, -128, -128, 127, 127, 127, 123, 69, -128, -128, -33, 5, -128, -128, -90, -44, -7, 33, 0, -15, -13, 63, 127, 127, 117, -119, -128, -128, -38, -128, -112, -44, 48, -88, -128, 17, -22, 0, -45, 37, 34, 60, -81, -128, -45, -59, -118, -128, -39, 123, 93, -11, 86, 96, 27, -75, 23, -2, -81, -27, 116, 127, 69, -85, 121, 127, 36, 13, 93, 6, 17, -128, -128, -128, -74, -29, 127, 127, 63, 0, -70, -128, -128, -65, 68, 127, -21, -128, -128, -128, -128, -100, -128, -128, -116, -60, -13, -17, -128, -128, 74, 127, 88, -128, -128, -88, -33, -122, -128, 38, 121, 87, -128, -128, -107, 127, 127, 86, -15, -44, -37, 66, -18, -34, -47, -128, -92, -81, -96, -90, -128, -128, -128, 48, 31, -18, -43, 39, 70, 127, 79, 127, 127, -55, -128, -128, -128, -1, -23, -90, 33, 127, 5, -128, -43, 8, 8, -128, -53, 103, 127, 127, 58, 127, 65, -128, -128, -86, 5, -11, -63, -26, -128, -34, -102, -21, 92, 127, 127, 127, 127, 80, -12, -13, 127, 127, -128, -128, -17, 127, -60, -128, -128, -128, -128, -108, -128, 42, 127, 100, -45, -58, -75, 43, 37, -107, -54, 127, 33, -70, -74, -85, -66, 49, 127, 127, -109, -22, 29, -12, -128, 21, 47, -57, -11, 127, 127, -16, -128, -97, 127, -2, -128, -128, -128, -59, 127, 127, -64, -128, -128, 88, 127, 127, 45, -121, -112, -32, -117, -28, 127, -48, -128, -12, 17, -91, 31, 13, -5, -128, -113, -6, 127, 127, -18, 3, 90, -32, -128, -116, -73, -102, 8, 127, 127, 127, -12, -122, -32, 123, 124, 8, 48, 127, 127, 127, -47, -128, -128, -128, -128, -88, 127, 127, 111, -128, -128, -112, -42, -54, 103, 87, 6, -73, -49, -128, -128, -71, 95, -22, -128, 32, 127, 10, -7, 127, 127, 127, 34, -100, -128, -68, 36, 102, -122, -128, 127, 127, 127, -128, -69, 106, 124, 49, -34, -128, -29, 119, 65, -113, -58, 127, 127, 12, 69, 127, 6, -108, 48, 80, -42, -80, -24, -117, -128, -128, 52, 108, 127, 127, 127, 66, 76, -63, -128, -128, -114, -91, -50, 44, 127, 31, -128, -128, -128, -128, -1, 98, 111, 127, -39, -128, -128, -26, -74, -119, -128, -58, 44, 60, 10, 3, -86, -128, -128, -101, -128, -128, 5, 127, 127, 76, -91, -39, 16, 27, 31, 31, -78, -29, -128, -97, -57, -28, -34, 76, 43, -128, -128, -73, 8, 43, -128, -128, -128, -71, 100, 127, 75, -28, 127, 127, 109, 127, 127, 116, 13, 127, 127, 123, -75, -7, 65, 101, -107, -38, -58, -52, -81, 74, 86, 127, -92, 10, 96, 127, -64, -73, 2, 45, -128, -128, -128, -76, -100, -117, 127, 85, 47, -95, -66, -73, -28, -123, -71, 127, 127, 127, 127, -127, -128, -128, -128, -28, -28, -128, -128, -43, -48, 103, 127, 68, -128, -128, 42, 127, 13, -128, -128, 52, -6, -39, -128, 119, 127, 22, -128, 112, 127, 127, -128, -128, 29, 127, 93, 24, 127, 127, -47, -36, 90, 127, 58, 76, -59, -128, -122, -106, -69, 127, 127, 127, 101, 22, 0, -12, -22, -71, -23, -128, 13, 5, -128, -128, -76, 22, 57, 18, -114, -8, 127, 55, -128, -128, 27, 65, -5, -74, -24, -128, 2, 127, 96, 15, -5, -128, -128, 64, 127, 0, 127, 127, 37, -128, -128, -48, 117, 39, -128, -11, 81, 127, 127, 127, -39, -128, -80, 127, 10, -128, -7, 117, -71, -128, -128, 28, 127, 107, -93, -6, 127, 127, 10, -128, -124, 59, 16, -128, -128, -128, -118, -93, -31, 36, 22, 11, -128, -128, -128, -128, -73, -13, 65, 71, -29, -128, -87, -3, -23, 127, 127, -127, -128, 64, 127, 31, -57, -76, -128, -128, 45, 127, 127, 127, 127, 127, 127, 127, -103, -128, -128, -54, 71, 60, 44, 127, 118, -75, -66, 127, 127, 47, -80, -128, -15, 31, 11, -49, 37, -52, -128, -128, 76, 127, 107, -128, -22, 127, -33, -117, -43, -39, -128, -64, 102, 127, 22, -128, -69, 127, 114, -128, -39, -34, -128, -128, -128, -128, 29, 127, 127, 109, -121, -128, -53, 127, -2, -128, -95, 127, 127, 100, -29, 53, 119, -128, -109, 69, 90, -128, -116, 108, 47, -128, -45, 127, 127, 106, 127, -108, -128, -128, 18, 127, 127, 127, 65, 80, 127, 127, -64, -128, -128, -5, -108, 48, 127, 127, -128, -128, 32, 127, 127, -18, -128, -91, 127, 127, 127, 127, 127, 127, 52, 127, 127, 103, -128, -100, 127, 127, 127, -102, -128, 28, 127, 127, 39, 49, -18, -128, -128, -24, -12, -42, 87, 93, 42, 76, 127, 26, 0, -24, 95, 101, 54, 23, 37, 54, 37, -128, -128, -98, -98, 69, 111, 21, -128, -128, -27, 34, -127, -128, -38, -128, -128, -32, 127, 5, -128, -119, 127, 127, -10, -93, 54, 127, 127, 127, -93, -128, -8, 66, -128, -128, -128, -107, -95, 81, 127, 127, 127, -5, -70, 79, 127, 127, -79, -128, -128, -44, -5, -128, -128, -128, 2, 127, -6, -128, -128, 27, 121, 92, 33, 127, 127, 91, -68, 45, 37, -18, -85, -64, -128, 34, 74, -37, -128, -128, 88, 26, -88, 68, 127, 96, 12, -52, 18, 55, 127, 12, -128, -128, -117, 93, -33, -128, -36, 33, 50, 101, -48, -128, 81, 127, 127, -128, -128, -128, 70, 36, 16, -17, -128, -128, 127, 127, 127, -5, -53, 11, -55, -70, -128, -55, -128, 33, 127, 127, 127, 96, 127, 79, -18, -12, 92, 54, 55, -73, -128, -128, 127, 111, -118, 33, 127, 127, -128, -128, 100, 124, -106, -128, -128, -128, 28, 3, -128, -128, -17, 86, 60, 127, 127, 127, 127, 127, 36, -32, -127, 29, 119, 127, 127, 127, 114, 122, 106, 1, -38, -1, 2, 79, -59, 7, -101, -128, -106, 127, 127, -32, -128, -65, 76, -43, -34, 21, 10, 127, 60, -128, 13, 127, -34, -128, -113, -39, 37, 127, 127, -128, -128, -128, -118, -107, -117, -16, -128, -113, 33, 127, -22, -128, -86, 28, 26, -124, -44, -16, -6, -63, 13, 37, -128, -76, -95, 127, 127, 39, -55, 3, 127, 79, 81, -50, -128, -128, -128, 13, 127, 80, -59, 49, 127, 74, -128, -128, -128, 108, 127, 127, -73, -76, 96, 49, -47, -128, 11, 127, 127, 127, 127, 26, -128, -128, 27, 36, -128, -128, -13, 65, 127, 127, 37, -128, -101, 59, -109, -116, -6, 29, -109, -128, -128, -63, 53, 58, -128, -128, -128, -128, -128, -128, -128, 85, 127, 127, -65, -6, -47, 127, 103, 127, -28, -48, -128, -23, 36, 38, -123, -128, 1, 127, 127, 97, -57, -38, 32, 124, 50, 127, 127, -128, -128, -128, -33, 74, 127, 90, -50, -103, -128, 107, 127, 127, -2, -100, -121, -49, -11, -86, 86, -74, -64, -63, 127, 23, -128, -128, -27, 127, 127, 90, -27, -128, -112, 127, -2, -128, -128, -128, -128, -128, 108, 127, 127, -95, -128, -128, -18, 21, 127, -45, -128, -128, -85, 127, 127, 3, -116, -71, -76, -39, 127, 127, 127, 127, 93, 43, 113, 91, -69, -128, 26, 49, -66, -2, 127, 127, 64, 78, 76, -78, -58, 47, 102, 38, 79, -128, -128, -128, -128, 74, 127, 127, 114, 127, 127, 127, 127, 60, 85, 68, 127, 127, 71, -128, -47, 127, 39, -128, -128, -81, -117, -128, -80, 24, 127, 33, -128, -128, -128, -49, 127, 127, 127, 10, -128, -128, 43, 112, -128, -128, 8, 127, 21, -128, -53, 127, -1, -98, 58, 71, -66, -128, -128, -102, -58, 11, 98, 6, -128, -52, -66, -70, -24, 127, 44, -128, -86, 127, 127, -80, -128, -74, 32, -102, -91, 29, 71, -78, -128, -128, -128, -95, 102, 127, 106, -128, -86, 127, 85, -68, 96, 50, -123, -128, 80, 127, -43, -128, -16, 127, 127, -28, -5, 127, -7, -11, -53, 29, -91, 95, 39, 6, 27, 127, -12, -114, -128, -44, 28, 70, -91, -97, 127, 127, -50, -128, -128, 127, 127, -122, -128, -128, -66, -88, -24, 127, 118, 11, -128, -128, -49, 92, 59, -119, -128, 88, 50, -42, -128, -128, -128, -52, 21, 127, 127, 127, -69, -128, -128, -128, -8, -50, -128, -128, 8, 127, 127, 69, -92, -128, -128, 33, 127, 97, 91, 127, 127, -128, -128, -10, 71, 38, -128, -128, -128, -98, -128, -128, 57, 127, 127, -57, -128, 65, 127, 127, 92, 108, -50, -13, 127, 127, 92, -128, -128, -128, -86, -109, -92, -18, 79, 101, 87, -128, -59, 26, 37, -116, 70, 127, 127, 23, -98, -128, -128, -128, -128, -128, -60, 113, 127, 127, 50, -27, 43, 69, 101, 127, 127, -128, -39, 127, 127, -44, -63, -76, 42, 127, 127, 127, 48, -79, -128, -128, -2, 36, 111, 127, -31, -128, -102, 109, 127, 39, -101, -128, -128, -128, 3, 127, 127, -75, -128, -128, -128, 0, 93, 100, 59, 66, -97, -128, -109, 88, 80, 100, 127, -127, -128, 52, 127, -68, -128, -95, 117, 34, -16, -21, -38, 17, 103, 112, 127, 101, -121, -11, 127, 127, 127, -109, -128, -18, 90, -21, -13, 127, 127, -123, -128, -124, 93, 79, 21, 113, 127, 127, 45, 107, -116, -128, -128, 127, 127, 15, -128, -122, 127, 108, -2, -11, 86, -74, -28, -127, -128, -96, 59, 92, -128, -128, -128, -18, -128, -128, -28, 127, 127, -100, -128, -66, 3, -96, 3, 43, 48, 22, -26, -128, -15, 127, 127, -128, -128, 3, 127, 65, 119, 68, 70, 17, 127, 103, 107, 13, -81, -10, 101, -8, -18, -43, -128, -106, -128, -128, -128, -128, -68, 96, -5, -128, -47, 44, 78, 111, -100, -128, -128, 23, 54, 127, 127, 28, 22, -101, -128, -128, 127, 127, 127, -3, -16, -44, -65, 103, 127, 127, -116, -128, -43, -52, -128, -128, -128, 68, 127, 122, 32, -43, -26, 22, 127, 127, 73, -117, -128, -91, -128, -128, 49, 127, 39, 23, -65, 6, -50, 116, 127, 127, 127, -44, 15, 68, 10, -29, -6, -128, -128, 127, 127, 127, 76, -17, -103, -128, -128, -118, 127, 127, 59, -92, -128, -128, -69, -33, -128, -128, -128, -7, 65, 127, 127, 127, -112, -128, -80, -81, -122, -128, -58, 127, 127, 26, -57, -23, 117, 127, 66, -128, -128, 127, 127, 127, -10, -117, -86, 127, 127, 102, -128, -128, -128, -128, -80, -15, 68, 127, 79, -91, 0, 127, 127, 93, 127, 127, 68, -15, -1, 10, 15, 127, 127, -58, -128, -128, -128, 32, 127, 18, -128, -128, -128, 124, 28, -128, -108, 127, -27, -116, -27, 66, -128, -128, -92, -1, -65, -76, 1, 127, 34, -128, -128, -107, 87, 95, -60, -102, -128, 74, 127, 39, -8, 127, 127, 55, 71, 127, 127, -48, 55, 127, 0, -128, -128, -64, -79, -113, -34, 127, 127, -29, -128, -50, 111, 127, 127, -5, -128, -128, 50, 127, 118, 42, -53, -45, 24, 69, 127, 127, -28, 42, 127, 127, -128, -128, -128, 0, 27, 53, 28, 127, 106, -55, -59, 5, -27, -102, 79, 122, 31, -71, 55, 111, 12, 87, 79, -52, -128, -128, -108, 127, 127, 127, 127, -33, -118, -13, -69, 24, 2, 106, -10, 47, 111, 127, 3, 101, 119, 98, 127, 34, -1, 127, 127, 127, 53, -121, -128, -27, 111, 127, 127, 107, -52, -128, -128, -17, 33, 97, 127, 127, -12, -6, 49, 116, 102, 93, 87, 59, 127, -54, -128, -128, 29, 24, 31, -17, 36, -15, -127, 16, -80, -119, -92, -65, -116, 127, 127, 29, -128, -128, -38, 48, 127, 127, 113, 43, 8, 52, -65, 96, 127, 112, -128, -128, -128, -53, 75, 33, 121, 127, 127, 13, -128, -106, -1, -79, -111, 13, 127, 127, 18, -75, -69, 32, 38, -121, -128, -128, 63, 127, 127, -128, -128, -128, -29, 31, 0, -128, -98, -69, 127, 64, 15, 3, 127, 97, 28, -37, 13, -76, -70, 127, 123, 92, 121, 127, 100, 127, 95, 59, 127, 127, 127, 48, -15, -32, -65, -98, 123, 127, 50, -128, -128, -24, -68, -123, -103, 79, 127, 127, 127, 48, -128, -102, 3, -65, -58, 127, 68, -59, 3, 23, -128, -128, -108, -128, -128, -128, 43, 17, 22, 27, 127, 10, 63, 113, 127, 127, 87, -70, -91, -85, -92, -128, -116, 127, 127, 87, -128, -107, 6, 127, 127, 127, 127, 127, 102, -42, -128, -128, -117, -28, 59, 8, -128, -128, -128, 102, 127, 127, 69, -34, -128, -48, 127, 2, -128, -128, 127, 107, -109, -57, 127, 127, -27, -128, -39, 127, 73, -71, 10, 75, -57, -128, -128, -128, 21, 117, 95, 27, -74, -128, -128, 43, 127, 127, -108, -128, -49, 127, 127, 47, 26, -10, -128, -69, 33, 127, 127, 2, -128, -128, -128, -91, -128, -91, -45, 38, 13, -102, 87, 16, -128, -128, -128, 8, 127, -1, -128, -116, 127, 127, 43, -28, -103, -128, -128, 103, 49, -58, -13, 5, 63, 127, 127, -54, 33, -16, -127, -128, -124, -6, 123, 5, 5, 21, -12, -6, 127, 2, 7, 38, 127, 27, -80, -128, -128, -128, -5, 127, 127, 2, -69, 102, 127, 127, 127, -10, -128, -128, -85, -66, -128, -128, -128, -118, -64, -3, -48, -128, -31, 127, 32, -128, -93, 127, 127, 122, -3, -28, 127, 127, 28, -66, 49, 60, -44, 69, 127, -34, -106, 57, 85, -53, -102, -128, -90, 127, 127, 127, -106, -128, -128, -128, -128, 43, 57, -71, -117, -74, 127, 127, -58, -128, -48, 127, 127, -111, -96, 74, 114, 42, -37, 101, 127, 127, -88, -26, 123, 127, 18, -22, 31, -38, -80, -128, -47, -10, -57, -80, 98, 122, 55, 23, 50, 34, -44, 0, 127, 127, 127, 112, -128, -47, 127, 127, -78, -113, -17, 127, 76, -107, -31, 127, 33, -117, -100, -44, -128, -127, 127, 127, -26, -29, 112, 127, -128, -128, -128, -128, -128, -109, 121, 127, 90, -8, 6, -66, 31, -12, 91, 12, -128, -128, 33, -74, -128, 76, 127, 102, 97, 127, -16, -18, 65, -11, -128, -128, 127, 127, 127, 127, -128, -128, -11, 22, -6, 106, 127, 81, 23, 11, 127, 127, 127, -44, -128, -128, -60, -128, -8, 127, 63, -128, -128, 59, 92, 31, -109, -13, 50, 127, 127, 10, -81, 33, 59, 116, 127, 127, -12, -123, -50, 43, 127, 2, 65, -91, 111, 127, 127, 15, -123, -128, -60, 127, 127, 111, -80, -128, -42, 127, 127, -33, -128, -128, -54, -111, -128, 79, 127, 127, -128, -75, 127, 93, -128, -128, -128, 119, 109, 29, 37, 102, -78, 7, 5, 59, -42, 70, 33, 16, 58, -95, -86, 76, 54, -128, 0, 127, 52, -68, -26, -128, -128, -128, 63, 26, -121, -117, -128, -128, -128, 127, 127, 127, -11, 13, 36, -113, -128, -128, 98, 122, 85, 43, -53, -128, -111, -121, 28, 127, 127, 10, -57, -92, -128, -32, 127, 123, 38, 80, 127, 127, 127, 127, 127, 127, 27, 3, 127, 121, -128, -128, -88, -128, -44, 127, 127, 76, -128, -128, 127, 127, 23, -69, -128, -128, -96, -75, 55, 38, 16, -128, -31, 55, 15, -118, 44, 44, 116, 78, 127, 52, -69, -128, -128, -109, -102, 0, 66, 127, 33, -2, 127, 127, 43, -128, -128, -17, 97, 127, 127, -53, -58, 79, 68, -128, -128, 96, 127, 63, -80, 68, 127, 73, -117, -128, -128, -74, 127, 127, 127, -95, -128, -128, 42, 127, 11, -128, 47, 127, 59, 21, 127, 127, -102, -111, -43, -122, -128, -95, 95, 127, 127, -3, -33, 49, 127, 127, -92, -128, -128, -128, 5, 127, 127, 127, 101, 60, 85, 29, -44, 68, 54, 74, 127, 127, -42, -87, 63, 127, -92, -5, 54, 127, 127, 127, 47, -6, -128, -128, 95, 112, -16, -54, 127, 127, 127, 127, 70, 12, 70, 29, 26, -28, 8, 37, 127, 127, -96, -128, -128, -39, -45, 33, 127, -117, -128, -16, 127, 127, 124, 22, -128, -128, 23, 127, 127, 86, 127, 87, 31, -111, -6, 90, -7, -128, 63, 127, 127, -96, -128, -10, 91, -44, -128, -128, -128, -13, -5, -128, -128, 38, -98, -123, 123, 127, -73, -128, -128, 34, 123, -38, -103, 91, 127, -8, -128, -128, -128, 27, 127, 96, 71, 12, 58, -27, 42, -93, 76, 127, 107, -128, -108, 18, -27, -64, -80, 59, -86, -128, -128, 31, 96, -57, -128, 96, 127, 127, -6, 58, 106, 76, -128, -128, -128, 44, -53, -85, 53, 12, -128, -52, -43, -109, -128, -44, -11, -93, -128, -74, 127, 127, 81, -3, 10, -12, -128, -100, -128, -128, 45, 127, 127, -23, -76, -87, -74, 53, 22, -60, 16, 8, 15, 127, 114, 116, -63, -128, -128, -49, 85, 68, 6, 28, -71, 112, 69, -128, -128, -57, 127, 127, 0, -128, -128, 68, 127, 127, -36, -90, -107, -39, -78, 127, 127, 127, -103, -128, -92, 33, 127, -108, -128, -128, -23, 127, 127, 127, -18, -128, -111, -75, -128, -128, -128, -43, 26, -116, -128, -128, -43, 44, 127, 127, 80, 12, -22, -58, -101, 127, 127, 57, -128, -93, 122, 127, 127, 28, -128, -128, -91, 127, 127, -112, -128, -128, -78, 111, 69, -54, -128, 108, 109, 127, -42, 91, 7, -102, -28, 127, 118, -58, -128, -128, -48, 100, 114, 127, 127, -37, -38, -17, 43, -48, 127, 24, 127, 6, 13, -2, 127, 55, -128, -96, 31, 15, -128, -128, 74, 127, 64, -128, -128, -64, 108, 127, 127, 127, 127, 127, 102, -85, -117, 74, 47, -102, 5, 127, 76, -124, -128, -128, -52, -116, 23, 59, -128, -116, 90, -36, -128, 127, 127, 68, -128, -128, -128, -128, -128, -103, 127, 127, 17, -128, -128, -42, 60, -39, -128, -128, -128, -73, -21, 127, 75, -34, -128, -26, 127, 127, 127, 23, 36, 24, -128, -128, -111, -49, 73, 113, 118, 28, 127, 127, 127, -80, -128, -128, -15, 58, 78, -85, -10, 78, 127, 102, -23, -109, -128, -128, 5, 127, 22, -128, -128, 127, 127, -109, -18, 127, 127, 127, 127, 127, -64, -128, -85, 86, 29, -74, -34, -54, -1, -114, -97, -12, 90, 127, 28, -128, -128, 44, 45, -66, -98, 58, 127, 127, 114, -128, -128, -68, -128, 21, 50, -39, -16, 106, 52, -68, 127, 127, 11, -49, 34, 49, 95, 123, 91, 79, 127, 127, 127, 127, -50, -128, -128, -91, -128, -128, -128, 103, 127, 127, 49, -128, -128, -117, -128, -123, 122, 28, -28, 68, 124, -128, -128, -36, 127, 127, 47, -78, -128, -121, 127, 127, 21, -128, -49, 127, 107, 127, 127, 127, 127, 91, 124, 116, 68, -23, 127, 127, 127, -108, -128, -27, 127, 44, -128, -128, -106, 53, 75, -6, -112, -122, -128, 1, 127, 21, -12, 23, 127, -87, -128, -128, -128, -128, 127, 127, 127, 36, -60, -52, 121, 127, 127, -26, -33, -22, -128, -128, -90, -102, -128, -128, -22, -16, -90, -119, -69, -128, -80, -32, 127, 127, 76, -128, -128, -128, -128, 18, 127, 27, -128, -128, 117, 76, 42, -31, -54, -128, -42, 127, 58, -128, -128, -101, 52, 122, 122, 66, 49, -128, -128, 10, 101, 6, -128, -128, -128, -128, -128, -55, -103, -128, -128, -68, -39, -92, -68, -98, -121, 87, 44, -128, -128, 81, 127, -69, -128, -128, 31, 127, 127, 127, 29, -128, -128, -32, 85, 48, -91, -98, 114, 27, -128, -107, 127, 63, 13, 127, 127, 127, 50, -128, -128, -53, 127, 127, 127, 109, 32, 69, 127, 127, 64, -26, -128, -86, 127, 127, 23, -128, -128, 98, 127, 127, 127, 0, -128, -128, -128, -128, 10, 127, 127, -108, -85, -128, -128, -32, 100, 54, -73, 8, 8, 73, -100, -128, -3, -6, -79, -128, -118, -52, -66, 38, 34, -128, -128, 127, 127, 127, 59, -44, -43, -10, -12, -18, 49, -54, -128, -128, 34, 93, 28, 5, 106, -13, -57, -128, -38, -31, -128, -128, 0, 95, -108, -128, -68, -57, -54, 10, 10, -108, -92, 127, 80, -103, -1, 127, 127, 8, -27, 80, 127, 58, 49, 113, 127, 49, -128, -128, -128, -5, 127, 127, 85, -85, -128, -128, 127, 127, 103, -43, 11, 127, 127, -118, -128, -86, 33, -6, 31, 127, 127, 65, 15, -58, -128, -128, -128, -128, 11, 127, 127, -69, -86, -48, 27, -47, 69, 21, 66, 18, -75, -128, -64, 54, -8, -92, -128, 33, 69, 59, 85, 90, 36, 124, 127, 2, 54, 127, 127, 44, 127, 127, -6, 45, 127, 54, -128, -128, 70, 127, 127, -47, -128, -13, 101, -128, -128, -111, 64, 27, -38, 122, 22, -128, -128, -112, 31, 127, 103, 127, 127, 103, -116, -27, 127, 91, 96, -8, 32, 37, -128, -128, -11, 127, 127, 127, 117, -33, -113, -74, -38, -78, 42, 121, 127, -24, -128, -128, -128, -128, 36, 127, 127, -38, -128, -128, -42, 79, 127, 127, 74, -5, 97, 127, 47, -116, 100, 127, -33, -128, -2, 53, 86, 22, -128, -128, -69, -17, -109, -28, 117, 127, 78, 127, 127, 127, 127, -57, -37, 127, 127, 122, 118, -96, -128, -7, 127, -1, -128, -128, -128, -121, 81, 127, 17, -106, 101, 127, 127, 127, 68, -68, -128, -128, -128, -128, -128, 45, 91, 76, -29, -117, -128, -128, -128, -128, 5, 102, 112, -116, -128, -60, 127, 127, 78, 24, 90, 50, 47, -1, 26, 127, 127, 127, -128, -128, -48, 52, -39, -111, 118, 76, -17, 127, 127, 127, -32, -128, 42, 109, 2, -49, 1, -16, 127, 127, -79, -49, 28, 97, 54, -85, -92, -15, 127, 127, 127, 127, 127, -98, -128, -33, 127, 127, 127, 127, 28, -100, -57, -15, -81, -128, -16, 119, 127, -24, -28, 109, -55, -128, -2, 127, 127, 34, -26, 10, -38, 106, 119, 127, 113, 127, -50, -101, 122, 127, 43, -88, -80, -128, -128, -128, -103, -128, -123, 117, 127, -7, -128, -128, 127, 127, 113, 70, 117, 107, 112, -79, -128, -65, 123, 96, -3, 124, 127, -128, -128, -70, 127, 127, 127, -107, -128, -128, 118, 127, 86, -32, -117, -128, -128, -75, -128, -128, -128, -33, -11, 55, 63, 80, 28, 112, -44, -123, -128, 59, 127, 127, -86, -8, 127, 127, -116, -128, -128, 127, 127, -43, -13, 0, -95, -128, -70, 69, -8, -64, -128, -128, -128, 119, 118, 70, -3, -128, -128, -128, -18, -59, -1, 127, 117, -32, -124, -113, -128, 127, 127, 127, 42, -33, -128, -123, -31, 36, -100, -128, -128, -93, -128, -34, -117, 27, 100, 80, -74, 33, 127, 24, 90, 98, -118, -114, 76, 127, 127, 7, -55, -74, -128, -103, 5, 127, 31, -128, -128, -128, 22, 8, 12, 112, 127, 5, -101, -128, -128, -57, 0, -128, -7, 29, -3, -128, -128, -128, -128, -119, 98, 65, -128, -128, 71, 106, -68, 45, -39, -38, -111, -38, -29, -128, 70, 58, 23, 15, 127, 127, 114, -128, -128, -128, 127, 106, -127, -128, -123, 81, 127, 127, -128, -128, -106, 85, 36, -128, -128, -39, -128, -128, -33, -90, -128, -128, -128, -128, -10, 127, 54, -128, -128, 127, 95, 43, -50, 111, 127, 127, 127, 127, 121, -47, -12, 47, 17, -43, 70, 92, -128, -128, -128, 37, 127, 55, -68, -128, -128, -128, -78, 127, 127, 127, -73, 15, 80, 32, -8, -58, -128, -10, 127, 80, -107, -43, 50, 127, 118, 11, 121, 127, 50, 23, 97, 127, 127, -100, -128, 69, 127, 127, -75, -128, -128, -58, -74, -128, -128, -128, -12, -32, 73, 127, 127, 127, 127, 127, 108, -127, -128, -128, 127, 127, 85, -15, 78, 80, -128, -128, -50, 75, 49, -128, -128, -5, 127, 127, 8, -128, -128, -128, -76, 0, -50, -69, 114, 127, -128, -128, -128, -23, -5, -109, -43, 127, 127, 5, -101, -97, 96, 103, 127, 127, 127, 65, 127, 127, -93, -128, -48, 127, 127, 43, -128, -128, -128, -128, 0, 127, 127, 127, 26, 109, 127, -75, -128, -128, 88, 64, -71, -113, -100, 123, 39, -7, 53, 68, -121, -15, 127, 127, 15, -106, -128, -29, 73, -54, -128, -48, 63, -106, -128, -128, -128, -68, -128, -128, -121, 85, 127, 81, -78, -73, -64, -52, 39, 60, 117, 32, -128, -47, 127, 127, 92, 8, -128, -128, -128, -128, -118, -52, 69, 127, 127, 127, 127, 119, 44, 39, 10, 17, 55, 37, -101, -13, 127, 37, -128, -80, 127, 117, -74, -128, -76, -117, 71, 127, 127, 127, -71, -128, -128, -128, 127, 127, 127, -87, -128, -58, -128, -128, -128, -23, 68, -64, -128, -5, 127, 127, 18, -54, -17, 64, 16, -88, -128, -128, 58, 127, 127, -114, -128, -128, 38, 127, 127, 1, -119, 29, 111, -7, 18, 100, -92, -79, -114, 121, 95, 124, 98, 33, -128, -28, 2, -128, -128, 73, 90, 127, 113, 127, -95, -128, -128, 91, 127, -27, -37, -117, 16, 36, 127, 109, 26, -78, -128, -128, -22, 7, 119, 127, -128, -128, 17, 127, 113, 113, 69, -52, -128, -128, -128, -128, 44, 92, -11, 15, -12, -123, -108, 122, 127, 58, 127, 127, 127, 127, -29, -128, -128, -128, -71, -70, -118, -43, 42, 117, 118, 81, 127, -78, -119, 31, 127, 106, 95, 76, -103, -15, 127, 88, 50, 127, 78, -128, -128, -22, 13, -128, -43, 127, 31, -29, -13, -128, -47, 127, 52, 38, 127, 127, -12, -12, 48, 97, -103, -36, 111, 127, 117, -81, -38, 127, 122, -128, -128, -54, 119, 52, -128, -128, -128, -128, -128, -128, -128, 48, 127, 127, -128, -128, 34, 127, 127, -27, 17, -86, -54, -43, 127, 42, -48, 7, 111, 66, 65, -116, -128, -128, -112, 127, 127, 73, -128, -107, 96, 36, -10, 127, 127, 31, 127, 127, 106, 127, 127, -32, -128, -128, -73, 127, 127, 69, 0, 127, 118, 13, 16, 127, 127, 127, 127, 36, -5, 22, 45, -27, -42, -127, 18, -124, -113, -128, -114, -75, 127, 127, 11, -128, -128, -128, -13, 127, 127, -48, -128, -128, -24, -17, 127, 127, -23, -128, -96, -49, 21, -55, -128, -117, 48, 127, 8, -128, -39, 49, 49, 36, 0, 85, 127, 38, -128, -45, 127, 66, -128, -27, 127, -39, -47, 127, 127, -116, -128, -17, 127, 127, 108, 27, 12, 87, 127, 127, 127, 127, 68, 5, 42, 116, 88, -68, -127, -113, -43, -32, -43, -13, 123, 127, 53, 86, 127, 127, 93, 111, 28, -73, -70, 32, -3, 39, 127, -53, -128, -122, 0, -26, -43, -57, -128, -128, -65, 42, 127, 87, -17, 95, 118, -128, -113, 127, 127, 127, 0, -85, 43, 127, 127, 55, -31, -91, 1, 127, 127, 127, 53, 68, 18, -15, 17, -52, -128, -128, 23, 127, 127, 96, -98, -128, 16, 127, 127, -117, -128, -38, 118, 102, 6, -50, 64, 127, 127, -6, -128, -128, 29, -7, 44, -87, -128, -128, 69, 127, 127, -80, -128, -128, 70, 127, 76, -31, 127, 127, -2, 13, -59, -69, -70, 57, 28, 45, 98, 127, 127, 127, 18, -45, -128, -128, -16, 6, -128, -128, 52, 48, -47, -34, 127, 127, 26, -31, -11, 7, -15, -128, -128, -128, -32, -63, 1, 127, 127, 102, 85, 113, 17, 113, -28, -128, -128, 127, 127, 92, 34, 15, 127, 127, -15, -128, -128, -124, -32, 127, 16, -102, -80, 16, -128, -128, -53, 127, 127, 26, -95, -128, -128, -55, -31, -63, -128, -78, 36, -127, -128, -85, 54, -54, -128, -128, -128, -128, -128, -97, -11, 26, 70, 127, -26, -113, 1, -102, -128, -128, 37, -43, -128, -48, 127, 127, -109, -128, -128, 12, 27, 127, 127, 127, 127, -28, -128, -128, 127, 127, 127, 127, 42, -81, -114, -60, -23, -128, -43, 127, 127, 47, -47, -128, -128, -103, -128, -128, -5, 127, 127, 127, 127, -128, -128, -103, 32, -112, -128, -43, 124, 127, 5, -38, 98, 127, 127, -70, -96, 33, 55, 6, 85, 81, -78, -55, 106, 127, 127, 38, -128, -128, -8, 49, -27, -113, 44, 0, 21, -24, 34, 54, 79, 13, 127, 127, 127, 74, -112, -78, -21, 71, 127, 127, 127, 58, 95, 122, -54, -128, -128, 55, 71, -60, -42, 117, 127, 78, 1, -22, -42, -112, -32, -3, 48, 106, 47, 12, -128, -128, -80, -124, -76, 50, -86, -18, 127, 80, -10, 127, 127, 127, 95, 2, -66, 1, -54, -106, -128, -128, -81, 127, 127, 78, -70, -128, -128, -128, 43, -64, -128, 55, 127, 127, 65, 33, -128, -121, -55, -8, 5, 43, -128, -128, -36, -48, -128, -70, 127, 127, 24, 12, 2, -1, -128, -128, -128, 68, 127, 127, 97, -5, -69, -71, 76, 36, 11, 16, -70, 21, 49, -85, -78, -48, -69, -128, 48, 127, 109, -128, -128, -34, 23, 127, 127, -78, -128, -128, 71, 127, 85, -16, 45, 64, -1, 114, 45, 96, -79, -128, -100, 88, -34, -128, -87, 34, -107, -128, -128, -112, -128, -128, 38, 127, 33, -128, -98, 75, -13, -69, 13, 107, -66, -60, -128, -81, -71, 127, 127, 127, 127, 127, 16, -28, 63, 1, -128, -128, -117, -54, 53, 127, 127, 127, 10, 85, 85, -91, -128, -75, 127, 127, -48, -80, -116, 2, 101, 127, -65, -128, -79, 107, 127, 127, 64, -123, -128, -90, -8, -42, -36, -128, -86, -53, 57, 107, -70, -128, -128, 10, 127, 127, 49, 71, 95, 71, -128, -103, 119, 127, -21, -76, -128, 57, 127, 127, -11, -128, -47, -60, -50, 1, 88, 13, -57, -18, -71, 106, -26, 8, 127, 127, -2, 127, 127, 1, -128, -103, 127, 127, 75, -16, -117, 17, -55, -91, -108, 127, 127, 127, 107, 26, -27, -88, -26, 127, 127, -97, -128, -128, 47, 17, -97, -11, -106, -128, -128, -48, -16, -64, 119, 127, 101, -128, -90, 45, 32, -43, 17, 11, 127, 127, 12, -128, -128, -128, 48, 127, 48, -128, -128, -80, -128, -123, 50, 127, 127, 127, 127, 48, -128, -128, 101, 92, -31, -50, 127, 90, -45, -128, -5, 127, 127, 127, 59, 127, 127, 127, 119, 64, 71, -10, -116, -59, 81, -87, -128, -128, 16, -12, 49, 127, 90, -5, 1, -47, 127, 127, 122, -31, -81, -81, -74, -58, -128, -123, 106, 127, 69, 127, 37, -22, -128, -128, 53, 127, 97, -102, -128, -128, -128, -100, -37, -2, 127, -17, -128, -128, -128, -128, -128, -128, -107, 113, 108, -128, -128, 127, 86, -128, -128, 127, 127, 127, 118, -78, -128, 58, 127, 81, -42, -24, -26, 31, 127, 93, -128, -128, 34, 127, 127, 73, -81, -12, 54, -128, -68, -128, -128, -128, 66, 127, 81, -74, -55, 10, -121, -96, 37, 127, 74, -128, -128, -47, 44, -108, -128, -95, 127, 127, -24, -128, -117, -44, -128, -128, 55, 7, -128, -128, 64, 127, -52, -128, -75, 127, 127, 64, 53, 54, -128, -128, -128, -128, -44, 18, -22, -38, 87, 58, -43, 45, 45, 103, 118, 29, -128, -128, -128, 127, 127, 127, -36, -128, -128, -38, -11, 26, 127, 127, 127, 127, 127, 54, -69, -54, -109, 66, 127, 127, -119, -128, -128, 127, 127, 36, -128, 7, 127, 127, 26, -128, -128, -75, 127, 10, -128, -128, -27, 42, 127, 63, -48, -128, 42, 127, 127, 57, 127, 127, 127, 27, -128, -128, -36, 127, 127, -8, -128, -128, -128, -91, 57, 92, -128, -128, -128, -71, 127, 127, 95, -128, 0, 127, 127, -38, -128, -128, 38, 127, 27, -31, -7, 6, -121, -44, 127, -3, -74, 66, 127, 127, 18, -95, 86, 127, 103, -27, 60, 59, 34, -85, -53, -59, 87, 127, 39, -101, -59, -128, 49, 127, 127, 107, 1, -74, -73, -93, 8, -5, 38, -128, -29, 127, 127, 7, -128, -118, 127, 127, 112, 118, 127, 127, 127, 127, 127, 37, -53, -42, 13, -32, -39, 124, 127, -86, -128, 27, 127, 16, -102, 21, 127, -36, -65, 116, -63, -128, -128, -75, -128, -106, -24, 6, -8, 88, 127, 65, 65, 127, 8, -128, 15, 127, 127, 123, -63, -112, 39, 75, 16, 107, 127, 2, -48, 69, 127, -49, -128, -71, 85, 92, 127, 59, -15, -128, -45, 127, -92, -128, -8, 100, -22, -42, 12, 119, 117, 127, 127, 127, -100, -128, -34, 127, 76, -128, -128, -66, -117, -128, -78, 93, 127, 122, 60, 68, 21, 16, -63, -15, -44, 17, 11, -29, -128, -128, 102, 127, -37, -128, -128, -79, -92, 29, 127, 127, 68, 12, 2, 16, 127, 127, 15, -128, -75, 127, 93, -128, -121, -106, -64, -80, -3, 2, 100, 37, -66, -128, -32, -23, -121, -90, -74, 45, 10, -128, -121, -90, -17, 54, 127, 127, 127, 127, 50, -128, -128, -128, -128, -128, -128, -128, -114, 90, 127, 127, 127, -17, -128, -128, -23, 127, 127, -128, -128, 16, 127, 127, -128, -103, 127, 127, 52, -10, -98, -85, -128, -33, 127, 127, 127, 127, 127, 18, -128, -21, 106, -98, -128, -128, 78, 127, 26, 43, 127, 127, -5, 85, 127, -128, -128, -29, 127, 127, -128, -128, 66, 88, -102, -128, -70, -107, -128, -50, -55, 12, 127, 127, -23, -79, 11, 38, -38, -128, -128, -37, 123, 103, -29, 34, 114, 106, -59, -44, -38, -33, -128, -42, -63, -10, -128, -128, -128, 127, 127, -42, -128, -80, -43, -103, -92, -93, -12, -6, 127, 78, 74, -28, 108, 91, 81, -108, -88, -18, 38, -116, -128, -50, 127, 111, -63, -123, -119, -128, -27, 127, 127, 127, -53, -128, -23, 127, 127, -57, -128, -73, 127, 69, -88, -33, 10, -87, 5, 127, 127, 124, -80, -128, -128, 93, 23, -128, -119, -53, 93, 65, -44, -128, -128, -128, -128, -47, 91, 127, 127, -15, -128, -128, -128, 21, 127, 0, -128, -128, 103, 127, 127, 68, -28, -90, -66, 54, 127, 32, -39, -127, 38, 127, 127, -78, -80, -43, -80, -123, -128, -128, 108, 127, 127, 127, 97, -128, -128, 7, 127, 127, 127, 127, 127, 106, 43, -106, -128, 0, 127, 127, 127, 127, 127, -3, -123, 32, 127, 127, 98, 127, 127, 127, 86, 57, 73, -39, -92, -128, -128, -128, -128, -85, -58, -42, 79, 127, 116, -98, 93, 127, 58, -7, 127, 127, 127, 101, -65, -128, -117, -17, 47, -54, 87, 127, 127, -12, 28, 78, -76, -128, -43, 127, -7, -128, -128, -78, 127, 127, 55, -114, -102, -23, 127, 122, 127, 127, 101, -128, -128, 127, 119, -109, -63, 127, 127, 127, 39, -128, -128, -36, 127, 127, -68, -55, -18, 28, 106, 29, -128, -34, 127, 127, 7, -3, 28, 57, -92, -128, -128, 112, 73, -128, -113, 65, 53, -8, -43, -128, -107, 119, 44, 36, 127, 31, 1, 103, -55, -128, -128, -128, 31, 53, -15, 91, 127, 127, 60, -52, -128, -128, -128, 50, 127, 17, -128, -128, -100, -10, -60, -128, -73, 127, 109, -78, -92, 6, 69, 127, 127, 127, 127, 127, -75, -128, -128, 7, 127, 127, 127, 63, -49, -88, 79, 127, 127, 26, -90, -93, 2, 68, -128, -128, 53, 127, -52, -128, -108, 47, -42, -108, 17, 28, -90, -15, 127, 127, -109, -128, -116, -38, -109, 127, 22, -113, -128, 91, 127, 127, 12, 75, 127, 101, 17, 10, -128, -128, -128, 64, 57, -53, -78, 127, 127, 127, 78, -18, 81, 127, 0, -128, -128, -18, -96, -128, -128, -12, -1, -128, -128, -128, -8, 65, 38, -64, 21, 106, 127, 127, 47, -118, -101, 57, 63, 0, -29, -128, -128, -42, 12, 1, -29, -18, 117, 127, 127, 15, 73, 121, 63, -128, -128, -128, 8, 79, 91, 127, 91, -8, 44, 76, 32, 121, 49, -103, 17, 127, 24, -128, -128, -57, 127, 127, 91, -128, -128, 50, 127, 114, -128, -128, 0, 116, 26, -128, 33, 85, 23, -127, 66, 127, 127, 122, 127, 127, 31, -12, -1, -86, -128, -128, 98, 127, -45, -128, -128, -11, -58, -17, 27, 107, 127, 127, 127, 28, 0, -107, -128, -128, -128, -3, 127, 127, 73, -66, -128, -128, 93, 49, 0, 98, 127, -18, 32, -24, -76, -128, 48, 127, 102, -128, -128, -128, -128, -128, -128, -113, 12, -1, -96, -63, -128, -128, -128, -128, -59, -66, 11, 93, 15, -128, -66, 127, -7, -128, -128, 52, 127, 97, 10, 21, 127, -121, -128, -128, 16, -73, -128, -128, -128, -128, -128, -98, -10, 34, -21, -76, 55, 127, 127, 90, -128, -128, 34, 127, 127, 127, 48, 45, -98, -128, -42, 85, 53, -128, -85, 102, 127, -71, -128, -116, -37, -128, -128, 8, 64, -128, -128, -123, -128, -113, -7, 106, -122, -128, 127, 92, -63, -124, 75, -27, 127, 127, 127, -13, 44, 127, 33, -43, -114, 0, 39, 36, 23, 50, -21, -128, 2, 17, 24, 98, 127, 127, -17, -74, 3, 127, -10, -128, -57, 127, 127, 127, -93, -128, -128, -47, -128, -10, 127, 117, 11, 23, -2, 3, 65, -2, -75, 17, 127, 63, -128, -50, 127, 127, 22, 44, -37, 68, 127, 127, 127, 123, -36, -109, 13, 127, 69, 127, 127, 127, 127, 1, -128, -109, 127, 127, 127, -128, -128, -90, 81, 8, 85, 112, 60, -128, -128, -96, -3, -44, 15, 127, 127, 22, -114, -128, -118, -128, -50, -100, 13, 127, 127, -113, -128, 2, 6, -128, -128, -69, 80, 127, 127, -76, -128, -128, -128, -128, 127, 127, 39, -128, -85, -21, -128, -87, 127, 127, 59, -66, -47, 50, 127, 127, -7, 31, -58, -128, -68, 127, 127, 127, 127, 127, 60, 127, 87, -36, -128, -128, -128, -87, 80, 54, -73, -128, -128, 37, 127, -48, -128, -114, -8, -70, -100, -128, 113, 127, 127, -55, -59, 127, 127, 124, -79, -42, 108, 127, 27, -128, -128, -58, 76, 127, 8, -90, 23, 127, 127, -75, -128, -124, 55, 127, 119, 28, -69, -80, 48, 127, 127, 57, 38, 127, 127, -21, -43, 112, 96, 13, 17, 127, 103, 114, -121, -128, -128, 0, 127, 127, 127, 76, -87, -128, -128, -65, 45, 24, -128, -23, 127, 127, -59, -128, -52, 68, -53, -128, 47, 127, 113, -128, -128, 42, 127, 127, -117, -128, -128, 71, 100, -2, -123, 49, 107, 47, 5, 32, 57, 16, -128, -128, -65, 127, 127, 127, 116, 68, -75, -128, -54, 109, 70, -116, -128, -128, 78, 127, -18, -128, -128, -8, 100, 127, 79, -128, -128, 127, 127, 127, -100, -21, 127, 127, 127, -103, -108, -26, 24, -81, -39, -128, -128, 44, 127, 29, -128, -128, -86, -128, -108, 127, 127, -36, -128, -91, 93, 75, 13, -26, 33, 127, 102, 74, -7, -22, -49, -128, -80, 2, -100, 24, 32, 15, -128, 33, 127, 106, -33, 39, 93, 127, 80, 52, -12, 127, 127, 60, 23, -73, -128, -128, -48, 63, -17, -100, -29, -128, -128, -101, -128, -128, -102, 11, -16, -5, 114, 122, -75, -76, 64, 74, -21, -55, -109, -60, 0, 127, 121, 88, -128, -128, -128, 7, 127, 127, 90, -10, 64, 127, 58, -128, -128, -128, -128, -23, 127, 127, 127, 49, -63, 28, 123, -109, -128, -128, -119, 17, 127, 127, 80, -8, -8, -128, -128, -128, -106, -128, -128, -50, 127, 127, 127, -42, 68, 127, 127, 91, 127, 33, -26, -128, -128, -116, 127, 127, 43, -128, -128, -128, -102, -22, -11, -33, 44, 44, -6, -66, 69, 66, -86, -86, 127, 127, 6, -128, -128, -123, -128, -128, -76, 121, 127, 68, 12, 127, 127, 97, 71, 100, 107, 68, -87, -92, 127, 127, 87, -122, 2, 127, 127, 48, -63, -128, 10, 85, -128, -128, -128, 69, 71, 34, -86, -108, -128, 32, 127, 127, 96, 127, 118, 57, -93, -128, -119, 27, -108, -128, -54, -69, 0, 117, -23, 12, 127, 118, -128, -53, -128, -128, -128, -53, 23, 32, 34, 5, -100, -128, -103, 127, 127, -57, -114, 3, 127, 127, 127, -48, -128, -128, 127, 127, 127, 0, -128, -128, -128, -39, 59, 76, -10, -71, -124, -59, -69, 71, 127, 98, 11, -65, -128, -128, -16, -63, -128, -95, 91, 122, 127, 108, 127, 53, 121, -60, -128, -128, 33, 127, 43, -128, -128, -28, 87, -50, -128, -128, 71, 127, 127, 127, 127, 63, 13, 92, 86, 122, -127, 24, 127, 127, -8, -44, -81, -128, -111, 87, 127, 127, 121, 127, 127, 96, -47, -7, -2, -26, -128, -45, -17, -69, -128, -91, -128, -7, 28, -18, 113, 127, -85, -128, -111, 11, -86, -128, -81, 107, 127, 17, -128, -121, -65, -128, -128, 37, 127, 127, 102, -111, -101, 127, 127, 123, 60, 127, 127, 127, 127, 118, -69, -128, -128, 36, 70, 3, 21, -2, -88, -68, 90, 17, -87, -27, 76, 69, 37, -34, 127, 127, 27, -71, -50, -79, -128, -128, -58, 42, 76, 12, -128, -128, -36, 12, 11, 127, 127, 5, 1, 112, 44, -128, -128, 38, 106, -6, -128, -33, 127, 127, 64, -91, -16, 50, 127, 57, -106, -128, -128, -128, -44, 127, 121, -128, -128, -48, 114, 102, 55, 111, 15, -100, -59, -75, -128, -96, -128, -108, -64, 13, 23, 60, -31, 34, 33, -88, -128, -128, -55, 71, 127, 127, 58, 23, -18, -128, -27, -22, -53, -113, -36, -22, 37, -59, 39, 127, 127, -12, 44, 102, 10, -128, -122, -79, -128, 0, 127, 44, 109, 127, 127, 127, 11, -128, -128, 0, 116, 13, -128, -128, 0, -63, -128, -128, -73, 85, 127, 127, -128, -128, -34, 75, -57, -128, -128, -1, 127, 127, 127, 127, 16, -28, -128, -90, 17, 81, -26, -71, -34, 21, 127, 127, 68, -23, 70, 88, -55, -1, 22, -45, 13, 26, -76, -128, -128, -119, -31, 123, 127, 127, 112, 59, 93, 127, -16, -128, -128, -128, -76, 127, 127, 29, -68, 48, 127, 48, -86, 74, 127, -8, -128, -128, 39, 103, 127, 37, -26, -47, -73, -128, -128, -45, 127, 127, -43, -128, -42, 127, 73, 91, -88, -128, -71, 127, 127, 127, 127, 86, -124, -128, -128, -69, -76, -128, -128, -5, 127, 52, 32, 127, 127, 11, -116, -128, 27, 100, 127, -13, -127, -113, 127, 58, -128, 23, 127, 127, 102, 28, -34, 127, 127, 127, 127, 88, -28, 68, 127, 92, 45, 5, 96, -39, -128, -121, 127, -32, -128, -128, -43, -3, -103, -128, -128, -128, -101, 64, 119, 70, 81, 127, 32, -128, 2, 127, 127, 21, 0, -107, -128, -108, -128, -52, 127, 127, 127, 16, -44, 124, 127, 118, 103, -76, -100, -39, 127, 127, 86, -128, -128, -12, 127, 127, 27, -128, -128, -17, 127, 69, -128, -128, -128, -128, -128, -128, 69, 127, 54, 86, 127, 127, 38, 70, 109, 127, 127, 127, 127, 28, -100, -71, 13, 26, 127, 80, -68, -71, -71, -128, 2, 127, 127, 111, -87, -128, -128, -8, 127, 92, -128, -34, 103, -73, -128, -24, 37, -31, -108, -128, -34, -59, -112, -108, 92, 121, -13, -128, -128, 0, 111, -113, -128, 5, 44, 52, 74, 114, -42, -92, -29, 80, 37, 53, 127, 127, 127, 95, 52, -71, -12, 23, 2, 50, 13, -79, -57, 38, 52, -3, -98, -128, 106, 127, 55, -128, -128, 44, 127, 15, -128, 29, 116, -22, -79, -90, 39, 127, 127, 127, 127, 103, -123, -128, -111, 55, 98, 127, 127, 114, 52, 86, 59, -93, -128, -128, -128, -73, 87, 127, 127, 127, 127, -63, -128, -128, -121, 127, 127, 127, -17, 79, 127, 49, -22, -91, 127, 68, -128, -128, 73, 127, 86, -128, -113, 127, 127, 127, -102, -49, -45, -128, -102, 29, -102, -128, -112, -128, -128, 8, 117, 127, 36, -18, 127, 127, 42, 95, 127, 127, 127, 54, -54, -108, -128, -81, 127, 127, 127, 127, 121, 85, 119, -1, -54, 52, 127, 85, -128, -128, 55, 29, 57, 127, 127, -44, -128, -128, 50, 127, 127, -128, -128, -111, -22, -128, -128, 65, -26, -31, 81, -34, -128, -18, 127, -97, -128, -70, 127, 28, -128, -128, -116, -128, -127, 81, 127, -53, -128, -128, 65, 68, -17, 23, -128, -128, -116, 23, 65, 127, 127, -7, -101, 23, 91, -128, -128, 95, 127, 52, -128, -128, 33, 127, 127, 127, -60, -106, -114, -128, -128, -59, 29, 3, -92, -128, -92, -42, 47, -88, -10, 127, 127, -45, -60, 127, 127, 32, -13, 127, 127, 42, -32, -29, -114, -54, 10, 49, -128, -128, 98, 127, 127, 45, -53, -21, 127, 98, 79, -128, -11, 127, 127, -128, -128, -127, 0, -10, 7, -128, -111, 75, 127, 36, -24, -34, 5, 39, 127, -2, -121, 80, 127, 127, 15, -75, -44, 36, -6, -78, 21, 13, -128, -81, 52, 114, -36, 76, 127, 127, 127, 1, -91, -102, -71, 127, 127, 106, -128, -128, -109, -128, -128, -88, -18, 112, 127, 127, 127, -13, -59, 109, 117, -79, -128, -100, -128, -59, -128, -128, -128, -117, 66, 71, 0, -74, 90, 97, 127, -57, -128, -128, 127, 92, 6, 103, 127, -90, -128, -128, -80, 28, 96, 127, 44, -50, -32, 88, 15, -74, -16, 127, 107, -95, 15, 127, 102, 52, -101, -124, -128, -128, -71, 127, 45, -128, -128, 0, 36, 122, 127, 102, -3, 127, 127, 127, 65, -33, -128, -128, -101, 127, 127, 60, -76, -128, -128, -116, -68, -52, 127, 127, 13, -85, -59, 21, -95, 42, 59, 127, 37, -128, -128, 116, 127, 69, -87, -128, -128, -107, 116, 127, 127, -128, -102, -17, -128, -128, 52, 127, -36, -128, -12, 68, 58, 87, 127, 127, -122, -128, -21, 127, 0, -91, -128, -128, -119, 80, 43, -128, -112, 38, 127, 74, -39, -60, 12, -43, 85, 127, -85, -128, 71, 127, 57, -128, 6, 127, 127, -65, -128, -128, -54, 127, 127, 22, 52, 127, 107, -128, -116, 74, 27, -121, -106, -88, 68, 127, 71, 8, 127, 127, 68, 70, 28, -69, 57, 90, -128, -128, 117, 127, -17, -128, -128, -8, 86, -37, 39, 127, 127, 11, -29, -128, -128, -128, -128, -119, 21, 98, 107, -24, -128, -128, 87, 127, 118, -96, -128, -128, -128, -128, -128, 127, 127, 74, -93, 39, 127, -103, -128, -87, 13, -59, -79, 68, -49, -128, -53, 29, 127, 127, -107, -128, -121, -33, -66, -128, -128, -86, -28, -128, -128, 37, 22, -16, 127, 127, 22, 98, 26, -128, -128, 43, 127, 127, -76, -49, -39, -17, -128, -106, 60, 122, 32, 71, 127, 112, 60, -49, -128, -65, 92, 127, 127, 127, -3, -86, -112, -114, -128, -88, 71, 2, -128, 10, -39, -16, -108, 8, -23, 127, 66, 38, -85, -101, 28, 127, 127, -59, -3, 74, -128, -128, -38, 127, 123, 121, 127, -71, -123, 127, 127, 127, -91, -128, 79, 127, 127, 43, -93, -128, -34, 127, 127, 10, -128, -75, 5, -13, -3, 38, 49, 74, -79, -59, 54, -58, -31, 87, 127, 127, 127, -8, 5, 118, -16, -128, -128, 12, 85, 127, 33, -128, -47, 127, 127, -23, -18, -48, 50, 88, 127, 127, 127, 49, 13, -16, -128, -114, -78, 6, -128, -128, -128, -80, -15, 5, 127, -78, -128, -128, 53, 112, 38, 55, 127, 127, 127, 98, 54, -100, -128, -128, 127, 127, 127, 31, -87, -128, -128, 127, 96, 38, 127, 127, 79, 91, -44, -128, -101, 127, 127, 127, -39, -128, -128, -128, -18, 127, 108, -128, -128, 102, 127, 118, -36, 127, 127, 48, 17, 1, -1, 34, 2, -109, -6, -95, 98, -18, -5, 31, 127, 101, 87, 123, 127, 1, -52, -53, 95, 5, -127, -80, -128, -93, -45, 3, -128, -111, -128, 2, -48, 64, 33, -127, -81, 107, 121, -5, 43, -128, 111, 127, 127, 127, 53, -98, -113, -8, -91, -128, 11, 73, -124, -66, 127, 127, 108, -111, -128, -128, 59, 127, -90, -128, -7, 59, 5, 117, 58, 16, 26, 15, 118, 91, 127, -8, -128, -128, -128, 55, 106, 98, 117, -42, -7, 90, 54, 127, -2, -12, -42, 36, 74, 106, -48, 36, 127, 50, 13, 15, 17, 59, 127, -10, 68, 127, 127, -128, -87, 127, 87, -118, 64, 127, 127, -10, -128, -128, -21, 127, 127, 53, 21, 32, 70, -60, -73, -119, 60, 127, 127, 66, 68, 18, -38, -128, -128, -128, -80, -5, 45, 127, 54, 0, -128, -64, 44, 127, 127, 127, 124, -128, -128, 26, 68, 24, -128, -128, -124, -57, -128, -106, -128, -128, -128, -6, 111, 127, 71, 98, -128, -108, -88, 11, 43, 112, 127, 127, 127, -24, -111, 48, 127, 127, -128, -128, -128, 26, -18, 13, 127, 70, -29, -128, -128, -128, 73, 27, 29, -37, 90, -37, 116, -15, -128, -128, 90, 127, 127, -36, -128, -90, 73, -91, -128, 0, 93, 39, -32, 90, 15, -128, -38, 127, 2, -128, -128, 52, 127, 127, 127, 3, 91, -28, -128, -128, -68, 12, 27, -98, -128, -128, -128, 55, 127, 127, -2, -128, -42, 127, 127, 31, -122, -76, -1, 127, 127, 127, 127, 58, -52, -15, 127, 127, 98, -106, -128, 48, 127, 127, 29, 47, 127, 17, -128, 26, 127, 53, -57, 69, 127, 1, -69, -24, 23, -76, -47, -38, -128, -128, 37, 127, 127, 127, -36, -128, -128, -80, -112, -47, 18, 65, -24, -34, 28, -34, -107, -97, 90, 118, -27, -128, -128, 5, 127, 101, 32, 127, 54, 28, -93, 50, 113, 127, -13, -128, -128, 127, 127, 127, 127, 127, -128, -128, -68, 44, -27, -76, -64, -45, 66, 127, -63, -42, 37, 78, 54, 127, 127, 73, 54, -8, -123, -91, 42, 55, -74, -106, -37, -54, -85, -128, 123, 127, 127, 69, -128, -128, 52, 127, 2, -128, -128, -128, -29, 88, 6, -98, -10, 31, -90, 50, 5, -128, -128, 119, 127, 127, 69, 26, 8, -33, 113, 127, 127, -128, -128, -128, -70, 127, 127, -101, -128, 59, 127, 127, 74, 127, 108, 107, 48, 79, -50, -128, -128, 37, 86, -128, -128, 127, 127, 28, -111, 71, 107, 17, 54, 63, -128, -107, -53, -5, -128, -128, -128, 59, 127, 127, 57, -128, -128, 127, 127, -119, -128, -69, -42, 108, 123, 127, 92, 127, 127, -80, -74, 69, 28, -128, -52, 124, -50, -128, -71, 24, 90, 85, -80, -128, 127, 127, 127, -26, -52, -124, -49, -38, 13, -102, -128, -123, 3, 26, -38, -128, -32, 80, -93, -116, -49, 3, -23, -106, -121, -128, -1, 86, 102, 92, 107, 54, -31, -34, -33, 68, -1, -128, 101, 127, 127, 127, 32, -128, -128, -128, -29, 127, 127, 95, 113, -29, -78, 127, 127, -33, -128, -98, 86, -23, -128, -128, -128, -118, -73, -7, 127, 119, 0, -78, 6, -23, 103, 127, -50, -76, 127, 127, 49, -8, -29, -128, -128, -128, 34, 127, 127, 39, -24, -128, -112, -6, 22, 73, -22, 116, 127, 127, 96, -71, -128, -128, 17, -128, -128, -127, -95, -74, 64, 127, 127, 111, 69, 90, 113, -33, 97, 112, -42, -128, -70, 127, 127, 127, 97, -100, -33, 69, 24, -100, 29, 127, 127, 127, 86, 127, 59, -124, -128, -114, -32, 127, 127, 127, 28, 43, -113, -85, 27, 127, 15, -128, -28, 127, 50, 33, -54, 5, -45, 36, -38, -36, 13, -78, -63, -18, 127, 106, -1, -74, -128, -128, -58, 127, 109, -27, -128, -73, 13, 80, -128, -128, 127, 127, 38, -128, -128, -54, -48, 127, 17, -59, -109, 127, 127, 47, -17, 127, 127, 127, -128, -128, 38, 71, 0, -16, 7, -106, -64, 23, -128, -128, 27, 127, 127, 127, 127, -59, -128, -112, -55, -65, 5, -88, -80, 127, 127, -97, -74, -49, -128, -128, -128, -74, -13, 127, 109, 127, 116, -11, -128, -86, 92, 29, -16, 65, 103, -42, -92, -31, 73, 127, 90, -87, -18, 1, -18, 45, 79, -103, -112, 127, 127, 127, -33, -113, -114, -123, 68, 18, 32, -18, 127, 127, 66, -128, -93, 12, 95, 127, -28, -128, -26, 127, 24, -128, -128, 127, 127, 127, 118, 36, -23, 74, -102, -128, -111, 127, 127, 127, 32, -128, -128, -128, -21, 127, 127, 65, 17, 12, -15, -79, -31, -75, -23, -16, 86, 116, 58, 86, -76, -87, -70, 127, 127, 127, 28, 64, 22, -128, -116, 127, 127, -128, -128, -16, 127, 127, -58, -128, -128, -16, -6, -128, -128, -7, -12, -128, -128, -128, -113, -121, -128, -128, -128, 64, 107, -31, -128, -32, -122, -128, 0, 127, 127, 63, -81, -85, 119, 127, -1, -39, -57, -86, -112, 37, 127, 127, 96, -55, -16, 45, 73, -96, -128, -128, -128, 75, 127, 113, -100, 109, 127, 28, -128, -128, -36, 8, 74, 76, 98, 78, -80, 42, 55, -128, -128, -90, 97, 124, 73, 16, -44, -128, -128, 127, 127, -1, -128, 127, 127, 24, -128, -88, 127, 127, 34, -128, -128, 23, 127, 127, 122, -44, -64, -128, 24, 44, 118, -128, -128, -75, 127, 127, 29, -48, 50, 127, 106, 127, 127, 79, 17, 68, 103, 78, 127, 127, -128, -128, -128, -24, -55, 60, 127, 127, -75, -128, -128, -111, 12, 127, 127, -44, -95, -106, 38, -81, 45, -42, 127, 116, 127, -2, 64, -39, -90, -128, 90, 113, -3, -60, -128, -128, 58, 127, 127, 7, 66, 127, -23, -128, -17, 127, 100, -68, 78, 127, 127, 79, 127, 127, 81, 127, 127, 93, 71, 127, 127, 39, -66, -128, -128, -33, 127, 127, 127, 127, 81, 37, 45, -38, -128, 121, 127, 73, -128, -119, 127, 127, 114, -93, -128, -128, -116, -69, 127, 127, 45, 38, 54, 54, -65, 54, 32, 36, 127, 127, -91, -32, 127, 127, -12, -96, -128, -128, 65, 127, 127, 53, 1, 96, 127, 127, -37, -128, -128, -107, 49, 127, 127, -128, -128, 23, 127, 127, -27, -128, -128, 113, 127, 127, 81, -12, -128, 78, 127, 52, -16, 0, -21, -128, -87, 107, 127, 93, -111, -70, 76, 127, 127, 127, -128, -128, 12, 127, 127, 127, -85, -128, -80, 127, 127, 36, 88, 127, 127, -24, -128, -52, 90, -47, -3, 127, 127, -74, -128, -128, 52, 65, -63, 6, -16, 54, -50, -75, 60, -128, -128, -60, 127, 127, 124, 127, 127, 127, -8, -63, 22, 127, 43, -8, -112, -128, 15, -49, 50, 127, 127, 127, 127, 127, 106, -53, -128, -65, 127, 93, -127, 121, 127, 42, -96, -91, -128, -128, -32, -117, -128, -128, -45, 47, 11, 53, 127, 102, 69, 70, -97, -128, -92, -128, -116, 92, 127, 127, 127, 78, -27, -128, -128, -90, -38, -17, 127, 26, -128, -128, -128, -70, 0, 127, 127, 12, -128, -113, -21, 21, 76, 127, 127, -8, -128, -66, 87, -17, -128, -96, -118, 52, 127, 127, 127, -128, -128, -28, 85, 79, 66, 68, -93, -107, 2, -54, 11, 7, -121, -11, 37, 13, -45, 32, -103, 31, 127, 22, -128, -23, 91, -128, -128, -24, 127, 127, 127, -128, -128, -76, 59, 100, 127, 127, 127, 86, -81, -128, -70, -53, -128, 86, 127, 76, -128, -128, 60, 70, -43, -81, 127, 127, 127, 127, 127, -108, -128, -12, 127, 1, -3, 73, 127, -10, -16, 23, 111, -79, -91, -36, -59, -128, -128, 53, 127, 127, -128, -128, -128, 3, -15, -23, 91, 127, 27, -119, -60, -70, -128, -128, -18, 127, 127, -43, -128, 23, 127, 127, -74, 28, 127, 88, -128, -128, 65, 111, -23, -128, -5, 127, 127, 108, 102, -39, -128, -128, -54, -128, -128, 127, 127, 127, 127, 43, -124, 76, 127, -17, -128, -128, -76, -8, -124, -100, -64, -128, -128, -113, -27, 127, 127, 127, 49, -100, -128, -95, -32, 127, 127, 127, 102, 55, -47, -128, -48, 127, 88, -128, -128, 73, 127, 127, -101, -128, -28, 127, 127, -15, -43, 127, 127, -52, -128, -79, 127, 127, 127, 127, 12, -122, -80, -59, -64, -64, 127, 127, 127, 108, 27, -128, -128, 42, 127, 127, 127, 109, 26, -54, 18, 127, 127, -60, -128, 17, 127, 47, -98, -7, 55, -48, -49, -128, -128, 24, 127, 117, -128, -18, 127, -43, -128, -128, -128, -27, -78, -68, 96, 127, 127, -11, -2, 93, 127, 17, -1, -27, 3, -128, -128, -32, 127, 127, 127, 31, -128, -128, 13, 127, 21, -128, -101, -32, 100, 127, 127, 117, 65, -6, 34, 127, 58, -85, -26, 73, -128, -128, -101, 127, 127, 7, -128, -128, -97, -128, -128, 68, 121, 87, 21, 16, 38, 127, 127, 127, 127, 127, 44, -7, -80, -74, 57, 101, 90, 59, -78, -128, -128, -88, 50, 39, -93, -128, 71, 127, 127, 127, 127, 127, 127, 60, -128, -33, 127, 127, -128, -128, 15, 127, 127, 70, 18, -78, -128, -128, -124, -103, 118, 127, 127, 97, -128, -38, 127, 71, -128, -128, -128, -88, -45, -128, -33, 127, 127, 29, -128, -128, -128, 5, 127, 127, 127, -34, -128, -128, -128, -128, 47, 127, 127, 127, 127, -76, -65, 60, 127, -28, -128, -73, 127, 127, 53, 58, -112, -128, -73, 127, 127, -118, -128, 64, 127, 48, -128, -128, -92, 127, 127, 127, -116, 7, 127, 127, 127, 80, 127, -17, -128, -128, 16, 71, -128, -128, -70, -2, 44, 90, 127, 117, 127, 122, 60, -54, 6, 127, 127, 87, -29, -69, -128, -128, 127, 127, -73, -88, 53, 13, -128, -128, -128, -128, 0, 127, 109, -15, 42, 66, 31, -2, 114, 53, 127, 127, 127, 101, 16, -128, -128, -58, 55, -85, -128, -128, -128, -48, -18, 50, 127, 92, -128, -128, 52, 111, 116, 127, 127, 121, 127, 114, 6, 97, 127, 71, 28, 108, 122, 96, -128, -86, 64, 127, 50, 55, -27, -26, -128, -128, -71, 122, 118, 76, -10, -92, -128, -74, 16, -66, -128, -65, 127, 127, 111, 12, -128, 28, 127, -128, -128, -128, -39, -52, -81, -64, 55, 98, 127, 91, 127, 127, 127, 74, -112, -128, -44, 79, 79, 127, 39, -128, -128, -18, 73, 69, 33, 5, -96, -74, 26, 127, 127, -64, -23, 127, 127, 127, 112, -92, -128, -128, -68, -128, -128, -12, 38, -98, -111, 98, 127, 127, 59, -7, -103, -12, -128, -128, -128, 123, 127, 8, -43, 31, -70, -128, -23, 127, 127, 127, 127, -128, -128, -128, -128, -128, -106, 127, 127, -27, -128, -128, 33, 127, 127, 127, 60, 87, 71, -23, -128, -65, 95, 44, 127, 37, 70, -128, -128, -111, -3, -74, 2, 32, 53, -26, -112, -128, -28, 127, 80, -128, -128, -75, -36, 92, 127, 81, 36, 1, 0, -128, -96, 59, 17, -50, 52, -128, -128, -128, 103, 127, 59, -128, -6, 127, 31, -38, 127, 127, -53, -76, 88, 127, 6, -59, 85, 13, -128, -128, -53, -128, -123, 127, 127, 28, -31, 26, 55, 127, -91, -128, -128, -2, 88, 79, -48, -128, 1, 58, -95, -128, 29, 127, 127, -75, -128, -76, 58, 15, -23, -28, -128, -101, 114, 17, -128, -128, -128, -128, 22, 127, 95, -75, -128, 96, 91, 11, -100, -113, -128, -90, 65, 112, -107, -128, -76, -49, -128, -128, -5, 127, 127, 1, -107, -128, 111, 127, 95, -128, -57, 127, -34, -128, -128, -128, 75, 127, 21, 2, 127, 127, -128, -128, -70, 127, 127, 127, -42, -74, -102, 11, 93, -11, -128, -128, -128, -28, 127, 127, 127, 109, 44, -73, -21, 1, -49, -44, -45, -73, -1, 127, -3, -107, 10, 13, -29, 45, 127, -1, -13, 37, -2, -128, -85, 34, 123, 22, -47, 78, -57, -74, -128, -124, 68, 127, -128, -128, -74, 23, -22, -128, -128, -128, -76, -38, 16, 116, 38, -128, -128, 23, 79, -70, -128, -128, -128, -81, -123, -128, -111, 73, 8, -6, -28, 127, 127, -22, -128, -117, -45, -128, 54, 127, 88, -27, 59, 74, -39, 114, -3, 26, -64, 127, 127, 127, 10, 0, 57, -95, -121, -13, 127, 127, 127, 22, -128, -24, 101, -29, -102, -11, -10, -128, -128, -39, -24, 74, 127, 127, 78, 127, 127, 127, -31, -128, -128, -96, 100, 107, -17, -13, 127, 32, -47, 127, 113, -86, -28, -1, 78, -50, -128, -128, -128, -12, 127, 127, 38, 127, 127, -7, 22, -10, -128, -128, -127, -39, 101, 97, 71, -118, -21, -60, -106, -128, -79, -75, -128, -128, 127, 127, 127, 60, -71, -128, -81, 127, 127, -47, -128, -128, -128, 15, 127, 127, -128, -128, -36, -15, -108, -128, -106, -6, 127, 92, -128, -6, 127, 80, -128, -128, 127, 127, 127, 117, 127, 127, -31, -128, 0, 127, 127, 127, -45, -96, 66, 127, 44, -78, -95, -128, -85, -107, -39, 111, 127, 127, 73, 42, -21, -50, 117, 127, 127, -38, -124, -117, 43, -38, -37, 127, 127, 54, 0, -66, -101, 127, 127, 50, -11, 32, 22, -128, -111, -97, -122, -80, 87, 70, -57, -34, -128, -128, -31, 127, 18, -64, -48, 27, -128, 24, 127, 27, -128, -2, 127, 85, -59, -87, -128, -128, 18, 45, 5, -128, 5, 33, 17, -128, -128, -128, 127, 127, -21, -128, -128, -63, 122, 127, 127, -49, -63, 11, 127, 127, -128, -128, -16, 127, 127, 98, -128, -128, 2, 123, 3, -50, 85, 127, 127, 127, 127, 127, 127, 6, -128, -112, 43, -2, -80, 43, -8, -128, -103, 127, 127, 127, 121, 119, 59, -128, -128, -128, -64, 22, 74, -64, -92, -91, 127, 48, -128, -39, 127, 127, -6, 6, 127, 127, -128, -128, -128, 18, 119, 127, 127, 31, -27, 53, -33, -38, 100, 47, -128, -108, 49, -1, 55, 85, 68, -128, -128, 26, 127, 26, -87, -114, 28, 127, -12, -128, -123, 127, 127, 50, -128, -128, 23, 76, -47, 42, 127, 127, 31, -32, -65, 127, 127, 127, -128, -107, 0, -98, -128, -128, 63, 119, 127, 127, 78, -39, -13, 38, 16, 127, 103, -128, -128, -128, -65, 69, 127, 91, 0, 127, 127, 127, 93, -88, -128, 17, 113, -22, -103, 127, 127, 74, -128, -128, -128, -128, -13, 27, -13, -128, -102, -85, 98, 127, 127, 53, -128, -128, 127, 127, 127, 127, -11, -128, -128, 127, 127, 96, 71, -54, -76, 45, 113, 71, -119, -58, -88, -65, 39, 127, 127, 127, 95, -128, -128, -128, 127, 127, 59, -50, 127, 127, 91, 50, 87, -73, -113, -128, -32, 1, -13, -128, -93, 127, 127, 127, 11, 69, 60, -70, 52, 118, 124, 32, -60, -128, -128, -128, 2, 74, 58, -53, 80, 69, 106, -107, -128, -37, 36, -69, -116, 127, 127, 48, -47, 22, -100, -80, 127, 127, -121, -128, -48, -93, -109, -128, -128, 16, 127, 127, 27, 127, 127, 122, -128, -45, 127, -18, -128, 54, 127, 127, -127, -128, -98, -2, -34, -32, -16, -128, -128, -121, -8, 74, 48, -128, -128, -128, 80, 57, -69, -58, 69, -22, -128, -32, -54, 15, 3, -128, -128, -128, 45, 90, 127, 127, 42, -128, -81, -60, -66, -36, -117, -128, 21, 127, 127, 45, -128, -21, 23, 43, 21, 127, 0, -78, -48, -11, 38, 102, -36, -112, -128, -124, -122, 11, 127, 96, -36, 127, 127, 18, -52, -43, -128, -7, 127, 127, -34, 75, 127, -48, -128, -128, 48, -47, -128, -26, 127, 103, -54, 15, 127, 127, 109, 12, 42, -55, -128, -128, -117, 0, -13, -128, -29, 101, -112, -128, -128, -128, 21, 127, 127, 36, 34, -65, -31, -95, -116, 3, 52, 127, 127, 85, -38, 127, 127, 22, -18, 17, -52, -128, 17, 63, 31, -7, 127, 108, -128, -112, 39, -5, -63, -3, 127, -108, -128, -128, 124, 117, -34, -8, 112, -22, -128, -123, 127, 2, -128, -128, 127, 127, 33, -68, -18, 70, -7, 36, -7, 29, -33, 32, -21, -34, -17, 3, 8, -128, -128, 127, 8, -128, -128, 127, 127, -28, -128, -128, 43, 16, 81, -53, -45, 111, 127, 33, -128, -3, 111, -128, -128, -45, 69, 58, 127, 127, 127, -47, -68, 32, 98, -44, -128, -128, -28, 127, 127, -26, -54, -24, -37, -128, -21, 116, -97, -128, 119, 127, 112, 85, 66, 29, -85, -128, 63, 123, 127, 127, 74, 50, 106, 108, -122, -87, 65, 69, -33, -28, -124, -108, -21, -59, -24, 17, 127, 127, -47, -88, -128, 127, 127, 127, 114, 71, -76, -117, -28, -128, -128, -26, 127, 127, -128, -128, -37, 64, 45, 116, 127, 3, -8, -128, -128, -128, -21, 127, 127, 127, -76, -128, -128, -76, -64, -86, -107, -52, 127, 0, -128, -128, -128, -128, 90, 127, 65, -128, -17, 127, 11, -88, 34, 113, -128, -128, -128, 88, 127, 36, -122, -17, -31, 122, 127, 127, 127, 127, -47, -123, -128, -128, -128, -64, -68, -128, -128, -114, -128, -114, 127, 127, 127, 85, -38, -63, -60, 22, -27, -75, -128, -128, 32, 8, -128, -102, 127, 12, -128, -117, 10, 127, 127, 127, -128, -128, 75, 127, -75, -128, 15, 127, 78, 33, 33, -78, 64, 127, -109, -128, -17, 127, 127, -128, -128, -59, 127, 127, -100, -128, -128, 73, 127, 127, 127, 1, -119, 5, -3, -128, -128, -119, -68, -128, 10, 127, 45, -128, -128, 33, 47, 103, 122, 39, 127, 127, -27, -128, -117, 66, 127, 127, 87, 127, 127, -66, -128, -128, -121, -85, 127, 44, -60, -128, -128, -50, 97, 53, 33, 0, -36, 106, 127, 127, 121, 32, -75, -73, -111, 78, 127, 127, -128, -128, 22, 29, -128, -128, 23, 127, 127, -29, -128, -128, -128, -76, 100, 127, 55, -113, -127, -36, 13, -21, 6, 127, 127, -78, -109, 98, 127, 107, 26, -128, -91, -76, 107, -39, -79, -128, -3, 11, -36, -24, 3, 127, 122, -32, -73, 16, 114, 127, 54, -36, 2, 74, -69, -128, -128, 50, 127, 127, -7, -128, -73, 24, -42, -128, 98, 127, 118, -96, -113, -128, -58, -34, 127, 90, -128, -128, -128, -128, -117, 74, 127, 127, 127, 79, 21, -28, -113, -128, -128, 53, 127, 37, -91, -128, -57, 15, 127, 48, -128, -7, 127, 81, -80, 3, 86, 24, -106, -128, -128, 127, 127, 127, 127, 127, 34, 27, 90, 127, -112, -128, -121, -7, 78, 36, -128, -7, 127, 127, -74, -90, 80, 127, 90, 22, 15, -96, -59, 117, 127, 117, 127, 86, -96, -128, -128, 127, 127, 127, -15, -98, -128, -68, -45, -128, -128, -128, 85, 75, -21, -128, -44, 23, 24, -71, 64, 127, 15, -111, -128, -128, -107, -103, -128, -128, 6, -103, -128, -24, 127, 127, 70, 66, 37, 26, -128, -88, 127, 127, 127, -16, -128, -122, 75, -96, -128, -128, -66, -71, -48, -97, -128, 18, 127, 49, -128, -128, 18, 73, 127, 86, 13, -23, 65, -26, -128, -128, 58, 127, 127, -24, -39, 70, 112, 49, 31, -74, 93, 114, 127, 78, 127, 92, 39, -74, -11, 124, 127, -128, -2, 127, 76, -128, -107, 29, 39, 127, -22, 111, 127, 127, -22, -31, -36, -128, -128, 45, 100, 127, 78, 63, 80, 127, 127, 102, -109, -32, 127, 127, 5, 13, 71, 127, 79, 6, 43, 109, 68, -11, 127, 127, 8, -73, -16, 127, 127, -33, -128, -58, 85, 127, -71, -128, -128, -69, 32, 75, -97, -128, -128, -128, -98, 127, 127, 127, 15, 1, -23, 44, -8, -48, -38, 28, -128, -128, 34, 127, 127, -86, -128, -116, -128, -128, 15, -102, -128, -48, 127, 127, 49, -69, -22, 5, -12, -111, 113, 127, 123, 7, 103, 127, -60, -128, -128, -128, 75, 127, 39, -128, -128, 123, 127, 24, -7, 127, 111, 78, 113, 127, 76, -76, -50, 127, 127, 21, -128, -128, -128, -55, -128, -128, -128, 23, 127, 127, 64, 57, 127, 90, -128, -128, 127, 127, 127, -27, 81, 127, 127, -1, -65, 53, 127, 127, -93, -128, -128, 59, 127, 127, -128, -128, -33, 22, -128, -38, 127, 127, -37, -128, -108, 127, 127, 127, 127, 127, 18, 47, 113, 6, -128, -128, -128, -128, 127, 127, 127, 96, 108, 27, -43, -68, 74, -65, -57, 63, 111, -53, -128, -128, -76, 127, 109, -128, -128, -39, -39, -73, -10, 49, -42, 98, 127, 127, 55, 28, 50, 60, 71, -45, 7, 127, 127, -106, -128, -128, -128, 34, 127, 31, -128, -121, -10, -128, -128, 65, 38, -128, -128, 33, 53, 39, 127, 127, -48, -128, -96, 127, 127, -2, -49, -48, -128, -101, 127, 127, -91, -128, -16, -31, -128, -128, 39, 127, 78, -128, -128, -74, 13, -44, -75, 127, 91, -71, -128, 59, 108, 127, 79, -73, -59, -49, 7, 101, 127, 127, 48, -48, -21, 122, 123, -7, 49, 127, 107, -63, 92, 127, -64, -55, -128, -128, -128, -128, -73, 127, 53, -128, -128, -38, -15, 75, -2, -128, -54, 127, 127, 95, 118, 127, 70, -93, -128, 36, 127, 127, 127, -66, -128, -128, 79, 127, 127, -102, -128, -128, -128, -18, 17, 127, 127, 127, 127, 127, 6, -15, 127, 127, 127, -91, -128, -60, -128, 78, 71, 23, -121, -100, -124, -122, 57, 70, -75, -128, -63, 127, 22, 0, 127, 127, 27, -128, -128, -11, 0, -44, -53, 32, -128, -128, -119, 24, 127, 127, 76, -91, -128, -128, 127, 127, 47, -75, -128, -116, 42, 49, -128, -128, 22, 127, 47, 44, -128, -128, -128, 127, 127, 23, -128, -22, 127, 127, -88, -128, -128, -128, -88, 127, 127, 75, 0, 64, 127, 38, 111, 79, 127, 109, 127, 44, -74, 91, 127, 127, -93, -111, -71, -102, -34, 78, 127, 64, 91, 116, 53, 96, -97, -128, -85, 127, 127, -128, -128, -78, 127, 127, 59, 17, -29, -60, -96, -27, -3, 95, 8, 127, -8, -59, -117, -43, -93, -18, 127, 127, -17, -128, -128, 0, 114, 127, 127, -78, -128, -27, 64, -21, 127, 66, -66, -128, -49, 88, 97, 127, 127, 64, -86, -57, -22, -16, 93, 43, -121, 2, 10, -117, -78, 28, 22, -32, 59, -15, -128, -128, -128, -128, -128, -97, 127, 127, -8, -128, -128, 127, 127, 116, 38, 38, -108, -69, -31, 127, 127, 118, 44, -52, -119, 23, 69, -3, 50, 23, -128, -128, -3, 74, 6, -1, 127, 127, -128, -127, -33, -21, -128, -114, 16, 127, 127, 113, 29, 127, 127, 127, -76, -128, -128, 2, -36, -128, -128, 127, 127, 15, -128, -128, -6, 123, 127, 55, 13, -79, -11, -128, -114, -127, 53, -60, -75, -29, 127, 127, 86, -128, -24, 127, 33, -109, -49, 91, 22, 65, -15, -13, 54, -29, -70, -43, 33, -13, -24, 127, 127, -7, -80, -128, 91, 127, 127, -28, -128, 13, 127, 68, 70, 127, 127, -118, -128, 10, 127, -38, -128, 91, 127, 127, 124, 5, 63, 127, 101, 73, 127, 60, -60, -119, -60, -128, 6, -42, 119, 127, 127, 127, -5, -128, -128, -128, -68, -66, -95, -65, 64, 2, -128, -128, 0, 65, -109, -128, 32, 127, 97, -128, -128, 66, 64, 96, 127, 127, 16, 23, 31, 48, -121, -128, -128, -98, -39, 92, 50, -128, -128, 127, 85, -128, -128, -79, -76, 79, 127, -27, -128, -128, -128, -18, 11, -128, -128, 127, 127, 33, -66, 38, -36, -74, 127, 95, -95, -76, -128, -128, -117, 0, 22, 127, 127, 127, 42, 127, -7, -128, -128, -15, -102, 6, 127, 127, 23, 119, 70, -74, -122, -118, -26, 127, 127, -66, -128, -128, 127, 0, -128, -128, 17, 127, 59, -128, -128, 127, 127, 12, -101, 29, 127, 107, 102, 53, 86, -17, -98, -128, -60, 21, 127, 127, 47, -128, -81, 7, -15, 38, 127, 45, -128, -92, 22, 127, 95, 58, 48, 127, 65, -128, -59, 45, -122, -128, -5, 15, 127, 127, 127, 127, 127, 95, -48, -98, -128, -68, 71, 75, -76, -44, 48, -53, -128, -111, 127, 127, 13, -107, -68, -117, 39, -5, 31, -63, 44, -123, -58, -128, -12, 18, 23, 127, 127, 127, 8, -128, -7, 127, 28, -107, -38, 85, 10, -24, -128, 48, 127, 127, -108, -86, 13, 127, 127, 10, -128, -128, -128, -128, -45, 127, 54, -128, -128, -102, 75, 79, 127, 59, 0, -128, -128, -128, 0, 6, 26, -45, -24, -74, -128, -65, -34, 12, 127, 127, 123, -55, -128, -128, -123, -3, 90, 127, 127, 7, -60, -50, -27, -128, 26, -10, 38, 50, 127, -71, -128, -128, 34, 91, -59, -47, 127, 88, -47, -128, -128, -128, -128, -128, 26, 127, 127, 87, 127, 48, -17, -43, -78, -128, -128, -1, 58, -65, -121, 74, 127, 127, 127, 127, 16, -21, -70, -44, 127, 86, -128, -128, -128, -128, -108, -116, 74, 127, 127, -66, 34, 127, -12, -128, -128, -102, -21, -26, 50, -128, -128, -128, -128, -75, 26, 101, 38, 113, 21, 75, -39, -106, -128, 86, 127, 127, 127, 127, -18, -91, -42, 11, 22, 55, -32, -13, 127, -32, -128, -6, 98, -6, -128, -75, 1, 2, -13, 127, 127, 71, 95, 127, -57, -128, -28, 127, 127, -66, -128, -47, -24, 53, -47, -37, -34, 127, 118, -98, 29, 79, 0, -65, -55, -109, -86, -2, 119, 127, -13, -28, -7, -118, -128, -58, -91, 11, -21, 1, -8, 127, 127, -28, -66, 27, 36, 127, 49, 44, 96, 127, 127, 113, -128, -117, -95, -128, -128, 66, 127, 127, 127, 100, -128, -128, -96, 106, 127, 127, 54, -3, 34, -68, 73, 127, 127, 109, -27, -128, -128, -128, -128, -128, -121, -13, 0, -65, -18, 127, 0, -127, 29, 91, -31, -54, 116, 127, 127, -29, -117, 12, 113, 127, 127, 127, -128, -128, -90, 73, 127, 127, -86, -47, 52, 127, -36, -128, -93, 96, 76, 91, 127, 127, 96, 45, -26, -2, -24, -39, 15, 127, 45, 37, 127, 127, -128, -128, -128, 87, 127, 127, -17, -34, 121, 127, 127, 109, -85, -128, -111, -78, 6, -86, -66, 28, 39, -64, 34, 127, 127, -16, -27, -18, -24, -128, -128, -18, -128, -31, 127, 127, 127, -121, -128, 85, 127, 127, 127, 127, 127, 127, 34, -128, -119, 96, 119, 127, 60, 127, 127, 92, -118, -128, -128, -53, 127, 127, -71, -128, -128, -7, 127, 127, 60, -36, -71, -128, -18, -34, 5, -70, 15, -97, -95, -55, 102, -50, -107, 43, 73, 127, 127, 107, 127, 127, 76, -13, -112, -13, 101, 127, -54, -128, 6, 102, 97, 15, -127, -128, 3, 71, 127, 127, 127, 127, -26, -128, -128, -76, 47, 48, 97, 116, -65, -128, -128, -49, 107, 127, 66, 127, 29, 127, 127, 127, 57, -78, -128, -23, 127, 127, 127, 81, -43, -24, 127, 127, -58, -18, 92, -11, -128, 5, 18, 49, 12, -48, -90, 28, 117, 127, 127, -112, -128, -122, -52, -128, -128, -128, 80, 127, 127, -69, -128, -128, 127, 127, 127, 22, -42, -128, -128, -81, 63, 127, 87, -128, -128, -43, -21, 28, -26, 123, 39, -2, -123, -128, -128, -128, -60, 127, 127, -8, 58, 127, -53, 28, 127, 127, -13, -128, -128, -128, -76, 127, 127, 92, 45, 113, 127, 92, 111, -128, -128, -15, 127, -91, -128, -128, -26, -86, -42, 127, 127, 114, 96, -10, -128, -128, 103, 127, 33, -128, 119, 127, -3, -128, -128, 127, 127, 127, 127, 108, -88, -90, 39, 86, 112, 10, -49, 33, -96, 73, 127, 121, -128, -128, -119, -128, -128, 127, 127, 124, -128, -81, 127, 127, 127, 70, 73, 52, -3, -66, 127, 127, 90, -91, -128, -128, -76, 127, 127, 7, -128, -113, 127, 127, -75, -128, -128, 92, 42, -128, -128, -128, -128, -128, -31, 127, 85, -97, -112, -31, 44, -69, -128, 23, 127, 127, -128, -128, -127, -47, -98, 15, -32, -85, -87, 127, 127, 68, -90, -92, 50, 127, 127, -68, -116, -27, 39, -66, -128, -106, 80, 127, 127, 6, 11, -31, -69, 69, -45, -128, -128, 108, 127, 127, -5, -11, -23, -109, -17, -50, -98, 42, 127, 34, -128, -128, -73, 70, 123, 53, 31, 127, 81, 22, -128, -128, -124, -36, -92, -86, 0, 64, -128, -128, -34, 127, 127, 127, 127, 81, -60, 47, 127, 127, -27, -128, -128, -22, 127, 34, -128, -128, 28, 102, 8, -86, -87, 49, 45, 93, -107, -128, -11, 17, -128, -128, -49, -37, -128, -123, 127, 127, -76, -32, -93, -128, -128, -128, 121, 127, 127, -128, -128, 28, 2, 93, 101, 90, -42, 96, -5, -128, -128, -128, -128, 59, 127, 91, -128, -128, -122, -128, -128, -50, 75, 26, -91, -31, 1, -69, -128, -22, 127, 127, 127, 49, -128, -128, -128, -85, 116, 127, -71, -128, -57, 127, 127, 127, -33, -128, -106, 78, 66, -116, -128, -63, 102, 127, 127, 98, -128, -12, 127, 39, -128, -70, -23, -128, -128, -1, -93, -117, 58, 71, -117, -27, 127, 127, 123, 23, 0, 12, 21, -116, -128, -128, -109, -58, 68, 127, 38, -71, -32, 127, 127, 127, -39, -128, -128, -95, -26, -128, -128, 127, 127, 71, -43, 127, 127, 31, -100, -23, 101, 79, -86, -79, -38, -48, 127, 127, 127, 127, 127, 32, -16, -31, 16, 127, 95, -22, 119, 127, -128, -128, 0, 91, -65, -128, -128, -128, -128, -128, 109, 127, 127, 44, 8, -8, 34, 127, 127, -128, -128, -122, -117, -128, -128, -128, -106, 5, -13, -128, -128, 88, 127, 0, -68, -3, 127, 127, 124, -128, -128, -128, -23, -128, -128, -128, 108, 127, -29, -128, -128, 36, -47, -128, -123, -122, -7, 5, -128, -128, 50, 123, 28, 68, -45, -37, -128, -128, -128, -128, 3, 127, 127, 97, -98, -66, 45, 68, -87, -128, -128, -55, 55, 127, 127, 127, -42, 59, 127, 127, 127, -8, -128, -128, 92, 43, -21, -11, -52, -128, 59, 127, 127, -54, -119, -90, 43, -5, -12, 60, 76, -53, 34, 85, -88, -117, -90, -92, -69, 103, -128, -128, -128, -16, 97, -36, -128, -91, -12, -31, 127, 88, 127, 127, 127, 11, -128, -78, -42, -54, -128, -128, -42, -36, 37, -55, 70, 13, 50, 64, 127, 127, -36, -69, -128, -128, -128, 76, 127, 127, -11, 26, 127, 127, 127, 127, 127, 2, -92, 80, 127, 127, 127, 113, 127, 127, 127, 76, -128, -128, -10, 54, 95, 127, 21, -128, -128, -17, 127, 127, 121, 127, 60, 42, 44, 44, 73, 75, 111, -65, -121, 44, 127, -71, -128, -16, 127, 102, -128, -128, -73, -128, -128, 124, 121, -31, -128, -128, -128, 112, 127, 127, 47, -26, 75, 124, -128, -128, -21, 0, -88, -36, -3, -111, 0, 63, -26, -33, -22, -74, -118, -128, -128, -45, -117, -128, 12, 127, 127, 10, 68, 127, 74, 55, 63, 127, 98, 127, 93, 71, -96, -128, -128, -106, -49, -65, -128, -108, 17, 118, -75, -128, 80, 127, 127, 8, -128, -128, 122, 127, 127, -103, -32, 127, 59, 26, 71, 5, -128, -63, 127, 127, 3, -17, 32, 93, 42, 28, -128, -128, 108, 37, -75, -42, -27, -80, 127, 127, -34, -128, -128, -128, -128, 1, 127, 127, 127, 38, -128, -43, 127, 119, -128, -8, 127, 127, 23, -128, -128, -128, -109, 10, 127, 127, 127, -15, -128, 26, 127, 127, 127, 127, 127, 44, -128, -128, -128, -128, -128, -127, -128, -128, -64, 127, 127, 71, 12, 127, 127, 127, 60, 70, 5, -34, 112, 33, -29, 22, 127, -29, -71, 31, 127, 127, 23, -85, 1, 127, 127, -17, 21, 91, -17, -128, -55, 117, 127, 85, -73, -93, 16, 66, 5, 127, 127, 68, -128, -71, 127, 127, 97, 127, 127, 95, -59, -128, -128, -128, -76, 106, 127, 43, 23, 127, 127, 87, -3, -13, 6, 1, -90, 53, 3, -128, -63, -50, -118, -128, -128, 36, 127, 127, -6, -80, -49, 54, -59, -128, -117, -85, 73, 28, -106, -108, 127, 127, -124, -128, -128, -64, 95, 127, 127, 127, 29, 13, 12, -48, -128, -97, 127, 127, 121, -81, -128, -128, -60, 80, 68, -42, -128, -127, -59, 88, 127, 127, -24, -128, -97, -17, -128, -128, 29, -13, -128, -54, -88, 22, -81, -128, -7, 127, 88, -109, -117, -128, -128, -63, -15, -23, -96, 100, 127, 127, 127, -90, -128, -53, 127, 127, 53, 7, -7, 117, 95, -15, -112, -128, 49, 60, 45, 17, 127, 127, 127, 71, 23, -81, -66, -128, -85, -42, 92, 75, 22, 18, 44, 127, 28, 117, 127, 64, 6, -128, -128, 12, 127, 85, -128, -11, 112, -23, -128, 127, 127, 127, 69, 39, 108, 49, -106, -128, -128, -128, -37, 34, 119, 127, -24, 23, 127, 97, -128, -128, 10, 127, -65, -128, -16, 127, 127, 102, 23, -44, -128, -128, -128, -128, -22, 127, 127, 66, -47, -128, -122, -21, -95, -128, -128, -128, 34, 55, 121, 127, 43, -128, -79, 108, 74, -27, 103, 48, -128, -112, -36, 123, 31, -128, -128, -7, 127, 24, -128, 48, 127, 87, -75, 39, 127, 111, -6, -121, -128, -128, 44, 127, 127, 10, -119, -95, 45, 127, -128, -128, 27, 127, 33, -128, -128, -79, -128, -128, 81, 127, 101, -128, 10, 127, 127, -21, -71, -121, 38, 117, 123, 127, 127, 49, -128, -128, -66, -7, -80, -6, -65, 0, -52, -21, -91, -128, -28, 44, -52, 122, 127, 127, 92, 127, 127, -31, -100, 54, 127, 74, -98, -128, -68, -128, -128, -112, 127, 127, 8, -128, -128, -128, -128, 13, -17, -32, -71, 2, -128, -100, -28, -18, -128, -128, -128, -22, 8, -8, 32, 127, -42, -128, -128, 127, 127, 127, 92, 69, 21, 85, 127, 37, 8, -13, 127, 127, 11, -128, -128, -128, -128, 42, 127, 12, -102, -52, -13, -23, 127, 127, -128, -128, -128, 127, 118, -31, -13, 127, -47, -128, -128, -128, -128, -128, -18, 63, 64, -65, -53, 87, 127, -13, -128, -18, 34, -80, -128, -34, -68, -128, -86, 17, -98, -128, -22, 127, 127, 127, 36, -91, -117, -128, -128, 1, 127, 0, -128, -128, 54, 11, -123, -118, 1, -69, -128, -21, 127, 127, -33, -128, 27, 127, 127, -103, -128, -128, 33, 108, 127, 101, -96, 98, 127, 127, 127, 127, 118, 93, 60, 17, -93, -18, 127, 49, -39, 54, 36, -124, -128, 13, 88, 127, -100, -45, 7, 31, -128, -128, -128, 55, 108, 127, 5, -128, -128, 127, 127, 69, -15, 16, -45, -128, 5, 127, 127, 23, -128, -128, -39, 127, 127, -128, -128, -79, 127, 93, -90, 5, 127, 127, 127, -90, -87, 27, 13, -97, 52, 93, -49, 43, 12, -8, -128, 80, 127, 17, 29, 127, 127, 127, -24, -128, -128, -86, -58, -116, -48, -128, -122, 28, 127, 81, -128, -128, 10, 127, -11, -128, -128, 71, 63, -111, -93, -27, 93, 55, 13, -90, -50, 98, 127, 127, 127, 127, 127, 44, -128, -128, -128, 3, -38, -43, -98, -74, -59, 16, -43, -128, -128, 24, 11, 38, 109, 53, -60, 33, 53, 5, 127, 127, -42, -68, -53, 37, 118, 127, 127, 127, 34, -63, -52, -39, -111, -112, -8, -86, -128, -128, -2, 127, 127, -13, 32, 92, 127, 58, 106, 127, 85, -128, -91, -38, -109, -68, -21, -106, -116, -100, 101, 127, 127, 127, 127, 122, 0, 127, 127, 27, -128, -128, -103, 127, 127, 78, -128, 18, 127, 127, 8, 18, 127, 127, -128, -128, -8, 127, 127, 111, -95, -128, -91, 127, 127, 127, -75, -128, -128, -33, 65, 92, 79, 118, 127, 127, 127, 127, 29, -111, -32, 31, 59, 39, 119, 3, -116, -128, -128, 92, 53, -55, -100, -128, -128, 54, 116, -53, -128, -128, 79, 127, 127, -5, 49, 127, 127, -50, -44, 127, 81, -117, -71, 29, 27, 27, 112, 127, 12, -128, -87, -33, -54, -58, -17, 7, -90, -58, -114, 81, -59, -90, -27, 69, 64, 43, 48, -123, -32, 127, 127, -12, -128, -85, 127, 127, 127, 127, -96, -128, -111, 18, -50, -128, -39, -11, 127, 127, 36, -52, -128, -128, -128, -128, 16, 127, 24, -128, -64, -128, -128, -32, 127, -27, -118, 6, -47, -128, 113, 127, 17, -128, -128, -128, -24, 91, 100, 21, 53, -58, -128, -128, 127, 127, 127, -32, -114, 29, 127, 127, 127, 54, -95, -128, -21, 127, 127, -93, -128, -59, 102, 22, 11, 100, 124, 127, 33, -123, -60, 90, 127, 127, 5, -128, 48, 127, 12, -74, 58, 65, -128, -128, -95, 1, 127, 68, 88, 26, 64, -36, 93, 59, 76, 21, 55, -36, -33, -128, -128, -21, 127, 127, 97, -95, -123, -74, 78, 55, -108, -26, 127, 127, -57, 28, -47, -128, -121, 53, 57, -32, 21, -128, -108, 36, 127, 127, 127, 127, 21, -128, -128, -79, 7, 69, -15, 92, 26, -128, -128, -128, -73, -34, -128, -88, 127, 57, -128, 47, 127, 123, 32, 112, 17, -128, -128, -128, 127, 127, 127, -128, -128, -114, 116, 127, 102, 91, 127, 127, 127, 127, -12, -128, -119, -38, -49, 53, 127, 127, 127, 90, -16, 127, 127, -22, -128, -128, 127, 127, 127, 127, 127, 55, -103, -128, -128, -128, -33, 127, 127, -81, -128, -117, -34, -122, -75, -85, 106, 127, 127, -128, -64, 127, 127, -16, -128, -128, -53, 71, -23, -128, -128, -26, 127, 127, -7, -33, 118, 127, 0, 34, 117, -118, -128, 18, 58, -80, 42, 127, -26, -21, 127, 127, -63, -39, -107, -128, 122, 127, 127, -98, -80, 85, 127, 36, -97, -128, -58, -68, -106, -103, 113, 127, 127, 109, 97, -96, -38, 127, 53, -128, -128, 123, 69, -39, -21, 64, -31, -92, -36, 127, 90, 103, -70, -128, -128, -45, 127, 47, -73, -12, 17, 0, -24, -101, 123, 127, 127, 127, 127, 42, 65, 127, -97, -128, -108, 34, -128, -128, -98, -16, 127, 127, 13, -128, -128, -107, -103, 3, -114, -47, 127, 127, 5, 68, 80, -118, -128, -128, -128, -128, -123, -6, 68, -49, -128, -32, 96, -13, -69, -128, -128, -95, 90, 37, -12, 127, 11, -128, -128, 7, 127, 127, 47, -128, -87, 59, -8, -128, -128, -128, -128, -128, -128, -128, -49, -12, -79, -128, -27, 97, -8, -128, -66, 97, 64, -5, 11, -85, -70, -64, -128, -128, -28, 127, 80, 33, 127, 127, 127, 7, 11, 8, -29, -128, -128, -128, -60, 127, 127, 80, -49, -28, 95, 80, -128, -128, -86, 6, 28, -2, 127, 127, 127, 122, 127, 127, 127, 36, -86, -37, 108, -26, -128, -124, 107, 127, 127, -52, -119, -128, 26, 127, 127, 60, 103, -29, 1, 127, 116, -128, -73, -1, -128, -128, -128, -128, -128, 75, 127, 60, 85, 112, -27, -128, -10, -37, -128, -91, 63, 57, 127, 127, 121, -86, -128, -128, -59, 29, 127, 127, 3, -128, -128, -48, 127, 127, -128, -128, -128, -128, -92, -128, -78, -13, -52, 68, 127, 31, 70, 127, 123, 127, -44, -128, -128, 127, 127, 127, 88, -8, -1, -34, 87, -3, -128, -128, -23, 127, 127, 52, -44, -109, 37, 86, 28, 127, 12, -97, -7, 127, 127, 23, 10, 38, 21, 44, -1, -48, -128, -43, 127, 127, -11, 92, 127, 59, -128, -68, 91, 91, 24, 127, -85, -128, -128, -128, -128, -128, -128, -128, -34, -7, 127, 127, 127, 127, 127, -23, -128, -24, 127, 12, 2, 127, 127, 1, 127, 127, 127, 127, 63, -121, -54, 93, 127, -5, -36, -28, 127, 44, -128, -101, 21, 116, 26, 70, -1, -45, -128, -2, 13, -117, -3, 127, 127, 53, 76, -7, -128, -128, -17, -24, -128, -128, 52, 112, 70, 5, 18, 42, 111, 127, 16, 102, 127, 45, -128, -92, -5, -34, -79, -10, -128, 13, 127, 127, 127, 127, -128, -128, 8, 127, 34, 16, 66, 45, -128, -100, 38, -76, -128, -26, 11, -59, -23, 127, 127, 127, 127, 85, -45, 74, 127, 127, 127, 127, 127, 127, -31, -128, -128, 69, 127, -60, -128, -24, 127, -80, -128, 17, 127, 127, -50, -78, 74, 127, 127, 47, -102, 5, 127, -3, -63, 109, 127, -31, -12, 127, 123, -38, 79, 69, -128, -128, -50, 47, 106, 18, -66, -117, -128, -128, -43, -2, -59, 1, 127, 127, -68, -128, -128, 127, 127, 96, -128, -128, -128, -13, -11, -106, -128, -128, -128, -128, -128, -27, 23, -100, -128, 6, 127, 127, 127, 71, 22, 42, 26, -34, 92, 12, -80, -128, -128, -66, 32, 127, 127, 53, 45, 111, 34, -101, -128, -128, 1, 127, 24, -73, 74, 127, 127, 87, 107, 80, 111, -74, -128, -128, -128, -102, -96, -128, -44, 123, 45, -15, 127, 45, -128, -128, -48, 29, 98, 17, -128, -128, -28, 127, -7, -87, 50, -58, -128, 31, 127, 91, -128, -68, -112, 66, -54, -36, -38, 127, 97, -91, -15, 47, -8, -128, -128, -43, 0, 87, 60, 31, -128, -26, 38, -65, -128, -5, 31, 114, 112, 13, -123, -81, 127, 92, 33, -73, 22, 113, -55, -128, 22, 127, -17, -128, -128, -128, -128, 8, 5, 10, 116, 31, -128, -128, -91, 90, 127, 127, 127, 127, 45, -119, 24, 127, 85, -121, -127, 44, 98, 122, -43, 24, 127, 127, 127, 42, -128, -128, -128, -64, -60, -54, -128, -73, -88, 6, 17, 127, 127, 29, -128, -128, 127, 127, 52, -128, -128, 127, 127, 127, 127, 127, -75, -128, -128, 1, 43, 63, -128, -128, -128, 43, 38, 76, 10, -103, -128, -128, 15, 90, -69, -128, 69, 127, -16, -57, 91, 23, -128, -128, -85, 127, 127, 127, 116, -113, -128, -128, 0, 13, -117, -128, -55, 127, 24, -37, 79, 49, -111, -26, -15, 5, -128, -128, -42, -3, 91, 91, 127, 127, 127, 127, -57, -119, 26, 127, 127, 127, 127, -49, -90, -29, -63, -128, -59, 127, 127, 127, 127, 121, 127, -55, -128, -128, 127, 127, -47, -128, -128, 127, 127, 0, -128, -81, -58, -128, -128, -43, 127, 65, -97, -90, -11, -49, 116, 116, 16, -68, 97, 93, 55, -65, -31, 37, -10, -21, -52, -128, -22, -123, 0, 127, 127, 127, 127, 47, -128, 11, 127, 127, 127, 5, -3, 127, 127, -128, -128, -73, 28, -81, -81, 1, -124, -128, 26, 127, 90, -85, -128, -123, 102, 63, -108, -128, 26, 31, 127, 127, 92, -128, -128, 127, 127, 127, 127, 127, 127, 0, 17, 0, -128, -98, 66, 36, -128, -128, 43, 74, -76, -64, 60, 48, -50, -32, -23, 108, 107, -98, -95, -74, 127, 37, -128, -128, 49, 127, 127, 118, 127, 87, -128, -128, -106, 79, 53, -100, -112, -128, -112, -59, 5, -128, -128, -128, 127, 127, -13, -128, -24, -75, -75, 26, 100, 8, -66, 127, 127, 107, -128, -7, 85, -118, -128, -128, -128, -68, 101, 124, 0, -111, -31, -75, 37, 23, 127, 127, 127, 127, 111, 15, 10, 6, 8, -98, -128, -24, 118, -13, -128, -47, 79, 17, -21, -124, -128, -59, 71, -74, -123, 127, 127, 127, 127, 127, 81, 24, -128, -128, -68, -21, -21, -64, 127, 127, 44, -128, -88, 60, -22, -87, 48, -12, -47, -66, 88, 127, 127, -106, -128, -128, 127, 127, 127, 124, 11, -128, -128, 29, 102, 127, 103, 127, 127, 127, 32, 66, 59, -52, -128, -128, -128, 79, 26, -57, -16, 127, 127, -71, -128, -128, -95, 7, 127, 127, 127, 52, 127, 127, 127, 81, -116, -128, 8, 127, 127, 127, 127, 127, 117, 0, -118, -42, -55, -97, -128, -128, -119, 127, 127, 127, 106, 127, 127, 127, -12, -36, -71, -128, -106, 17, -63, 69, 127, 127, -128, -128, -128, -100, -26, 127, 127, 127, 43, 127, 127, 18, 127, 127, 127, 57, 53, 114, 127, 90, -45, -73, -3, 15, 127, 86, -57, -57, -57, 108, 127, 37, -117, 63, 127, 127, 15, -128, -128, -128, 90, 127, 48, -121, -55, 1, -37, 127, 127, 10, -128, -128, -88, -128, 86, 127, 127, -48, -102, -76, -86, -128, -128, -6, -53, -15, -53, 23, -97, -98, -128, -128, -12, -2, -68, -64, -64, -47, 117, 81, -23, 127, 127, 111, -15, -85, -103, -123, -103, 86, 127, 127, 106, 3, -29, -128, -128, 39, 127, 127, 121, 127, 119, 63, 6, 28, 91, 127, 127, -15, -107, -91, -7, 11, -18, -85, -49, -100, 79, 127, 127, 127, 79, 111, 127, 31, 48, 114, -3, -128, -128, -128, -128, -11, 6, 2, -128, -123, -128, 81, 127, 127, -128, -121, 127, 112, -128, -128, -53, 106, 127, 127, 127, 15, -128, -128, -116, 127, 127, 127, 127, 97, -8, -47, -26, 76, 127, 127, -98, -36, 127, 127, -128, -128, -128, -98, -13, -53, 16, 127, 118, -118, -91, 37, 71, -24, 22, -128, -128, -128, -128, -128, 108, 127, 36, -128, -128, -86, -116, -3, 70, 13, 8, -88, 39, -119, 8, 80, 127, -8, -128, 65, 127, 71, -128, -128, -90, -128, -33, 127, -34, -128, -128, -29, -39, -34, -128, 24, 118, 127, 15, -28, 49, 27, -128, -54, 42, 93, -98, -50, 29, 90, -122, -97, -69, 121, 38, -24, 57, 57, 31, 127, 107, -128, -54, 127, 127, 54, -28, -113, -128, -128, 101, 127, 127, 127, -1, -128, 26, 127, 127, 3, -1, -65, -128, -66, 1, 12, 49, 127, 127, 100, -128, -128, -108, 127, 127, 127, -28, -128, -128, 49, 109, -33, -128, -128, -90, 18, 15, -128, -128, -65, -108, 5, 60, -5, -128, -128, -12, 127, 119, 7, -18, -55, -128, 112, 109, 42, -128, -87, 18, 127, 127, 58, 107, 74, 113, 21, -118, -3, 33, -111, -128, 6, -26, -128, -128, -119, 74, 127, 127, 127, 127, -96, -128, 0, 127, -36, -128, -128, -74, 13, 124, 127, 127, 127, 23, -107, 36, 73, -128, -128, -86, -109, -68, 16, -123, 10, 127, 60, -22, 26, -33, -34, 69, -121, -128, -128, 43, 127, 127, -23, -38, 50, 88, -128, -106, 48, 127, 91, 79, -54, -34, 1, 80, 127, 127, -49, -128, -128, 60, 127, 127, 45, -88, -128, -128, 48, 127, 100, -24, 39, 12, -57, -93, 102, 37, 23, 113, 122, -37, -11, 127, 127, 90, 127, 5, -128, -122, -49, -49, -100, -42, 38, 127, 68, -119, -128, -128, -128, -26, -24, -13, 91, 127, 80, -128, -113, -16, -7, -24, -60, -128, -128, 68, 127, 17, -102, 15, 1, -128, -111, -128, 2, -33, -128, -128, 127, 127, -68, -128, -128, 113, 106, 0, -103, 47, -73, -128, -128, -128, -113, -109, -128, -128, 26, 127, 8, -128, -118, 63, 127, 127, -10, -85, -42, 98, 127, 17, -128, -128, 34, 127, 127, 53, -49, -128, -128, -66, 68, 114, 31, -92, -128, -128, -90, -119, -128, -128, -128, -95, -128, -128, -128, 85, 127, 127, 90, 107, 24, -128, -128, -128, -88, -1, 79, 127, 70, -102, -128, -128, 65, 93, -128, -128, -2, 127, 66, -92, 13, 63, 81, 127, 102, -5, -102, -29, 2, -1, -128, -5, -36, -128, -128, -128, 21, 127, 127, 8, -52, 50, 127, 97, 16, 127, 127, -2, -98, -128, -128, -128, -128, -128, -128, 76, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -96, 96, -2, -114, -68, 42, -43, -90, 33, -123, -45, 127, 127, 127, -34, -128, -128, -43, -12, -128, -70, -31, 127, 127, 27, 87, 2, -128, -128, -10, 127, -18, -128, -128, -128, -124, -92, -18, 127, 111, -128, -128, 55, 71, -128, -128, 64, 121, -113, -128, -128, -128, -128, -128, -90, 59, 12, -128, -100, 127, 127, -116, -98, -26, 127, 127, 127, -53, -128, -128, -128, -128, -108, -109, -128, -109, -92, 114, 127, 127, -16, -128, -101, 65, -17, -124, -128, 127, 127, -52, -64, 117, -69, -128, -128, -117, -2, 6, 21, -69, -128, -128, -118, -106, -16, 95, -11, -128, -78, 33, 76, 32, 66, 127, 127, 127, 127, 127, 127, 24, -76, -24, 100, 74, 0, 64, 127, 127, 127, 39, -119, -60, 36, 21, -114, -128, -123, 98, 75, 10, 3, 53, 127, 127, 127, -75, -128, -128, 17, -100, -128, -27, 31, -128, -128, 127, 127, 76, 96, 127, 127, -79, -128, -128, 118, 127, 127, -128, -128, -23, -106, -95, 27, -10, -128, -128, -128, -10, 127, 127, 57, -48, -49, -60, 127, 127, 127, 127, -16, -91, -128, -128, -128, 127, 127, 45, -31, -127, -128, -128, -11, 127, 109, 119, 69, 127, 49, 127, 127, 127, -50, -128, -128, -128, -121, -128, -70, -3, 70, 66, 127, 127, 117, -128, -128, -81, -21, 18, 43, 29, -65, -87, -128, -81, 0, 127, 127, 122, 127, 127, 39, 26, -44, -37, -123, 127, 127, -8, -95, 107, 113, -15, 74, 38, -95, 43, 127, 127, 117, -128, -114, 0, 53, -33, -128, -128, -70, 127, 127, -39, -121, -65, -97, 27, 127, 80, -128, -128, -128, -128, -128, -15, 127, 111, -128, -128, -66, 127, 127, 69, -95, -128, -128, 52, 127, 112, -128, -70, -38, 7, -36, 58, 31, 88, -3, -12, -1, -117, -128, -128, 47, 127, 127, -45, -128, -87, -18, -59, 0, 127, 127, 127, 81, -78, -128, -128, 118, 127, 127, -47, 29, 78, -102, -128, -128, 127, 76, -128, -128, 127, 127, 127, 17, -53, 66, 127, 127, 127, -10, -128, -128, -128, 127, 127, 36, -128, -16, 127, 127, 68, -42, -98, 6, -3, -128, -128, -116, -55, 57, 90, 44, 107, 23, 127, 18, -128, -128, -66, -121, -58, -15, -42, -128, -128, 44, 127, 127, 127, 127, 127, 127, -64, -128, -31, 92, 13, 27, 127, 127, 68, -128, -128, -117, -2, 127, 53, 33, -39, -128, -128, -18, 127, 127, 123, 127, -128, -128, -90, 127, 127, 18, -70, 93, 127, -97, -128, -124, 127, 127, -17, -128, -39, 127, 127, 54, 114, 127, 127, -31, -36, 127, 127, 127, 24, -23, 73, 88, 24, -11, 111, 127, 127, 127, 54, -98, -128, -128, -121, -88, -117, 23, 93, 127, 127, 127, 127, -17, -128, -128, 96, 127, -97, -128, 22, 127, 127, -68, -128, -44, 66, 65, 69, -116, -128, -128, -128, -128, -8, 69, 123, 127, 127, -55, -29, 33, -12, -128, -128, 60, 127, -12, -128, -107, 71, -69, -78, -21, -93, -128, -70, 63, -50, -128, -85, 38, 24, -55, 42, 34, -75, -128, -128, -90, 101, 13, -128, -117, -5, -27, 18, -80, -97, -128, -53, -95, -55, 93, -55, -116, 81, 127, 127, -128, -128, -116, -49, 24, 48, 127, 127, 121, -16, -22, -22, -74, -65, -86, -128, 76, 85, 58, -123, -33, -87, -128, -123, -80, -117, -128, -70, -128, -128, -128, -80, 91, -31, -128, -119, 13, 95, 109, -87, -128, -122, -128, -106, 39, 12, 54, 127, 8, -128, -10, 127, 121, 127, 127, 127, 108, -117, -128, -128, -128, -69, 52, -103, -128, -107, -23, 7, 2, -86, -128, -103, 69, 127, 119, 13, 102, 127, 127, 8, -128, -87, 57, 124, 127, 93, -73, -106, -15, -59, 16, 54, 78, 65, -119, -128, -109, 127, 127, -66, -128, -128, -71, -45, -128, -111, -54, 79, 60, 34, -96, 2, 3, -3, -128, 39, 38, 114, 127, 127, -80, 31, 127, 127, 127, 127, 39, -128, -128, -122, -113, 64, 127, 95, -128, -128, 29, -21, -128, -60, 33, -114, -128, -109, -128, -128, -22, 78, 70, 127, 127, 127, 37, 15, 88, 5, -68, 47, 127, 127, 63, -128, -128, -128, -128, -38, -18, -113, 33, 93, 68, -81, 13, -65, -13, 44, 127, 127, -54, -64, 42, 71, -128, -128, 21, 101, -79, -128, -128, -92, -50, -93, -106, -88, -23, 70, 127, 87, -128, -128, -128, -106, 22, 127, 127, 127, -11, -18, -107, -128, -128, -128, 127, 117, -69, -44, 118, 127, 2, -96, -128, -81, 127, 127, 127, 127, 127, 117, -16, -128, -128, -27, -128, -128, 93, 32, 36, 127, 116, -108, 16, 127, 127, 37, -103, 22, 34, -128, -117, 52, -58, -52, 127, 57, -128, -53, 18, -128, -128, -80, -34, 118, 127, 127, -128, -107, 127, 75, -49, 127, 102, -128, -128, 93, 127, 127, 127, -7, 5, 26, 58, -8, 68, -26, 73, 23, 65, -109, -55, 127, 127, 45, 11, -75, 117, 127, 127, 127, 127, 118, -128, -128, 55, 127, 127, -23, -101, -128, 2, 93, 31, 6, 127, 127, -33, -34, 127, 127, 33, -98, -128, -128, -128, 92, 127, 127, -103, -128, -66, -54, -128, -28, -42, -122, -128, -32, 0, -24, -16, -38, -2, 37, -3, 16, 75, 54, -17, -75, -123, -6, 59, 79, 0, -97, -86, -128, -128, 78, 66, 5, 127, 23, -128, -36, 127, 91, -128, -128, -10, 76, -18, -128, -128, -128, -55, -24, 17, 65, -59, -128, -128, 45, -88, -81, 63, 13, -128, -12, 127, 127, 73, 33, 32, -127, -128, -128, -68, 97, 103, 45, -128, 32, 6, -128, -128, -1, 127, 127, -10, 43, 13, -18, -128, -103, -119, 24, 93, 100, -128, -128, -128, -5, -63, -128, -128, 127, 127, 87, -79, -45, 127, 124, -128, -128, 31, 37, 127, 127, 79, -128, -128, -28, 12, 127, 74, 27, -68, -128, -128, 86, -1, -128, -128, -54, 127, 45, -128, -128, -128, 27, 127, 127, -26, -128, 1, 127, 127, 32, 81, -43, -128, -119, 58, -53, -71, 101, -1, 2, 24, 53, -128, 55, 101, 127, 90, 127, 37, -128, -128, -128, -128, -128, -6, 123, 127, -43, -128, -128, -75, -34, -69, -36, -27, 122, 127, 127, -69, -128, -128, -127, -128, -128, -128, -128, -128, -48, 127, 127, 90, -128, -128, -128, -128, -128, -113, 24, 127, 127, 127, 88, -27, -128, -55, -28, -123, -128, 95, 127, 127, 88, -75, -128, -123, 127, 127, 109, -23, 74, 74, -27, -24, -60, -128, -128, 47, 58, -58, -79, -33, -17, 48, -17, -91, -128, -128, -107, -118, -53, -113, -108, -54, 12, 13, 73, 119, 100, -128, -128, -53, 127, 127, 127, -36, -114, 53, 127, -29, -128, -122, 103, 102, 97, -76, -78, -102, 17, -64, -95, -96, -15, -37, -29, -11, 103, 127, 127, 5, -78, 32, 87, 109, -128, -93, -15, 88, -2, -101, -128, 7, -53, -128, -128, -128, -128, 49, 127, 127, 86, 59, 47, -38, 88, 127, 127, 85, -90, -18, -38, -80, -80, 88, -7, -128, 73, 127, 127, 127, -6, -100, -26, 76, -22, -98, 23, 127, 127, -8, -128, -128, -48, -123, -128, -128, -128, -100, -29, -50, -102, 16, 127, 127, -52, -24, 63, -12, -128, -114, -117, -128, 1, -59, 31, 127, 127, -26, -128, -59, 127, 127, 127, -55, -128, -128, -106, 11, 65, 127, 65, 45, -55, -29, 38, 127, 127, 69, -73, 6, 42, -96, -128, -108, -58, 2, 127, 127, 21, -43, 119, 127, -54, 8, 127, 127, 127, -11, -128, -59, 124, -47, -74, 0, 106, -52, 28, 34, 127, 85, 101, 86, 42, -16, -78, -128, -128, 78, 57, 16, -12, -103, -128, 119, 127, 127, 127, 127, -128, -128, -128, -8, -6, -106, 22, 127, 127, -65, 33, 127, 127, 17, 127, 127, -66, -128, -128, 102, 127, 0, -128, -128, -128, -96, 43, 127, 127, 27, -28, 15, 76, 96, 111, 118, 122, -128, -54, -10, 31, -10, 127, 127, 102, -11, -86, -128, -66, 12, 80, 48, 29, 78, 69, 68, 98, 74, -107, -128, -11, 127, 127, 70, 0, -88, -122, -73, 97, 127, 127, 127, 127, 127, 91, -75, -128, -128, -128, -17, -27, -7, 29, -49, -3, 127, 127, -32, -128, -128, 69, 127, 127, 15, -96, -44, 127, 80, 50, -128, -128, -70, -65, -124, -128, -86, -87, 21, 127, 127, -78, -128, -128, -12, -50, -39, 112, 38, -128, 47, 127, 53, -87, 33, 3, -128, -93, 127, 127, 119, 127, 127, 43, -128, -11, 127, 116, -92, -63, -70, 119, 36, 18, -57, 57, 127, 127, 102, -34, -76, -64, 23, 29, 124, 127, -7, -18, -49, -97, -52, -71, -64, 1, 8, -103, 97, 127, 127, -98, -128, -16, 127, 116, -43, -128, -36, 0, -21, 17, 42, -121, -54, 127, 127, 36, -54, -128, -3, 127, 21, -70, -16, 49, 44, 127, 32, 33, -6, -50, 53, 81, 69, 70, 52, -127, -49, 1, 127, 127, 50, -32, 37, 127, 49, -87, -128, -128, -128, -102, 112, 127, 127, 91, 28, -128, -118, -17, 49, 50, 127, -128, -128, -128, -128, -128, 50, 116, 122, -13, -50, -128, -26, 1, -73, 8, 127, 101, -79, 21, -8, -128, -128, -128, -16, -76, -128, -103, 108, 114, -33, -32, 37, 88, 118, 127, 118, -128, -128, -76, 37, -21, 53, -45, -80, -128, -112, -95, -128, -118, 127, 123, -85, -128, -95, -16, -123, -13, 108, 127, 96, 38, -128, 10, 95, -68, -128, 29, 121, 13, -128, -128, -36, 21, 127, 127, 24, 33, 127, 127, 49, -128, -63, 127, 114, -114, -23, 39, 2, 39, 127, 127, 127, 7, -2, 127, 127, 127, 121, 80, 2, 59, 127, 127, 127, 121, -68, -128, -22, 96, -11, -128, -128, -128, -112, 122, 127, 127, -50, -59, -109, 29, 88, 127, 47, 5, -128, -128, -128, -8, -96, -26, -55, -24, -17, -24, -17, 31, 127, 5, -95, -128, -128, -37, 127, 127, -103, 12, 127, 127, 71, -113, -128, -26, 34, -108, -128, 18, 39, 108, -38, 47, -24, 127, -32, 55, 71, 54, -128, -128, -53, -128, -128, -44, 60, -63, -128, -38, -48, -3, 73, -2, -54, 97, 127, 86, -37, -111, -128, -93, 127, 127, 18, -128, -28, 111, 127, 65, -98, -128, 102, 127, 73, -128, -55, 1, -45, -90, 8, -7, 93, 3, -55, -78, -8, 24, -45, -18, -47, 127, 127, 58, -116, 28, 65, -128, -128, -128, -128, -39, 114, 127, 123, 88, 49, 13, 44, -108, -128, -128, -128, -128, -33, 3, -59, -128, -76, 113, 80, -128, -128, 91, 127, 22, -52, -128, -128, -128, 37, 74, -24, -128, -128, -128, -47, -18, -10, -38, -111, 38, 127, 127, -128, -128, -64, 85, 127, 127, 86, 37, 127, 127, -92, -128, -107, 79, 112, -2, -98, 119, 127, -128, -128, -49, -111, -128, -128, 60, 127, 118, -58, -78, -10, 127, 127, -128, -128, -128, -128, 13, 31, 43, 127, 127, 127, 127, 52, -128, -128, -3, 127, 127, 58, 45, -65, -128, -128, -1, 70, 43, -13, -7, 127, 127, -128, -93, 127, 66, -37, 28, 116, 23, 111, 66, 127, -36, -80, -128, -107, 22, 127, 127, -128, -128, -128, -10, 45, -12, -6, -12, 18, 33, -64, -128, 70, 54, -66, -60, 127, 127, -76, -66, -33, -55, -128, -100, -128, -64, 65, 127, 127, -88, -128, -128, 50, -58, -128, -128, -87, 127, 127, 127, 22, -128, -128, -128, -123, 73, 127, 127, 74, -65, -128, -121, -64, 52, 13, 109, -1, -21, -17, 127, 127, 127, -12, -128, -128, 8, 31, -92, -128, 11, 36, 70, 63, -5, 50, 76, 90, -55, 0, 127, -7, -76, -128, 53, 127, 127, 32, 10, -76, -128, -128, -128, 76, 127, 127, -38, -76, -81, -60, 86, 47, -16, 92, 87, 53, 7, 127, 22, -39, 69, 127, -16, -128, -128, -128, -63, 1, 90, 127, 53, -128, -128, -101, -111, 45, 127, -15, -75, 127, 127, 63, -128, -128, -68, -18, -113, -95, -47, 102, 66, -96, 0, 127, 81, 106, -112, -69, 23, 127, 117, -75, -128, -128, -128, -2, -15, -16, 76, 116, 127, 127, 37, -97, -17, 10, -93, -128, -29, 127, 127, -128, -23, 127, 127, 32, 53, 7, -128, -128, 103, 127, 127, -11, -128, -128, -57, 127, 127, -90, -128, -128, 127, 59, -52, -81, -38, -119, -65, 127, 127, 2, -128, -128, -69, -128, -128, 86, 127, 48, -108, 66, 127, -71, -71, 109, 127, 96, 7, 48, 116, 127, 80, -7, -23, -74, -121, 86, 100, 55, 119, 127, -76, -128, -128, 2, 127, 78, 36, -24, -70, -7, 80, -98, -96, 0, -128, -100, 93, 127, 127, 127, 71, 88, 127, -3, -128, -128, -128, -48, -103, -128, -128, -117, 21, 34, -64, -122, 15, -79, -122, -6, -57, -128, -128, -128, -128, -128, -23, 127, 127, -128, -128, -71, 127, 127, -64, -10, 0, -48, -28, 100, 80, 127, 127, -18, -117, 5, 127, 78, 0, 52, -16, 127, 127, 127, -80, -128, -128, 17, 2, 34, 36, 127, 127, 127, -13, -128, -70, 127, 127, 127, 127, 58, 6, 12, 76, 13, 127, 22, -58, -128, 78, 127, 66, -29, 0, 52, 127, 127, -42, -128, -117, -23, -68, -116, -128, 50, 127, 22, -128, -128, -128, 17, 127, 57, -1, 32, 44, 3, -42, -23, 57, -96, -38, 127, 21, -128, -43, 127, 127, 86, 111, -12, -69, 119, 88, -128, -128, -128, -128, -128, -91, -75, 2, 66, 87, -54, 11, -128, -128, -128, -70, -86, -128, -128, 31, 8, -78, -128, 28, 48, -34, -128, -128, 101, 16, 12, 15, 127, -128, -128, -128, -23, 121, 127, 80, 58, -44, -128, -128, 0, -3, -37, 68, 22, -65, -128, -128, -128, 127, 127, -8, -128, -32, 127, 127, 116, 100, 127, 127, -73, -128, -113, -85, -128, -128, 127, 127, 57, 93, 39, -42, -74, 39, -31, -33, -116, -128, -66, -128, -6, 7, 107, -103, -109, -65, 127, 127, 96, -70, -76, 29, 64, 127, -6, -107, -64, 74, -17, -128, -128, -102, 73, 127, 127, 127, -53, -90, -97, 53, 48, 24, -128, -76, -18, -29, 24, 57, 29, 127, 121, 73, -42, 21, 127, 127, -119, -128, 18, 127, 10, -128, -101, 78, 92, 59, 127, -39, -128, -38, 127, 127, -71, -128, -128, -7, 127, 113, -128, -128, -128, -113, -109, 127, 127, 11, -52, -23, -8, -107, 23, 10, -55, 107, 127, 127, 127, 127, 101, 0, -74, -102, -12, -92, 63, 1, 26, 8, -75, -27, 127, 127, 5, -128, -128, 127, 127, 73, -128, -128, -93, -57, 76, 92, -106, -103, -27, 127, 127, 5, 58, 127, 127, -21, -128, -128, -128, -22, -16, -65, -128, -74, 32, 57, 95, 127, 6, -128, -128, 123, 127, -65, -128, -128, -128, -78, -22, -45, -128, -24, -102, -109, -121, 118, 127, 127, 8, -63, -23, 127, 127, -21, -39, 76, 127, 21, -28, 100, 127, 127, 74, -12, -57, 127, 127, -16, -127, -128, -128, -70, 127, 127, 24, -128, -106, 53, -128, -128, -128, -128, -95, -68, -65, 42, -47, -66, -18, 10, -128, -128, 76, 127, 127, 127, 127, 63, 0, 127, 127, 127, 78, 39, -128, -128, -70, 119, 95, 11, -10, -69, -108, 49, -6, 109, -71, -128, -128, -58, 85, 24, -122, 2, 127, 127, 71, 127, -34, -128, -128, -98, 79, 127, 127, 22, 42, 58, -8, 21, 111, 127, 13, -21, -81, -18, -65, -22, 8, -38, -1, -21, 3, -122, -128, -128, -128, 93, 127, 97, -128, -128, -128, 111, 127, -21, -128, -128, -68, 116, 127, -1, -128, -128, 21, 123, 109, -128, -128, -79, 127, 69, -53, -128, -121, -80, 79, 113, -106, -128, -43, 63, 117, 127, 127, -33, -128, -88, 113, 127, 127, -38, -128, -128, 127, 96, 3, -50, 21, -74, 79, 127, 74, -128, -128, -5, 101, 127, -47, -11, 127, 127, 68, -128, -128, 109, 127, 73, -124, -42, 111, 127, 114, 127, 34, -128, -128, 71, 127, 55, -128, -128, -50, -17, -74, -54, 127, -63, -128, -70, 8, 31, 5, -32, -128, -128, -128, -128, 127, 127, -31, -128, -43, 86, 12, 50, 127, 95, -23, 65, 66, -64, -128, -118, 0, -128, -128, 27, 127, 121, 15, -36, -103, -108, -122, -76, -6, -128, -128, 27, -5, 66, 127, 127, -54, -128, -128, 73, -23, -96, 90, 127, 31, 58, 127, -48, -128, 39, 127, 112, 91, 76, -29, -128, -113, -128, -128, -128, -28, -15, 60, 127, 119, -79, -128, -128, 127, 23, -70, -128, 47, 127, 127, -97, -128, -107, 127, 127, -31, -128, -128, 6, 127, 127, 127, 78, 28, 97, 8, 42, 65, 127, 127, 127, -101, -117, 29, 127, 79, -12, 64, 127, 69, -5, -128, -128, -128, 91, 127, 127, -103, -118, -128, 55, 116, 127, 127, 127, 127, 127, -37, -70, -102, -45, 53, 127, 127, 103, 127, 65, -128, -128, -128, -128, -128, -128, 11, 127, 74, -128, -128, -27, 119, 11, -128, -128, 127, 127, 55, -106, -16, 54, 71, -8, -38, -50, -78, -128, -128, 2, 127, 127, 29, -16, 73, 48, -27, 31, -5, -6, 73, 127, 118, 38, -116, -43, -28, -87, -128, -128, -128, 24, 74, 58, 6, 32, 127, 127, 127, -128, -128, -95, 112, -32, -128, -128, 106, 98, 109, 71, 127, 127, -48, -128, -34, 127, 127, 122, -21, -128, -128, -27, 12, -37, 45, 66, 127, 37, -128, -128, -128, -128, -111, 87, 127, 127, 127, 16, -109, -95, -3, 47, 97, 92, 3, 107, 127, 32, -45, -128, -128, -128, -128, -128, 127, 127, 127, -38, -128, -69, 28, 87, 127, 98, -128, -128, -128, -18, 3, -127, -128, -73, 70, 127, 127, 24, -58, -128, -128, -12, 127, 127, 127, 76, -91, -128, -128, -96, 15, 69, 127, 127, -65, -128, -55, 127, 127, 75, 127, 6, -74, -81, -12, -38, -26, 127, -3, -121, -128, -7, 32, 27, -128, -128, -128, 5, 127, 127, 127, 6, 50, 127, 123, -36, -128, -128, -128, 2, 123, 127, -114, -107, 13, -102, -52, 103, 118, -12, 12, -128, -92, -52, 90, 127, 127, -54, -128, -22, 54, -128, -128, -70, 98, 127, 127, 87, -22, -33, 5, -50, 127, 123, 91, 127, 32, -128, -128, -38, 32, -1, 8, 127, -102, -128, -128, 43, 70, -124, -128, -32, 127, 127, -69, -92, 12, 127, 97, -73, -128, -98, -16, -37, -10, -32, 70, -128, -128, -90, 78, -128, -128, -128, 29, 123, 1, -73, 0, 10, -68, -16, 0, 8, -73, 28, 0, 64, -48, 95, -5, -44, -60, 127, -18, -128, -65, 127, 127, -128, -128, -34, 127, 0, 8, 119, -48, -63, 36, 52, -55, 127, 127, 11, -128, -95, 127, 127, 74, -24, -128, -128, -90, -5, 127, 119, 27, -1, 127, 127, 127, 127, 43, -128, -78, -2, 127, 127, 127, 116, 37, 92, 127, 108, -78, -124, -128, -3, -60, -128, -128, 73, 93, 103, 127, 127, -79, -128, -111, -28, -50, -54, -128, 88, 127, -128, -114, 127, 127, 127, 127, 45, -128, -128, -36, 2, -28, -118, -32, 127, 127, 127, 37, -128, -128, -128, -29, 59, 48, 107, 122, 100, -42, -96, -128, 78, 127, 97, -128, -128, -22, 43, -95, -128, -128, -128, 74, 127, 114, -3, 106, 127, -128, -128, -66, 127, 127, -13, 75, 127, 127, 33, -128, -128, -128, -128, -128, -128, -59, 127, 127, -7, -15, -128, -128, -128, -128, -128, -128, 11, -5, -24, -103, -1, -128, -97, -101, -15, 26, 58, -114, -128, -128, -31, 44, -49, -88, 88, 96, -128, -128, -128, -55, 29, -29, -101, 127, 127, 127, -64, -58, -8, -128, -15, 92, 49, -128, -74, 127, 127, -70, -128, 12, 127, 55, -88, -128, -65, -65, -128, 2, 55, 18, -106, -52, -86, -124, -98, -116, 8, 112, 17, -128, -128, -128, -128, -128, -109, -45, -71, -58, 15, 127, 127, -5, 37, 127, 127, -128, -128, -59, -128, -113, 21, 127, -21, -128, -108, 3, -128, -128, 27, 127, 127, -34, -38, 127, 127, 127, -81, -128, -26, 127, 127, 127, -59, -128, -107, 127, 127, -57, 11, 127, 127, 127, 71, -47, -128, -128, 22, 127, 127, -16, -101, -53, 90, -95, -128, -128, -42, -128, -128, 127, 127, 127, 17, 70, 119, 10, 18, -103, -128, -107, 78, 81, 5, -128, -97, -128, -81, -17, -93, -128, 48, 127, 106, 17, 127, 127, 1, 58, 127, 32, 44, -15, 73, -18, -43, -53, 34, -73, -128, -128, -128, -128, -128, -29, 127, 127, 15, -128, -128, -124, 127, 127, 127, 127, 127, 127, -47, -128, -73, 86, 42, -34, -15, 109, 79, 127, -88, -128, -128, 0, 100, 28, 12, 3, 127, 127, 37, -128, -128, -22, -58, -34, 127, 127, -113, -98, -7, -112, -128, -113, 3, 127, 127, 127, 127, -7, -128, -64, 127, 74, -128, -128, -128, 38, 81, -52, -128, -86, -13, 3, 78, 24, -95, 127, 127, -60, -47, 127, 127, 127, 127, 127, 112, 15, 8, 127, 127, -29, -128, -18, 127, 98, -43, 13, 127, 33, 31, -3, -44, -128, -109, -87, 127, 127, 127, -54, -128, -128, 116, 127, -7, -128, -128, -119, -11, 121, 127, 127, 97, 42, 33, 127, 127, -74, -128, -128, 127, 127, 91, -128, -112, 29, -124, -128, -59, 127, 18, -127, 127, 127, -73, -128, -128, 33, -8, -8, -88, 36, 50, 127, -128, -128, -128, 58, 127, 127, -15, -128, -128, 36, 127, 22, -114, -39, 55, -128, -106, 127, 117, -58, -128, -128, -128, -128, -75, 26, 55, -63, -128, -128, 8, 59, 127, 127, 22, -128, -127, 18, -128, -127, -34, -116, -128, 127, 127, 127, 92, 127, -44, -33, -29, 17, 127, 127, 101, -54, 26, 59, -103, -122, -68, 75, 73, -64, -128, -128, -27, 76, 11, -119, -34, 50, 113, 127, 21, -87, -128, -127, 7, -45, -6, 127, 48, -128, -66, 87, 123, -43, -6, 80, -128, -23, 127, 79, -17, 127, 88, -128, -128, -128, -34, 3, 106, 70, 17, -128, -128, 0, 127, 70, -119, -50, -73, 127, 127, 97, -85, -50, 11, -101, -85, -34, 127, 127, 124, -5, -65, 127, 127, 127, -80, 26, 98, -45, -114, 37, 22, -44, -47, 38, -128, -128, -128, 92, 127, 127, 8, -44, 8, 127, 127, 109, 127, -37, -27, 63, 127, -98, -128, -128, -75, 127, 127, 85, -33, 31, -15, -114, -128, -128, -78, 23, 26, -73, -128, -128, -114, -128, -92, -85, 33, 57, 127, 65, -63, -96, 37, 54, -106, 100, 127, 127, 78, -54, -128, -79, -33, -59, -111, -66, 121, 80, -18, 81, 127, 24, 127, 127, 127, -93, -128, -128, 97, 114, 116, 127, 127, 18, 85, 34, 15, 55, 22, -128, -101, -54, -128, -32, -128, -57, -57, 47, 22, 127, 127, 127, 122, 127, 54, 108, 76, 6, -113, -68, -128, -128, -2, 127, 127, -81, -29, 127, 86, -128, -128, -80, 127, 127, 17, -128, -6, 127, -88, -87, 64, 127, 87, 127, 112, 23, -128, -111, 18, 18, -71, -15, 127, 68, -128, -108, 68, 48, 32, -23, -128, -80, 13, -124, -128, 127, 127, 98, 127, 127, 127, 127, 60, 93, 65, 22, 18, -2, 34, 127, 127, -32, -15, -103, -128, 52, 127, 127, 127, -2, -128, -128, -128, -90, 113, 127, -15, -128, -34, 107, 37, -128, -128, 11, 127, 127, 127, 108, 121, -43, -128, 1, 127, 127, 127, 127, 127, 127, 127, 127, -23, -114, 22, 117, -55, -26, 127, 127, -85, -128, -73, 60, 45, -13, 103, 127, 127, -71, -64, 127, 127, 107, -128, -128, -55, 74, -58, 1, 12, 1, -79, 119, 127, 44, -18, 27, 85, -78, 11, 95, 127, 127, 70, -128, -128, 28, 127, 127, 127, 38, -128, -98, 127, 3, -128, -128, 80, 73, 17, -27, 127, 96, -28, -128, -87, 37, 127, 118, -103, -86, 12, 90, 63, 75, -81, -128, -128, 63, 127, 127, -11, -1, -128, -128, -128, 127, 127, 55, -128, -24, 66, 127, 59, -113, -128, -128, 127, 127, 96, 127, -58, -128, 10, 127, 127, -113, -128, -128, -128, -15, 121, -48, -116, -39, -128, -90, 127, 103, -128, -128, -123, 127, 127, 103, 18, -112, -75, -29, 127, 127, 127, -80, -128, -39, 116, -32, -86, 127, 127, 127, 124, -98, -128, -128, -63, -69, -102, -128, -59, 17, 127, 127, 127, -59, -128, 18, 127, 33, 71, 127, -42, -128, -128, -34, 103, 107, 6, -6, 127, 127, -71, -128, 24, 127, 127, 0, -101, -128, -128, 127, 127, 12, 8, 127, 127, -15, -17, -5, -128, -128, -128, -128, -128, -29, 71, -101, -128, -13, 81, -75, -42, 127, 127, -100, -102, 64, 127, 28, -128, -128, -127, 16, 127, 86, -128, -128, -128, -128, -97, 127, 95, -15, 11, -34, -128, -128, 2, 127, 127, 124, -22, 60, 52, 127, -17, -128, -90, 17, 28, -76, 127, 127, 127, 42, -29, -59, -128, -128, -128, -1, 127, 127, 127, 127, -102, -128, -128, -128, 15, 37, -101, -128, -128, -37, 127, 127, 127, -3, -128, -128, 69, 86, 127, 87, 42, -76, 71, 127, 127, 92, -76, 7, 106, 44, -33, 127, 127, -1, 70, 127, 27, 64, -11, -101, -128, -128, 73, 48, -76, -54, -109, -128, -128, -121, 22, 63, -13, -81, 37, 53, -128, -128, -128, -57, 102, 127, 93, -128, -60, 127, 127, 15, -128, -76, 37, -128, -128, -96, 117, 127, 85, -128, -128, -26, -32, 3, 113, 127, -128, -92, 66, 117, -66, -98, 123, 127, 64, -128, -128, 36, 127, 127, 127, 127, -34, -128, -57, 12, -75, -128, -127, -128, 0, 113, 127, 81, -108, -79, 3, 65, -16, 33, -28, -128, -128, -48, 7, 100, 127, 127, -54, -6, 2, -128, -128, 87, 127, 5, -128, -42, 127, 127, 127, 127, 127, 10, -49, -78, 78, 78, 103, -78, -123, 2, 127, 127, 127, 65, -7, -45, -15, 15, 11, -11, -128, -87, 121, 55, -85, -128, -78, 100, 127, 127, 68, 121, 127, 127, 114, -128, -128, 48, 123, -128, -128, -117, -58, -128, -128, -128, -79, -123, -66, 24, -29, -58, 118, 127, 108, -79, -73, -24, 0, 58, 109, 8, -26, -76, 42, 119, -2, -128, -128, -92, 11, 127, 127, 127, 10, -98, -128, -128, -108, -23, 47, 111, 2, -128, -128, -128, -47, 18, 37, 112, 127, 127, -11, -1, 53, -15, -69, -57, -128, -128, -49, -29, -128, -79, 91, -87, -128, -38, 6, 0, -48, -128, -128, 97, 32, -101, -128, -116, -128, -88, -128, -107, -54, -60, -128, -128, -128, 79, 39, -103, -128, -71, 127, 127, 127, 127, 112, -87, -128, 6, 127, 107, 36, 0, -29, -98, -7, 112, 118, -79, -128, -6, 127, -7, -111, 17, 102, 81, -13, -123, -128, -128, -128, 10, 65, -26, -128, 0, 32, 15, -128, -128, -64, -49, -36, -121, -97, -128, -97, 127, 127, 5, -128, -128, 108, 127, 96, -2, -32, -53, 118, 52, -102, -127, -5, 127, 127, 2, -33, 0, -66, 2, -128, -97, 109, 65, 33, 122, 127, -68, 90, 127, -5, -128, -128, 54, 127, 38, -34, 127, 127, 127, 127, 87, -71, -128, -58, -128, -128, 24, 127 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
