-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
            18, -8, -8, 4, 14, -9, -14, 20, -15, 16, 9, -2, -3, -12     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -4, -23, 70, 97, -125, -115, 123, -86, -83, -65, 28, 89, -22, 29, 65, -105, -18, -124, 98, 24, -37, 84, -37, -12, -125, 6, 16, 107, 117, -77, -22, -83, 30, 112, -96, -95, 52, 36, -53, -113, 31, -62, 67, 88, 78, 18, 25, 83, 50, 55, 24, 112, -75, -35, 72, 56, -120, -122, 2, -25, -3, -127, -114, -115, -123, 26, -11, 91, -7, 53, 94, 45, -118, -36, 17, 17, 81, -49, 26, -58, -3, -2, -69, -92, -40, -70, 67, -96, -6, -115, 116, -80, 111, 41, 42, -71, -114, -76, -124, -62, 27, 72, -98, -42, -33, -52, 42, -74, 36, -68, 112, 93, 110, -63, 110, -128, -121, 108, -32, -21, 95, 50, -21, -36, -16, -49, 93, 91, -9, -45, -48, 43, -88, 73, -105, -126, -62, 44, 41, -45, -6, 93, 40, 56, -42, 121, 109, -103, -103, 103, -48, 95, 83, -37, 31, -33, -20, 127, -112, 86, -122, -26, -71, 127, -4, -70, -115, 113, -69, 84, 23, 27, -1, 10, 103, 43, 91, 48, 46, 109, 94, -78, -102, 73, 15, -4, 84, 18, -13, -84, -126, 23, 4, -105, -101, -53, -46, 8, -91, 79, -90, -97, -49, 120, 8, 46, 120, 70, 8, 79, -101, -28, 14, -105, 31, 57, 45, 90, 68, -47, -20, 59, -55, 47, 18, -3, -123, 16, 42, 53, 116, -103, -18, 108, 107, -35, 47, -16, -68, 94, 112, -39, 85, -9, 74, 103, -19, -127, -20, 30, -3, -58, 117, 69, -92, 47, -25, 65, 49, 9, -39, -41, 78, 99, -62, 84, -86, 84, -34, 106, 40, -4, 30, -96, 87, 56, -4, -37, 8, -119, -113, 37, 53, -13, -88, 88, -58, -34, 113, -79, -100, -52, -82, -23, 97, 65, -30, 84, 7, -117, 60, 124, 122, 120, 105, 55, -105, -30, 72, -13, 41, -101, -96, 126, 104, -57, 108, -96, -97, -87, 22, 29, -21, 110, -32, -109, 1, -9, 31, -72, 21, 74, 74, 107, 26, -90, -50, -8, 118, -113, 98, 17, -60, 114, 60, 97, 100, -44, -17, -75, 122, -38, -6, 13, 77, 106, 8, -77, -94, -57, 2, 9, 16, -18, -63, -78, -3, 110, -4, -30, -75, 91, 54, -31, -57, 4, 117, -76, 86, -44, 80, 46, 79, -68, 68, 17, 64, -124, 85, -90, 60, 103, -117, -33, -17, 91, 85, -60, -19, -92, -68, 108, 13, -109, 97, -107, 72, 104, 51, -48, -4, -112, 36, 0, -77, -52, 118, -57, 90, -68, -44, -80, -114, -65, -61, -82, 95, 109, 85, 62, 65, 21, -18, -7, 60, -39, -54, -43, 74, 105, -36, -96, 39, -81, -63, 82, -85, -90, -43, 108, -31, 96, -80, 113, 96, 18, -76, -13, -90, -58, 20, 91, -6, -44, 82, -66, 114, 116, 118, 97, -108, 35, 45, -33, -58, 70, 6, -68, 7, -23, 121, 112, 11, -121, -125, 67, 26, -12, -59, 121, 91, 0, -38, 64, -94, -126, -39, -64, 104, 28, 109, 4, 68, -18, -99, 56, -26, 47, -45, 126, 119, 65, -25, 71, 32, -113, -32, 55, -103, 48, 14, 4, -66, -22, 103, 60, -46, 6, 52, 41, 82, -4, 88, 64, -53, 21, 111, 64, 118, -45, -70, 37, -112, -38, 102, 95, 82, -114, -42, 3, -38, 3, -123, -53, -58, 80, 39, -73, -30, 72, 65, -12, 32, 126, -3, 31, 76, -120, 85, -63, 104, 26, -18, -112, -38, 75, 84, -63, -125, -87, -78, 8, 94, 66, -27, 122, -84, 84, 25, -3, 36, -51, 26, 1, 53, 113, -2, 25, 121, -21, -88, -61, 51, 20, 63, 10, 97, -96, -23, 58, -30, -103, 2, 87, 85, -37, 125, 59, -12, 74, 76, 105, -80, 126, -124, -9, 66, 29, -5, -27, -60, 46, 2, 67, 27, 32, -33, -117, -101, 1, 82, 29, -78, -116, -54, 3, -124, -104, -89, 49, -98, 58, -38, -97, -67, 30, -67, -2, 45, 61, 82, -3, 67, -19, 74, -27, 94, 107, -15, -70, 71, -79, 48, 5, -128, 69, -22, 116, 88, -45, -80, -58, 123, 100, 28, -95, 46, -41, 3, 16, -124, -94, 35, 115, -122, 5, -127, -122, -13, -120, 97, -92, 93, -89, -120, 10, -102, -22, 85, -67, 61, -126, -70, -98, -49, 3, 72, 67, 111, -42, 72, -122, -124, 8, -107, -109, 99, 5, 53, 74, -85, 8, -94, -49, -120, 53, -16, 85, -96, -62, 88, 54, 72, -20, -127, 97, 28, 9, -16, 44, 32, -89, -24, -19, -61, 14, 61, 51, 52, -87, 62, -117, 2, 62, -105, 0, 64, -84, 55, 6, 120, 73, -6, -122, 124, -128, -7, -16, -9, -41, 1, -35, 84, 44, -126, -93, 77, 16, 29, 99, 16, -113, 52, 49, -62, 7, -14, 85, -15, 42, -79, -50, 87, 49, 96, 46, 89, -86, 87, -99, -126, 69, -1, 29, -7, 95, -2, 50, 82, -55, 24, 93, -77, -11, -21, -34, 98, -106, -53, 100, 121, 50, 33, 111, -110, -91, 101, 17, 64, 27, 25, -15, 41, -10, -47, -52, 83, -103, 84, 106, -61, 47, 111, 70, -31, -98, -50, -116, 29, 73, 43, -48, 92, 118, -42, -69, 86, 110, -88, -10, 7, -100, -95, 83, 71, -23, -78, -90, -72, 12, -14, -79, 121, 79, -90, 31, -18, -52, 61, -92, -106, 82, -84, -25, -44, -17, -21, -64, 108, 59, 65, -118, -97, 111, -59, 22, -18, -20, -13, -51, 113, -61, -24, -66, -94, -91, 33, -73, 5, -53, 5, 7, 20, -121, -81, 20, -128, -117, -99, 24, 112, -89, -100, -127, -89, 90, 14, -59, 74, -60, -77, -128, -88, -67, 68, 68, -44, -89, -20, 58, -40, -72, 127, -112, 35, -8, 15, 28, -119, -112, -102, 73, -96, -32, 79, 81, -61, -81, -52, 106, -104, -128, 11, 110, 88, 111, -22, 107, 121, 67, 5, -52, 32, -115, -2, -82, -118, 46, -123, 50, -88, 127, -42, 45, 68, -54, -104, -102, -5, 10, -62, 101, -79, 117, 67, 10, -5, -75, 76, 54, -55, -43, 113, -128, 33, 66, -102, -52, -30, 109, 82, -21, -55, -99, -37, -15, -110, -88, 77, -69, 87, -126, 51, 76, -104, 33, 91, -29, 78, -47, -42, 91, -109, -98, 72, -126, 37, -120, -110, 62, -61, 62, -1, -110, 78, -11, 82, 121, -27, 27, -21, 81, -78, 120, -37, 89, 22, -97, 92, 24, -110, 15, -41, -97, -9, -23, -78, 75, -128, 73, 81, -120, 104, 89, -40, 93, 116, -118, -11, -128, -38, 100, -126, -103, -10, -60, -42, -11, -28, -46, -104, -46, 74, 91, -92, 17, -111, -92, -71, 127, -109, 57, -35, -23, 67, 37, 126, -70, -84, 47, -95, -18, -53, -69, 105, 102, -73, -42, -91, 81, 97, -74, 17, -98, -53, 112, -90, 29, -126, -47, -28, 68, -73, 8, 43, -66, -116, -116, -110, -14, -114, 12, 9, 84, 7, -121, 62, -64, -23, 109, 25, 1, 99, 17, -35, -6, 12, -45, -82, -89, 55, -3, -32, 103, -72, -125, 55, -8, 94, 56, -122, -98, -118, -92, -112, -3, -47, 119, 34, 90, -123, -50, -5, 53, 97, 30, -66, -38, -44, 2, 88, 12, -97, -62, 4, 109, 53, 40, 127, 36, -2, -83, 115, -14, 42, 46, 106, 39, -120, -27, -74, 126, -82, -71, 124, -9, 98, -5, 85, 27, -69, -43, -57, 98, 89, 9, 87, 60, -79, 30, -48, 55, -66, -67, -77, 79, 70, 29, -22, 38, 23, -127, 23, 63, -28, 12, 51, -36, 23, -41, 123, 13, 116, -108, 109, 76, 15, -125, -94, 34, -12, -63, -48, -85, -77, 22, 27, 20, -90, 2, -108, 116, -106, -28, 66, 51, -55, -75, -101, -76, 73, -114, -56, -65, 38, 93, 58, -37, -103, -82, -72, 5, -18, -83, 127, 35, 6, 101, -36, -48, -44, 69, 90, -2, 52, 115, -2, 24, -112, -97, -74, 96, 116, -72, 82, 103, -32, 17, -64, 91, 120, 84, 66, -122, 8, -9, -96, -128, -109, 34, 69, -30, 50, -89, 43, -35, 45, -107, -120, 105, 87, -39, 75, 95, -122, -79, 43, -20, 112, -18, -124, 28, -100, -105, 88, 1, -26, 72, -17, -71, 45, 126, 40, 47, 97, -79, -8, -88, 12, 70, 20, 26, 88, -56, 118, -10, 68, -40, -63, -59, -49, -52, -75, -49, 64, -60, 77, 104, -49, -4, -118, 61, -120, 96, -51, -30, -7, 62, 30, 86, -66, 44, 70, 8, -51, 74, 9, 90, -107, -7, -115, 118, 27, -27, 79, 112, -38, 118, -73, 76, -28, -24, -63, -24, -70, 99, 102, -100, 114, 122, -90, -88, 127, -92, 17, 52, 62, 42, -7, 45, -41, -95, 118, -127, 94, -15, 73, 84, -118, -55, 78, 74, -76, -35, -17, -80, -4, -18, -22, 31, 41, 23, -48, -72, -110, 112, -32, -27, 36, 23, -25, 73, 117, -117, -55, 13, 0, 98, -40, 99, 120, -11, 36, 72, -17, -90, -86, -86, 99, -20, 36, -103, 65, 16, -28, -64, -85, 59, 6, -61, 84, 71, -107, 70, 57, 95, -126, 82, 68, 64, 50, 20, 124, 98, 63, -67, 75, -5, -23, -102, 18, -44, -60, 72, -78, 104, 107, -15, -82, 82, -126, -16, 93, 121, -63, -116, 4, -37, -83, 47, -44, 103, -67, -63, 3, -15, -59, 101, -91, -63, -79, -39, -3, -70, -116, 125, 107, 122, 99, 4, 107, -106, 0, 29, 25, -56, 21, 21, 77, -65, -90, 75, -123, -25, -59, 14, 5, 37, 24, -41, 19, 25, -89, -21, -41, 99, -60, -96, 66, 87, 1, 51, 9, -35, 1, -55, 55, 6, -15, 0, -81, 126, 109, -84, 115, 24, 62, 62, 1, -41, 106, 1, -85, 95, 64, -127, 31, 108, -70, 78, -36, -4, -51, -11, -39, -82, 51, -13, -125, -47, 124, 75, 4, 16, 21, 49, 72, 112, -101, 101, 33, -15, -96, -121, -109, -97, -123, -17, 102, 64, 19, 54, -22, -105, 37, 70, -62, 24, 30, 103, 32, -29, 59, 101, 12, 127, -54, -103, -123, -111, 91, 50, -100, -108, 34, 10, -44, -8, -61, -31, -80, -109, -59, -48, 84, -128, 70, -101, -61, -48, -86, 99, -23, -17, 20, 125, 113, 74, 18, -14, -100, -86, 72, 19, 99, 63, -33, -34, -6, 81, -31, 54, 105, -32, 97, 15, 102, 4, -95, -87, 2, 83, -9, 2, 35, 44, -128, 29, -42, 105, -61, -19, -17, -52, 95, -43, 27, 33, -16, 109, -87, -45, 42, 116, -37, 51, -36, -118, -70, 84, 40, -115, 87, 51, -27, -40, -92, 25, 77, -70, 67, 127, 10, -93, -83, 74, 46, -98, 53, 98, 54, 37, -101, 82, -49, 121, 101, -30, -14, 59, -105, -39, 63, 3, -87, -117, -14, 91, -37, 118, -51, 81, -110, 4, -102, -82, -102, 90, -4, -54, 86, -115, 74, -24, 116, -89, -104, 7, 12, 80, -22, 59, -33, 66, 10, 122, -29, 73, -124, -4, 33, -17, -17, -12, -69, -110, -19, 36, 20, 37, -103, -112, -25, 13, -30, 91, -78, 91, -7, -51, 15, -25, 31, -77, 84, -107, -119, -43, 17, -23, -25, -30, 118, -54, -82, -5, 59, 36, 91, 84, -31, 1, 98, -93, 74, 112, 86, -97, 84, -14, -127, -68, -19, -17, -20, 2, 5, -28, 127, 36, 79, 18, 110, -124, 51, 116, -10, 10, -99, -4, 6, -2, 46, 15, -76, -54, 37, -119, -28, 50, -59, -16, 121, 21, 11, -101, 89, -25, 56, -57, 48, 109, -117, -27, -121, -50, 16, -127, 100, 59, -78, 80, 96, 17, -88, 36, -92, 84, 17, 76, 47, 53, -1, 41, -38, 83, -29, 18, 80, 90, 48, -4, -64, -41, 48, -58, 15, -10, 21, 69, 41, -47, 66, 14, 16, 107, 57, 119, 93, 1, -23, 15, 115, -97, 22, -59, 65, -55, 13, -82, 56, -68, 99, 33, 82, -62, -90, 11, -97, -43, -73, 26, 53, -31, 72, -35, -1, 119, -85, 125, 16, 121, 116, -118, 52, -27, -108, 101, 7, -83, 40, -97, 58, 42, 53, 30, -104, 93, 63, 34, 17, 127, -49, 77, -126, -76, -27, -87, -38, 104, -51, -56, 19, 30, 115, -46, -57, -80, 3, 57, -33, 69, 89, -54, 66, -98, 76, -31, 102, -60, 79, 55, -72, 112, -82, 26, -30, 0, 103, 44, -16, -11, -77, 94, -120, 28, 3, -80, -77, -94, -68, -121, 117, -118, -31, -49, -9, 57, -127, 89, 70, 47, -89, -104, 85, -42, 28, 5, -28, 35, -76, 93, -7, -96, 25, -86, -37, 121, 78, -1, 19, -38, -40, -120, 77, 104, 124, 92, 22, -38, 118, -85, -16, 70, -43, -83, 112, 75, -8, 15, 19, -47, 46, 84, -114, -22, -34, -101, 19, -124, 76, 47, 102, -115, 65, -114, -110, -62, -82, -70, -112, -96, 100, 10, 88, 10, -108, -87, 96, 92, 0, -16, -28, -47, -122, 63, -67, 35, 77, 56, -44, 19, -61, -15, 78, -14, -103, 48, 37, -7, 105, -64, 27, 54, 47, 116, 109, -88, -10, 77, -125, -77, -19, -122, -14, 94, -60, -20, 120, 69, -64, -86, 23, -98, 108, -121, 100, 103, 46, 64, 18, 90, -30, -95, 51, 101, 98, 62, 54, -6, -14, 10, -31, -66, 65, 82, -79, -83, -68, -49, -119, 48, -17, -56, -19, 7, -123, -35, -35, 65, -39, 24, 21, 61, 125, -11, -3, 42, -127, -114, -44, 86, 37, 1, -119, 56, -53, 54, -24, 25, 17, -5, -127, 2, 79, -67, -103, 84, 26, -85, 74, 64, 110, -23, 51, 9, -12, -100, -70, -1, 94, -43, 74, 6, -128, 12, 14, 113, -19, -61, -116, 121, -53, 73, 74, -108, 99, 99, 36, 16, -2, -48, 80, -37, 124, 3, 33, -24, 35, 31, 62, -94, 5, -34, 86, -74, 1, -87, -116, 63, 68, 86, -126, 78, 115, 80, 68, 1, 58, 40, -73, -62, -96, 6, -27, -91, 124, -39, -126, -110, -23, -108, 50, -83, -91, 27, -75, 69, 13, -105, -49, 109, -79, 119, 117, -66, -65, -77, -68, 17, -82, 8, 118, 38, -12, -47, -120, 91, 47, 114, 111, 125, -21, 89, -24, 21, 80, 81, -102, -123, -78, 37, 82, -39, 79, -127, 105, -110, 30, 119, -10, 91, -45, 8, 104, -46, -107, -2, -82, -24, 119, -53, 94, 38, -2, -40, -23, 40, -107, 39, -113, 85, -99, 121, 16, 72, -69, 10, -36, -117, 0, -23, 69, 36, -51, -45, 61, -23, 43, -62, -1, -19, -7, 126, 29, 109, -45, 89, 60, -121, -1, 14, 95, -63, -67, -25, 41, 23, -40, -33, -22, -51, -16, -66, 64, 92, -106, -72, -50, -47, -107, -113, -97, -59, -38, -105, 47, 23, -14, 104, 31, -76, -8, 115, 5, -114, -14, -64, -13, -57, -101, -63, -116, -29, -17, -2, 112, -46, -15, 44, -19, -64, 77, -19, -32, -127, 102, 13, -105, -122, -92, 21, 107, 72, 21, 125, 10, -93, 82, 104, 13, -33, -25, 68, -121, 124, -21, -79, -116, 3, -15, 87, -87, -11, -6, 90, 80, -23, 119, -23, 70, -101, -31, -35, -103, -113, -7, -50, 13, -111, -89, 65, 83, 99, 56, -86, 39, -46, -20, 105, 113, 102, -9, 73, 88, 54, 62, 29, 63, -27, -9, -128, 90, -120, 97, 3, 57, 47, -9, 58, -79, 26, -20, 47, -99, -55, -55, -94, -123, 9, -11, -101, -100, 100, 120, -116, -59, -128, 50, 115, 114, -100, 37, 83, 6, 87, -8, -122, 70, 103, -120, -54, 24, -40, 80, -89, -65, -44, 54, 108, 29, 85, -45, 25, -4, 59, -56, -40, -59, 22, -102, -121, -21, -76, -115, -109, -11, -55, 11, -28, 40, 120, 2, 16, -5, 38, 63, -124, -114, -102, -99, 16, -3, 31, 77, 110, -31, -109, 97, -35, 48, -123, 62, 52, -35, -48, 33, -67, -113, -115, -50, -86, 111, 21, -4, -32, -53, -103, 68, 37, 11, 31, -57, -119, -77, 103, -111, 13, -106, -31, 32, -18, 49, -6, -125, -7, 60, 115, -27, 28, 42, 101, -18, -83, -70, -57, -68, 77, -25, -68, -112, 88, -86, -54, 127, -77, 72, -76, 89, -94, -111, -33, 35, 87, -30, -96, -44, 48, -35, -86, -115, -80, 14, 55, 12, -81, 80, 98, -91, -80, -47, -21, -118, -50, -117, -90, 107, -80, -24, -39, 11, -30, 109, 92, 95, 15, 112, -106, -40, 111, -40, -69, 104, 46, -60, -28, 105, 16, -110, 20, 11, -7, -30, -113, -120, 83, -102, -34, 67, -44, -91, 107, 92, -98, 46, 23, -22, 30, 36, -4, 82, -107, 78, -128, -98, -90, 70, 41, -28, -128, 104, 106, 40, 69, 46, 49, -122, 115, -94, 11, -86, -91, -13, 31, -116, 38, 47, -122, 11, -21, 74, -14, -89, -104, 108, 49, -79, -28, -58, -119, -38, 117, 53, -12, 25, 29, -122, -72, -69, -62, -69, -38, -125, 97, 54, -37, 36, 43, -53, -106, -102, -101, -51, -111, 26, -19, -31, 87, -126, -128, 18, 101, -2, -122, 118, 1, -25, 47, -108, -53, 118, 42, -8, 62, -34, -12, 40, 105, -93, 53, -117, 10, 47, -128, 120, 66, 36, 72, -112, 19, 94, 74, 121, -80, 38, 126, 120, -48, -126, -97, -32, 125, -124, 73, 121, 79, -109, -90, -111, 10, 78, -49, 24, -61, 12, -6, 82, -121, 127, -39, -80, -46, -127, 97, -12, -8, 51, -2, 36, -113, -115, 58, -104, -52, 2, -53, -67, 24, -18, -122, -105, -109, 111, 64, -45, 18, -72, -74, -68, -96, -1, 95, 43, 24, -68, -40, 24, 110, -32, -124, -49, -86, -8, 97, -124, -86, -45, -31, -125, -78, -95, -59, 61, -99, -86, -101, 89, 46, -50, 96, 45, 36, 62, 66, -101, -21, 3, 3, 92, 20, -64, -92, -32, -118, -55, -115, -56, 95, 49, -121, -58, 24, 16, 126, 122, -85, -46, -124, 21, 25, -56, 15, -126, 43, 113, 51, 69, 15, 75, -90, 24, -78, 121, 94, 97, 63, 98, 119, 42, 93, -61, -106, -80, 88, 83, 123, -57, -111, 53, -67, -87, -122, -117, 97, 118, 114, -2, -24, -114, 46, 126, -26, 8, -57, -112, -9, -114, -95, -48, 94, 38, 15, -2, 57, 66, -3, -16, -69, 42, -101, 82, -119, 71, -28, 34, -91, -109, 4, -111, -38, -64, -123, -108, 27, 71, -22, -57, -118, -11, -73, 127, -9, -87, -85, -54, 22, -20, 82, -94, -121, 5, -97, -46, 127, -59, -52, -4, -33, 85, -3, -106, -64, -105, -90, 0, -105, -58, -110, 124, -114, 102, 92, 59, -18, -121, -113, 12, 96, -47, -9, 28, -69, 88, 120, -109, 28, 83, 89, 31, -96, 116, -7, -107, 108, -37, -22, 74, -82, 9, 124, 52, -1, -26, -99, -118, 22, 108, 66, -61, -99, 47, -61, 104, -24, 53, -11, -63, -41, 90, 76, 22, -107, -12, -59, -61, -92, 117, 125, 48, 95, 9, -95, 123, -101, -28, -109, -31, 116, 11, -47, -108, -7, 50, -79, -69, -6, 57, 127, -11, 2, 62, 0, 73, 52, -86, 4, 108, -109, 25, -93, -5, 63, 49, -89, -47, -72, -127, -46, 56, -62, 76, 25, 92, -28, -118, -83, -27, 35, 20, 107, -47, -57, 94, -111, -100, 74, -68, 105, 33, 7, 17, -83, 75, -20, -77, 50, -6, -28, 77, 51, 97, -70, -119, 102, 73, 90, -46, 63, -114, -2, -17, -61, -29, -79, 81, 15, 10, -7, -59, -110, 0, -60, 49, -119, 74, -33, -94, 21, 106, 95, 118, -108, -101, 96, 75, -104, -52, -106, 108, -51, -118, 33, 2, 56, -27, -62, -67, -46, 87, 118, 115, 109, -74, -123, -100, 111, -109, -36, -98, -66, 54, -88, -108, 82, 120, 29, 46, -17, -32, -54, -94, -13, 43, -3, 38, 47, -74, -67, 96, 94, 22, -10, 124, 31, -99, -84, 35, -126, -14, -14, 97, 81, 109, 22, 12, -128, 126, -90, -7, -80, 79, 22, -112, -110, 19, 125, 29, 55, -75, -108, -88, -69, -12, -115, -59, -97, 126, 46, -17, 101, 109, -125, 123, -44, -116, -38, 41, -93, 4, 115, -64, 127, -60, 95, -125, 59, -53, 41, -115, 3, -15, 94, -53, -61, -91, 66, -13, 97, -79, -30, 62, 115, 72, -7, -50, -36, -93, 13, 47, 47, -109, -97, 11, -88, 73, -62, 0, -51, 16, -65, 121, -100, -106, -22, -115, -14, -18, 39, 110, -96, -15, -87, -105, 70, 100, 121, 3, 111, -105, 96, 51, -81, 27, -65, -105, 121, 57, 127, 51, -74, 14, 28, 74, -123, -67, -69, -126, -56, 30, -69, -45, -73, -33, 123, 89, -51, -47, 22, -62, 6, 94, -58, 51, -43, -72, -73, -108, 77, 54, -112, 76, 22, 125, 15, 94, -112, 45, 16, -100, 49, 101, -7, -15, 94, 124, -37, 79, -87, -72, -66, -10, -52, -92, -90, -20, 9, -124, 100, 100, -105, -13, 2, -49, 62, -100, 56, 127, -88, -92, 29, -86, 92, 10, 113, 127, -65, -95, 124, 103, -87, 62, 107, 50, -114, 3, -37, 80, -53, 30, -81, 123, 11, 78, 12, -101, -13, 90, 29, 56, -29, 94, 19, 61, 124, 4, 89, 42, 61, -51, 95, 37, -81, -22, 27, -68, -81, -125, 16, 37, 31, -49, 42, 110, -65, 54, 111, -62, -93, 2, 59, 11, -20, 78, 65, 126, -123, -15, -103, -65, -57, 71, 76, -48, -77, 126, 98, 2, -115, 1, 53, 84, 90, 121, -23, 74, 115, -78, -67, 21, 10, 115, 89, -20, -12, 51, 29, -6, 73, -1, -71, 88, -64, -125, 4, -92, -6, 55, 121, 115, 119, 102, 126, 30, 101, -113, -76, -85, 63, -96, -51, 110, -61, -108, -51, 97, -36, 88, 12, -103, 100, 9, -126, -67, 62, 42, 117, 47, -74, -110, 62, 98, -28, -111, -28, -102, -81, 84, -14, -87, 4, 47, -47, -71, -27, -115, -40, 68, 63, -114, 123, 33, 6, 83, -118, 81, -122, -105, 96, 60, 119, 19, 66, 90, 121, 102, 118, -65, -104, 80, 35, -68, -81, -31, -24, -81, 42, 83, -85, -115, -20, -60, 78, 80, 57, -67, -124, -107, 39, 27, -29, -85, 59, 65, 42, -23, -103, -4, 93, -128, 10, -4, -91, -77, -14, -109, -71, -49, -8, -107, 82, 95, 109, 4, -56, 74, 28, -93, -46, 12, -49, -39, -91, 48, -62, 77, -79, 46, 46, 101, -5, 84, -5, -108, -34, -98, -82, 19, 74, -102, 24, -77, -20, -47, 9, 96, -112, 113, -104, 121, 15, 26, 16, -113, -43, 106, -37, -103, -105, -33, -10, -124, 97, -108, -51, -81, 46, 37, -82, 13, 120, 99, 45, 86, 74, 36, 87, 103, 7, 40, 35, -8, -117, -25, 47, -116, -37, 60, -98, 93, -15, 63, 106, 83, -42, 50, -117, -117, 98, 70, -90, 62, -118, -17, 0, 106, 91, -6, -13, 24, 73, -41, -118, 29, 82, -43, 78, -10, 113, -116, 121, 88, -96, 23, 119, 7, -111, 21, 100, 121, 64, 107, -117, 17, -87, 5, -22, 102, 80, -121, -77, 39, -56, 43, -46, -124, 90, -2, -4, -73, 32, 23, -34, 11, -2, 71, -66, -1, -79, 11, 60, 77, -94, 122, 113, -44, 17, -95, -106, 2, -111, -12, 127, -18, -80, 18, -6, -109, -33, 20, 54, -22, 36, -3, 11, 74, 84, 81, 66, 81, -124, 61, -125, 97, 102, -97, -63, 11, 98, 127, -87, -14, -46, -43, 67, 78, -56, 38, -26, 9, -115, -1, -70, 89, 103, 74, -20, -67, -17, 5, -6, 87, 80, -24, 52, -51, -3, 36, 111, 76, -40, -47, -103, 43, -34, -117, -74, 46, -97, -22, 70, 81, 44, -77, 81, 94, -63, 43, 65, -63, -17, 92, -128, -25, -8, -21, 25, -74, 105, -102, -81, 22, -119, 107, -56, -5, -49, 79, -74, -99, 68, -119, -48, 81, -112, 119, 62, -124, 93, -19, 69, -26, -24, -128, 91, -57, 92, -63, 74, -116, -116, 15, 47, -77, 72, 48, 118, -68, -122, 68, -63, 57, 18, 74, 11, 58, -80, -47, -51, -50, -79, 46, 6, -24, 99, -56, -1, 102, 22, -107, 14, -80, -114, 18, -81, -4, 27, -46, -18, 31, -100, 60, -2, -85, 101, -97, 84, -74, -112, 42, 113, -25, -47, -22, 60, 26, -73, -29, 84, 61, 41, -80, 84, 22, 64, -32, -6, 74, -91, 121, -101, -91, -102, 64, -28, -43, 120, 20, -61, -20, -82, -19, 115, -122, 20, 90, 88, 125, 95, -90, -67, -29, -37, 80, 34, -28, -36, 113, -37, -57, 58, -75, -27, 38, -79, 52, 104, -4, -94, -22, 41, -8, -59, -22, -107, 0, 54, -42, -32, 59, 10, -6, -121, 15, -63, 81, 18, -19, -118, 121, -44, -93, -27, -124, 112, 69, 2, -27, -38, -15, -48, 56, -120, -53, 37, -59, 90, -38, 34, -19, 86, 75, -112, -43, -39, -125, 37, -86, -105, 53, 72, 118, 69, 14, -53, -115, 38, -79, -24, -85, -16, 99, 75, 36, -92, 40, -115, -114, 64, -55, 88, 9, 93, 101, -95, -98, -54, 122, 9, 95, 112, -80, 111, -128, -102, 62, 78, -2, -57, 85, -121, -7, -97, -58, 29, -5, -93, 122, -57, 16, -44, -87, 40, 103, -76, 9, 51, 95, 98, 98, 48, 83, 11, -124, 42, -52, -16, -77, 52, 20, -25, 10, -16, -6, -36, -74, -100, -91, -89, 22, -95, 70, 49, -79, 89, 111, -61, -23, -45, -73, 21, -70, -40, 28, 31, 118, 57, 96, 121, 15, -38, -56, -91, 73, 57, 4, 36, 78, -115, 46, 74, 44, -21, -19, 105, 50, -31, -107, -78, -106, 67, -32, 79, 15, 36, -114, -64, -109, 118, 107, 101, 126, 103, 86, -36, -71, -4, 105, -18, 95, 22, -6, -38, 122, 53, 5, -106, 120, -89, -97, -48, 89, 64, 123, -77, 102, -42, -113, 113, -77, 42, 125, -9, -30, -2, 3, 44, -14, 77, 30, -114, 103, -27, 80, 6, -72, -101, 117, 81, 22, -115, 76, 126, 102, -89, 2, -28, -77, 90, -107, -54, -44, 24, 0, 33, 110, 59, 89, 50, 25, 36, -127, 123, -117, 38, 83, 17, -110, -57, 57, 23, 20, -64, 56, -62, 40, -123, -83, -124, 6, -16, 46, -24, 15, -44, -70, 63, -5, 31, -40, -19, 109, -36, -90, -64, -44, -70, 107, -71, 105, -93, 119, -25, 122, -127, -37, 81, 17, 47, -81, 5, 114, 73, -50, -45, 10, 70, -114, -128, -83, -46, -46, -67, -55, 101, 46, 62, 127, 86, 11, -112, 49, 101, -125, 11, 99, 99, 19, -123, -9, 36, -78, 42, 15, 103, -111, -41, 42, 18, 125, 91, -128, 104, 31, -8, -56, -50, -40, 44, -21, 86, -27, 86, -99, 90, -93, 117, -60, -59, 25, 77, -6, 4, 45, 38, 105, 29, 15, 86, 57, -82, -94, 105, -51, 38, -27, 43, -13, 125, 55, 7, -97, -104, -32, 114, 23, 78, 88, 26, 21, -7, 81, -14, 93, -39, -93, 93, 112, 98, -85, 5, 40, 119, -32, -119, -82, -39, -118, -120, -100, -112, -89, 70, -97, 56, -28, -123, -9, -26, -39, 37, -114, 95, 116, -28, 111, -95, 28, -70, 93, -82, 101, -26, -76, 108, 125, -56, 67, -76, -23, -6, -43, 6, -19, -65, 109, -39, -56, -111, 33, 102, 15, -95, -73, -11, -105, 109, -66, 41, -90, 72, 88, -100, -42, -32, 89, -100, -59, -63, -77, 83, 67, 7, 115, 14, 30, 15, 36, 40, 80, -68, -4, 19, 56, -70, 79, 108, 64, 33, 123, -59, -58, -23, -94, 44, 127, 119, 117, -15, -6, 97, 93, 108, 101, 119, 81, -34, -21, -94, -22, 43, -123, -55, -67, -44, 41, 80, 57, 14, -109, -37, -96, 27, -67, -58, 123, 84, -92, 67, -66, -116, 68, -60, -32, 15, -30, -57, -20, -105, 39, -107, -73, -66, -16, -64, -120, 51, 10, 52, 28, 1, -101, 103, -88, -60, -98, -124, -73, 68, -15, 61, -124, -92, 108, 91, 26, -68, 84, 118, -90, -72, 34, 89, -21, 109, 78, 107, 112, 63, 28, 52, 108, 71, 10, -94, -68, -103, 116, -114, 82, 110, 36, 34, -27, 109, -121, -72, 94, -93, 110, 54, 82, -120, -77, 52, -83, -112, 36, -119, 51, 57, 123, 42, 36, -97, 124, 15, 54, -2, 93, 11, -111, 108, -71, 120, 64, 103, -95, -13, -42, 34, 89, -62, -20, 75, -107, -95, -68, 102, -37, 96, -70, -106, 28, -87, 18, 94, -39, -29, 32, -128, 23, 37, 27, -20, 16, 55, -126, -125, -48, -119, -118, -6, 114, 51, 61, 25, -121, -3, -55, 7, 100, -94, -12, 89, -14, -122, 28, 64, 105, 80, 23, -55, -102, 93, -2, 83, 17, -88, -48, -63, 3, -102, -127, -104, -68, -111, -18, -103, -30, 34, -73, -36, -97, -119, 7, 97, -52, -71, -36, 60, 55, 52, -83, -58, -62, -33, 127, -103, 11, 2, -15, 49, 29, 45, 70, 77, -121, 33, 67, 1, 115, -87, 19, 92, 41, -70, 109, -49, 80, 9, 38, 103, -92, 119, 85, -85, 74, 86, 10, 26, -35, -22, 118, 66, 19, -14, -37, 124, 24, -82, -30, 31, -15, 92, 123, 14, -117, -106, -65, -101, -78, -46, -37, -28, 38, 23, -128, 70, -87, -87, -24, 100, -41, 110, 17, 111, 100, 28, -4, -113, 49, 25, 27, 33, 10, -68, -91, 36, 61, -23, -9, 68, 110, -70, -103, 27, 105, 44, 2, -119, -127, -70, 124, 6, 0, 18, -27, 50, -99, -79, 19, 71, 73, 103, 37, -105, 8, 37, 116, -57, 16, -14, 65, 25, -37, 96, -81, 72, -61, -87, 69, 123, -110, 16, 125, -60, -66, 112, -115, -118, -71, -71, -13, -75, 33, 110, 42, -105, -73, 10, 49, 115, -11, -46, 88, -63, -18, 82, -42, 85, -25, -55, -32, 77, -106, 93, 57, -54, 71, 84, -19, 123, -37, -51, -126, 121, -125, -64, 98, -32, 44, -63, -122, -17, -15, 87, -89, 41, 94, 64, 46, 99, -75, 17, -85, -29, -36, -65, -92, 11, -20, -21, 52, 64, -96, -70, -22, -40, 101, -86, -57, 125, 61, -21, -123, -122, 22, -18, -69, -44, 43, -19, 42, -123, 14, 23, -66, -37, 24, -119, 4, -36, -53, 117, 103, -33, 18, -68, -57, 112, 9, 87, -40, 87, -2, -46, -42, 73, -73, 124, 92, -88, -116, 67, -58, 80, 103, -102, 75, -91, -49, -88, 11, -80, 83, 108, -86, 38, -43, -66, 34, -6, -102, -11, 75, 31, -103, -59, 126, 75, -51, -60, 74, -22, 26, 65, 5, 73, -58, 96, 102, -63, 119, -70, 84, 112, -112, 95, -45, -44, -64, -34, 41, 21, 97, 118, 72, -107, -23, -24, -8, -126, 21, 56, 48, 102, -125, -95, 111, -81, -2, -4, -37, 32, -68, 88, 52, 109, 93, -109, 69, 7, 95, 111, -48, 123, -71, 28, 29, -11, -118, 30, 56, -52, -83, -57, -16, -2, 105, -47, -49, 57, -119, 63, -104, -12, 47, -95, -80, -93, 35, -36, -120, -89, 18, -37, 57, 44, -3, -70, 39, -57, -69, -90, -70, -63, -108, -84, 33, 30, 37, -34, 55, -35, -95, 84, 13, 82, 71, 120, -34, -24, -66, 21, 44, -40, -103, 70, 124, -27, -92, -61, -48, -9, -63, 5, 31, -105, -126, -24, 80, 6, 74, 86, 120, -59, 18, -95, 96, 116, 92, -15, 24, -20, -22, -127, -103, 53, 115, -20, -34, -90, -39, -68, 44, 123, 60, -79, -87, 50, -66, -55, -10, 118, -75, 75, -48, 77, 3, 125, -65, -87, 76, 102, -25, 71, -115, -62, -39, -99, -2, 103, -42, 118, -27, -87, -4, -15, -118, 19, 68, 46, -30, -124, -106, 117, -31, 124, 79, -54, 79, 46, -60, -43, -29, -86, 16, -49, -119, -25, 84, -63, 31, 126, -119, -27, -10, -9, 124, 124, -48, -32, 116, 50, -43, 15, -110, -95, 77, -43, -44, -35, 52, 38, 11, -2, -18, 93, 11, -83, 0, -12, 26, 114, -68, -4, 27, -90, -11, 12, -34, -91, 32, 72, -110, 22, 43, 72, 55, 36, 127, 106, -67, 94, 94, -77, 91, -15, 73, 69, -65, -10, 89, 41, 67, 79, -86, -11, 61, 2, -23, 70, -4, 61, -13, -122, -16, 15, 45, 112, 44, -4, 122, 0, -9, 40, 126, 93, -44, 50, 2, -125, -114, -98, 30, -30, -86, 9, 67, 38, -52, -14, -103, 73, -10, -80, -84, -106, -57, 102, 76, 81, 59, 2, -53, -9, 116, 42, -8, 97, -5, -39, -6, 77, 118, -64, 4, 78, -81, -15, 6, -39, 103, -3, 5, 100, -31, 47, 17, 22, -62, 95, -65, -51, -105, -123, -81, -100, -55, 102, 93, -103, 119, -8, -117, -124, 111, -127, -34, -8, 55, -44, 110, -55, 81, 2, -69, -91, -3, -17, 56, 55, -65, -107, -60, -104, -2, -81, -67, 89, 97, 30, -121, -61, -127, 73, 61, -46, 16, 73, -113, -9, -116, -116, -77, -107, -122, 59, 73, 56, -83, 25, -21, -2, 73, -101, 40, -64, 112, -6, 35, 20, -22, 32, 29, 110, -107, -40, -25, 6, -123, -23, -8, 6, -71, 68, 74, 104, 113, 119, 15, -95, -125, -104, -26, -53, -122, 122, -45, 27, -3, 20, 18, -104, 34, -31, -50, -101, -33, 127, 84, -83, 101, -62, 97, 76, 54, 92, -27, 100, -4, 4, 122, -9, 94, 9, -105, -44, 61, 25, 61, 87, 9, -28, -32, -9, -14, -29, 73, 52, -90, -39, -52, 124, 97, -52, 2, -128, 111, 86, 107, 76, 18, 114, -109, 73, 22, 125, -59, 56, -50, 118, -32, -86, -97, -21, -117, 49, 7, -42, -98, 95, -20, 27, -67, -4, -72, -41, -104, -12, -59, 24, 110, -94, -54, -5, 83, -69, -85, -66, 86, 31, -59, 123, -93, 108, 57, 79, -44, 82, -8, 29, -25, -42, -76, -40, 10, -91, 83, 42, 11, 57, 100, 41, 111, -128, -91, 14, -8, 16, -35, -112, 36, 127, -35, 75, 55, 88, -11, 22, -78, -9, 43, -7, -47, -124, 26, 56, -6, -100, 58, 110, -91, 1, -99, -48, 111, -113, 121, -120, 35, 117, 115, 116, -18, -127, -43, -47, 11, -15, 30, -26, -108, -31, -101, -51, 74, 119, -12, -107, 52, -40, -121, 48, 97, -31, 16, 5, -85, -1, 33, 28, 117, -57, -57, 47, 51, -12, -121, -77, 10, -38, 18, -67, 86, 74, -8, -51, -67, 67, 74, 104, -104, -21, 59, -96, -15, 8, -54, -25, -127, -55, 101, 50, 15, 57, -116, 122, 83, -38, 11, -37, -29, -52, -100, 37, 118, 38, 100, -50, 18, -48, -92, -115, 9, 29, -19, -46, 37, 83, 46, 44, 38, 62, -102, 5, 121, 23, 68, -100, -28, -116, 101, -19, 72, 11, -77, 120, -41, -21, 110, 30, -56, 46, 96, -102, -71, -73, -88, 125, 37, 12, -7, 77, -35, 65, -128, -50, 17, 5, -62, -63, 19, -44, 10, -56, 83, 17, 86, -103, -93, 29, -127, -22, -13, -5, 72, 46, -102, 125, 75, -97, -77, -46, -127, -86, 17, 60, 52, -3, -76, 70, 11, -51, 23, -12, 116, 107, -91, -101, -60, -98, -87, -90, -78, -35, 85, 31, 67, -48, -28, -115, 37, -41, 60, 103, -96, 79, -119, 88, 107, 83, 9, 60, 21, -60, 121, -27, 39, 33, 57, 50, 87, -89, 23, 106, 82, 41, -89, 43, -36, -71, -120, -28, 14, 81, -33, -55, -50, 9, -38, -23, -117, 17, -76, 65, -10, 68, -25, 7, 86, -91, 115, 89, -68, -53, -55, -55, -32, 44, 94, 60, -102, -86, 97, -97, 42, -127, 80, 103, 11, -88, 50, -5, 81, -118, -86, 124, 67, 79, 22, 90, 82, -69, 15, -7, -79, 21, -15, -46, 24, -53, -121, -126, 92, 123, 72, 75, -82, 49, -51, 69, 68, -33, 118, 17, -70, -55, 70, 106, 15, -58, -116, 98, 100, -75, -37, -8, 21, -103, -84, 121, -48, -15, -46, -41, -16, -26, 80, -57, -25, -19, -56, 4, -18, 30, 90, 80, 8, -125, -52, -49, -15, -72, -57, 112, 88, -121, 124, 119, 12, -66, 99, -89, -48, -15, -110, 32, -70, -79, -57, -101, -119, -77, 17, -82, -63, -46, -110, -128, 59, 78, 59, -91, -98, -85, -63, 47, 26, -110, -34, -17, 118, -100, -88, -10, -77, 60, 72, -38, 109, -80, -89, 74, -35, -3, 84, 86, 73, -12, -18, -121, 48, 91, 15, 56, -66, -75, -47, 94, 66, -39, -55, -42, 0, 0, 5, 63, 9, 97, -5, -9, -48, 58, -114, -82, -83, 83, 18, 32, -83, 18, 19, -121, -126, -71, -3, 61, -99, 35, -109, -72, 123, -14, 118, -12, 53, 58, 51, -103, -68, -81, -21, -54, 60, 51, 78, -27, 62, 43, -32, -83, 21, -11, -67, -82, -86, 57, -13, -18, -94, -60, -26, 114, 59, 72, 6, -61, 33, 16, -116, -18, -69, -109, -19, -17, -116, 38, 110, -103, 70, -88, 71, 34, -24, 28, -33, 20, 58, 5, -9, -4, -15, -114, 96, 104, -67, 81, -97, -103, 89, 43, 42, 41, -88, -127, -92, 104, -5, 52, -24, -58, -75, 4, 100, -126, -25, 94, 91, 16, -99, 89, -109, 84, -82, -98, 51, 57, -43, -81, 15, 91, -12, 66, -77, 20, -113, 33, 3, -59, -84, -54, 108, 71, -113, -34, -30, -41, 96, -98, 35, 95, 114, 29, 91, -113, 48, 127, 72, 43, -1, 12, -118, -11, -58, 70, -78, -97, 122, -93, 21, -97, 98, 91, 16, -20, -10, 78, -32, -107, -99, -27, -62, 32, 115, 24, -92, 126, -52, -116, 57, -119, -33, -1, -44, -5, -40, -116, 33, -83, 71, -115, 43, 113, 36, -104, 12, -9, -19, 106, -112, 63, -41, -26, -74, -54, 83, -82, -50, -107, -118, 29, 123, 51, 95, -124, 42, 44, 46, -97, 94, -117, 87, 42, -5, -123, -8, -1, -85, 94, 118, -62, -16, -73, 8, 63, -20, -10, -96, -122, 95, -70, -22, -100, -44, 80, 84, -83, 61, 117, -83, -23, 119, -111, -42, 50, -118, -30, -22, 126, -109, 27, 3, 119, -120, 70, -6, -96, 10, 9, -54, 67, -27, 41, -105, -42, 82, 29, -111, 54, -44, -87, 20, -3, -112, -81, 127, -115, 96, 88, -1, 119, -26, -44, 71, -125, 126, -49, -31, -99, -34, 124, -99, -12, -115, -114, 70, -45, -27, 38, -64, 46, -108, -102, -122, -58, -59, 112, -47, -86, 87, 68, -51, 70, -122, -117, -47, -69, 30, 88, 96, -103, -126, -62, 2, -125, -118, -35, -45, 10, -3, 1, -8, -7, 7, -8, 2, 67, -114, 50, 15, 2, -100, -38, -121, -46, 43, -58, 63, 50, 111, -50, 11, -14, -105, -52, -89, 41, -87, -70, -93, -53, 11, 6, -95, -28, -92, -32, -51, 59, -117, 86, -3, -72, 49, -55, -80, 71, 82, -123, 78, -66, -123, 6, 48, -84, 113, -77, -84, 37, -126, 122, -5, 118, 78, 89, 25, -66, -55, -81, 95, 25, -110, -115, -22, 20, -77, -28, 24, 22, -27, 114, 101, 4, 99, 63, 68, -23, -102, 88, 97, 98, 88, 76, -114, -9, 98, 48, 14, -88, -51, 34, -98, -67, -112, -3, -12, 25, -112, 118, 96, -66, -44, -93, 45, 90, 40, -37, 18, 59, -39, 92, -50, 110, 3, 83, -47, 26, -52, 103, -101, -95, -95, -91, -43, -56, 60, 29, -7, -55, -126, -10, -68, 38, 99, 125, -1, 122, -27, 58, 8, -68, 75, -49, 98, 107, -126, 94, -46, 119, 109, -62, 89, -7, -67, 22, 100, 68, 18, -93, -110, 59, -12, 11, -5, 102, -52, 77, -8, -15, 80, 61, 96, 52, -44, 55, -110, 120, -36, -82, 51, 115, 26, 95, -54, 125, 94, 5, 28, -121, 4, -79, 83, 76, -80, -47, 20, -72, 25, 80, 44, -50, 95, 35, 40, -107, -38, -24, 56, 124, 80, 27, -82, 46, -64, -43, -71, 19, -13, 5, 61, -28, 24, 109, 10, 116, 98, -1, -65, -95, 87, 115, -32, 68, -47, -85, 89, -55, -100, 54, 65, 41, 27, -11, 42, -7, 47, -86, -1, -107, 47, 1, -98, 25, -64, -111, -121, -105, 3, 108, 5, 123, -35, 1, 125, 99, -13, -39, 11, 7, -67, -22, -123, 44, 27, 38, -19, 71, 90, -10, 124, 84, -40, 12, 35, 112, -41, 5, 89, 29, -22, 78, 19, 85, -125, -13, 53, 121, 115, 104, 126, 73, -22, -126, 109, 71, -47, 69, 118, -45, -48, 94, -48, 51, -75, -24, 64, 61, 14, -77, 5, -48, -31, 109, -22, -87, 122, 122, -33, 24, 0, 58, -87, 4, 8, -127, 111, 10, 27, -60, -82, 51, 22, -54, -46, -81, 1, 113, 88, 56, -115, -74, 1, -112, 26, 70, -34, 61, 46, -17, -21, -110, -82, -84, -125, -115, -39, 127, -27, 109, -57, 79, -47, 100, 79, -22, 98, 44, 69, 118, -96, -50, -11, 1, 30, 117, 23, 45, 110, 58, -90, 116, 104, 75, 8, -68, 102, -32, 125, 99, -43, 13, -6, 110, -62, -66, -10, -41, 20, -68, -73, 93, -57, 90, -79, 65, -61, -64, 110, 68, 97, 127, -9, -101, -21, -91, -2, -46, 77, 42, -64, 62, 5, -115, 60, -15, 93, 55, 117, 1, -110, 75, -77, -1, -36, -125, -92, -10, -12, -46, 121, 104, -22, 29, -3, -23, -39, 101, -86, -21, -39, 24, -111, 72, -102, 81, -89, -49, 74, -41, 35, -92, -53, 90, 7, -45, -41, -1, -9, 15, 30, 59, 31, -108, -102, -10, -52, 127, -37, 98, -23, 14, 96, 38, 28, -23, 37, -18, -86, -98, 94, -121, -119, -43, 96, 96, 59, 106, 122, 23, -120, -93, 30, 85, 54, -115, 67, 106, 10, 26, 2, 116, 123, 116, 50, 80, 65, -21, 95, -64, 63, 11, -122, -30, 79, -47, 97, 100, 113, 21, -86, 4, 27, 8, 48, 101, -62, -115, -7, 119, 34, -120, -23, 53, -2, -97, 24, -29, 76, 4, -93, -91, -46, -25, -112, 34, 33, 7, 48, 47, 124, 105, 60, -16, 71, 40, -99, 91, -117, -24, 119, -11, 104, 18, 63, -38, 89, -53, 115, 77, -25, 60, -87, 11, 107, -9, -27, -42, -36, -27, -79, 17, 99, -73, 7, 93, 1, 26, -21, -114, -60, 17, -86, 7, -27, -56, -48, -47, 98, 31, 92, -110, 98, 100, -82, 103, 42, -126, 102, 124, -55, -56, -126, -33, 56, -81, 49, -1, 51, -70, -120, -120, 49, 25, 31, 112, -80, -82, 90, -15, 8, -19, -8, -80, 107, -91, 85, 7, -14, 28, 106, 2, -54, -54, 50, -86, 12, 105, 117, 32, 67, 69, 6, -111, -4, -31, -8, 118, 58, 107, -71, 13, -82, -66, 6, -42, -97, 39, 48, 65, -107, 50, 92, -29, 27, 126, -46, 14, 2, 82, -20, 14, 72, 85, -112, -108, -96, -97, 115, -61, -9, 31, -26, -27, -62, 100, -109, 62, -95, 33, -127, 51, -32, 112, -105, -112, -14, -7, -112, 2, -34, 81, 36, -106, 8, -38, -52, -121, 46, -42, 50, 28, -72, 48, 34, -3, -118, 1, 55, -22, -58, 94, -69, 64, 68, -21, 121, 4, -3, -37, -55, 74, -14, 16, 114, 96, -117, 113, -114, -73, -6, -84, 68, -45, -20, 8, 124, -11, -88, 105, 20, -43, 31, -90, -18, 36, 84, 47, -26, -112, -44, 114, 13, 121, 48, 93, 68, -105, 110, 48, -97, 101, -16, 76, 46, 99, -81, -41, 29, -96, -25, 73, -104, 115, -18, -115, -7, 78, 4, -120, -33, 13, -16, -55, -72, -57, -16, 115, -2, 77, 3, -35, 54, 6, 10, -28, 20, -32, -7, -64, -46, 77, -110, -48, 127, -89, 3, -36, -30, 97, 55, -104, 43, -119, -30, -58, -51, -42, -62, -123, -32, 102, -80, 72, -37, -77, 28, 42, 108, 103, -40, 26, -26, 86, 20, 62, 79, -29, 6, -107, 97, -114, 82, -4, 116, 11, -87, -61, 44, -85, 25, 26, -10, 113, 27, -96, -54, -44, -109, -19, -98, 95, -98, -1, -55, 114, 113, 56, -27, -105, 25, -107, 126, 115, 74, 98, 72, 67, 56, 89, 20, 102, 22, 102, -23, 56, 56, -72, 121, -105, 47, -23, -19, -35, -75, -35, 64, -112, -74, -106, 61, -38, 89, 28, 3, -46, -12, 2, 5, -51, 70, -26, -58, 4, -27, 58, 77, -37, -32, -55, 20, -123, 70, 55, -36, 119, -11, -123, -42, 60, -84, 1, -74, -30, 44, -49, 118, 21, 93, 33, -58, 90, 49, 10, -68, 55, -11, 3, 16, 108, 75, 83, 81, 95, 114, 98, -49, -83, -44, 24, 72, 11, -38, 110, -106, 54, 50, -118, -74, 122, -24, 96, 122, 37, -45, -19, 30, -76, -73, 54, 121, -77, -90, -47, 28, 42, 28, 83, 107, 6, 76, -122, 106, -61, 53, 99, -123, 120, 48, -107, -84, 27, -38, -21, 55, -125, 120, 42, 122, -34, -90, 61, 109, 55, 38, -86, -46, -20, -57, 47, 54, 65, 112, -4, -6, -8, -105, -100, 124, -96, -74, 117, 52, -63, 48, 3, -36, 16, -97, -111, -32, 37, -63, -106, -40, 15, -83, -21, -19, 113, 86, -96, 45, 30, 104, 29, 69, -34, -15, 115, 64, -96, -76, -77, 23, 68, 90, 66, -106, -92, 83, -26, 72, -70, 119, -2, -97, 88, 69, -76, -109, 76, -84, 17, 9, 87, 24, 31, 95, -36, -42, -127, -73, -89, 122, 54, -58, 7, -59, 56, 61, -12, -71, -12, 24, -42, -30, 111, -95, 75, -113, -98, 96, -111, 117, 118, 121, 60, 87, 101, 19, -47, 41, 115, 70, 108, 3, -112, -84, 36, -120, 64, -75, -57, -89, 72, -4, -39, -46, -29, 70, 10, -48, -27, -21, -111, 77, 49, 16, -67, 36, -127, -126, -1, 73, 66, -92, 87, -8, -40, 80, 0, -97, -45, 89, 4, 24, 120, 94, -114, -82, 99, 46, -101, 121, 7, -72, 69, -16, -116, -79, 57, 59, 88, 91, -120, -14, -71, 15, 38, 124, -114, -37, 49, 125, 25, -56, -9, -7, 101, 117, -115, -85, -59, -24, 110, -113, 108, -11, -70, 13, 106, -128, 54, 51, -36, 97, -56, -8, -59, 64, 16, 86, -83, 31, 34, 44, 71, -62, 40, 86, -126, 27, 124, -86, 24, 0, 26, -50, 38, -111, 106, 12, -28, 94, -90, 27, -14, 126, 12, -82, -14, 16, 72, 1, 53, -122, -9, 115, -107, -40, -5, -16, -1, 47, 3, -121, -56, -27, -19, 23, -15, -27, -50, 37, -20, -46, -29, 55, 83, 74, 114, -59, -46, -96, -2, 114, 125, 51, 77, 41, 24, 54, 17, 42, 41, 72, 45, 44, 84, -45, 83, 49, 70, 127, 94, 115, 118, -53, -6, -58, -106, 33, 58, 62, -79, 53, 72, -29, -79, -95, -13, 107, -8, 63, 63, -7, 85, 44, 116, -83, -81, 110, -19, 113, 99, 105, -105, 74, -23, 74, 127, 66, 26, -83, 78, -62, -128, 49, 74, 66, 77, -27, -74, 5, -127, -65, 92, 113, -111, 110, -59, 103, 93, 108, -83, -10, -4, 27, 49, -38, -95, 43, -77, -50, -56, 16, 3, -60, -6, -63, 17, 64, 53, 39, 106, 104, 74, -98, -48, -118, -18, 74, -34, -26, -62, -47, -56, 3, 126, -87, -63, 100, -34, 61, -61, -123, 15, -47, -45, 63, 125, -120, 116, 33, -116, -75, -20, -79, 105, 6, -44, -31, 88, -10, -58, -56, -41, 73, 113, 18, -81, 54, 17, -123, -95, -11, -114, -102, -55, 0, -40, 22, -118, -49, -55, -121, 121, -64, 32, -21, 109, 102, 86, 24, 113, 72, 32, 95, -126, 28, -50, 61, -66, -3, -28, 79, 127, -103, 23, -46, 110, -71, 53, 65, -119, -37, -92, -103, 0, 18, -92, 111, 6, -75, -112, -92, 51, -103, -49, -52, -123, -63, -49, 82, 48, -6, -127, -22, -109, 46, 83, -89, -104, -12, -37, -42, 7, 32, 123, 84, -55, 42, 13, -82, -26, -91, -90, -114, -36, -115, -81, 118, -71, 79, 70, -77, -9, 56, 100, 75, -73, 89, 88, -74, 86, 57, -78, 55, 22, -52, 18, -118, -116, -91, 97, 98, -73, 57, 89, 13, 125, -127, -69, -26, -52, -64, -105, -115, -104, -4, 90, 91, 74, 111, 16, -51, -29, 66, -41, 112, -51, 43, -48, 83, 33, -15, -76, 7, -13, 16, 14, 58, -9, 78, -36, 47, 106, -15, -88, -40, -26, -101, 40, -41, 92, -50, -127, 35, -40, 103, 98, 113, -41, -38, 34, 24, 109, 29, -81, -36, -9, 17, 47, -45, 87, 66, 13, -7, 108, 2, -47, -69, -47, 24, 52, 6, -52, 63, 29, -106, 76, -40, 19, 27, 119, 115, -127, 110, 25, -40, 9, -68, 20, -70, 92, 123, 115, -23, 80, -11, 97, 24, -83, 88, 46, -118, -19, 112, -69, -62, 55, -66, -103, -36, 92, -88, -127, 63, -58, -128, -85, 84, -4, 92, -85, -30, -52, 58, 52, 32, 75, -16, 32, 92, 16, 13, -125, 80, 42, -26, -100, 21, -45, -3, -27, -85, 48, -61, -111, -43, -83, 91, 89, 107, 78, -90, 113, 83, -114, 31, 80, -24, 70, 44, 111, 17, -122, 70, -86, -62, -54, -47, -2, 116, -98, 23, -6, -1, 124, -88, 105, 92, 0, -8, 25, -62, 48, 19, -18, 35, -40, -32, 57, -92, -81, 53, 92, -36, -85, -23, 32, 36, -74, 94, -124, 117, -31, 20, 29, 112, 62, 38, 84, -21, 120, -76, -111, -16, 52, -42, 46, 13, 88, 102, -8, 5, -35, 122, -36, -128, -98, -2, -16, 114, 23, 35, 0, 120, 5, 23, 105, -107, -90, -107, 56, 36, 82, -15, -98, -128, -16, 58, -65, 35, -118, -6, -58, 56, 37, 20, -19, -51, 83, 6, 119, -89, 63, -7, -55, 89, -8, 105, 20, 118, 57, 105, -47, 26, -100, -92, -110, 124, -94, -68, -110, -110, 19, 61, -122, -22, 125, -7, 107, 123, -74, 73, 34, -12, -7, 83, -71, -60, -6, -32, -99, 117, 34, 44, 62, 119, -128, 109, -30, -71, 14, 44, -42, 17, -25, -64, -78, -66, -90, 10, -44, 63, -43, 29, -16, -69, -51, -41, -37, -121, -32, 5, -17, 81, 38, -87, 70, -68, -57, -105, 57, -125, 32, -94, 56, 62, 39, 78, 49, 43, -61, -71, -89, -75, -102, -108, 120, 78, 109, -68, -19, 106, 76, 26, 107, -23, -33, -117, 68, 59, -52, 12, 67, -70, -63, 61, 72, 120, -110, 115, -30, -121, 102, -47, -116, 14, -44, 119, 8, 2, 32, 16, -59, -59, -33, -24, 64, 95, 89, -78, 54, -64, -45, -100, -106, 20, -61, -97, -96, -54, 74, 75, 111, 91, -2, -88, -4, 18, -45, 17, -55, 103, -34, -88, 109, 70, -87, 69, 78, 126, -124, 75, -60, 73, 89, -10, 30, -57, 24, -25, -23, 72, -112, 82, -44, -71, 54, 27, -88, -12, 107, -46, 103, -119, -69, -121, -89, 104, 126, 62, 85, 89, -78, 76, 88, -95, 26, 65, -4, 108, 77, -25, -8, 89, 9, -122, 91, -77, -28, 43, -16, 125, 126, -73, 17, -85, 30, 9, 13, -14, 67, 18, 21, -42, -91, -20, 93, -89, -76, -44, -112, 123, 21, 1, -100, 6, 56, 24, 111, 20, -116, 29, -65, 16, -75, -58, 99, -99, 4, -54, -116, 35, -121, -53, -71, 96, 79, 3, 21, 112, 102, -70, -83, -32, -36, -98, -81, 81, 112, -24, 91, 19, 48, 76, -88, 71, -43, 113, 13, 72, -13, 11, -88, -83, 49, -76, -47, -62, 112, 9, -26, 72, -3, -103, 64, -49, -55, -82, -127, -72, -46, -18, -23, -24, -38, 108, 27, -87, 78, -10, 52, 19, -15, -102, 41, -124, 99, 33, 49, 47, -59, -17, -46, -47, 54, -17, 114, -94, -55, 79, 118, 106, 94, 78, -10, 94, 37, 18, -70, 0, -34, 41, -56, -32, -86, -42, 58, -26, 75, -38, -76, -68, -111, -122, -34, 109, -22, -25, -73, -101, 116, 62, 103, 67, -33, -1, -49, -100, 11, -2, -103, 84, -26, 83, -91, 99, 2, 70, 86, 67, 121, 118, 64, 25, -115, 120, 86, 40, -69, -125, -121, 30, 9, 7, -42, -32, 10, -57, -78, -123, 56, 7, 40, 123, 109, 68, 100, 66, 56, 110, -125, -112, -78, -19, -20, 71, -21, 22, 63, -50, 57, 0, -68, -1, 127, -12, -4, -107, 75, -44, 35, -104, 26, -60, 63, -111, 88, -77, -19, 72, 74, -125, 24, 78, 59, 94, 73, 13, -38, -18, -64, -26, 89, 54, 110, -66, -59, -55, 99, -96, 110, -19, 37, -117, -88, 80, 13, 90, 116, -65, 123, 81, -83, 56, -77, 59, 54, 75, 89, -67, 79, -117, -81, -43, 35, -112, 123, -97, 89, 115, 3, 115, 99, 87, -97, -87, 8, -75, -116, -64, 29, -76, 87, 76, 119, -44, -91, 100, 107, 12, -47, 100, 51, 43, 78, 75, 25, -113, -118, -8, 123, 11, -36, -57, 118, 1, 32, -66, 107, 13, 93, 33, -92, -44, -73, 61, 26, 104, 91, 8, -119, 124, -125, 48, 112, 123, -18, 97, -41, 32, 17, 42, 35, 125, -124, 127, -111, 120, 100, -94, 117, 59, -112, -99, -25, -34, -58, -89, -30, -69, -116, 33, 115, 78, 2, -101, -4, 83, -33, 11, 20, 16, -112, -84, -90, -121, 119, -69, -70, 97, 31, 6, 11, 46, -112, -16, -53, 109, -94, 61, 51, 14, 112, -124, -89, -72, -66, -63, -41, 122, -19, -64, -100, 53, 125, 38, -85, 44, 126, 98, 107, 76, 32, -35, -79, 73, -58, -33, 51, -79, -81, 79, 29, 122, 55, -88, -17, -98, 88, -91, 62, 5, 23, 100, 114, -39, -115, 31, -71, -60, -30, 108, 115, 122, 58, -77, -99, 5, 115, -53, -18, 43, -51, -49, 3, 15, -93, -24, -49, 111, 43, 122, -102, -10, -16, -123, 36, 29, 42, -41, -8, -47, -20, 72, -68, 39, -24, 59, -121, -52, 123, 114, -126, 11, -20, -87, -71, -127, 42, -90, 83, 84, -115, -41, 95, 104, -9, 92, -79, -48, 6, -15, -37, -49, 50, -61, 120, 26, -120, 105, -73, -104, -88, -85, -1, 99, -75, -57, -114, 45, 81, 111, 39, -90, 86, -103, -82, -16, -42, 85, 105, 17, 39, 126, 88, -19, 99, 42, 46, -42, 68, -126, -121, 46, -73, -52, -47, -20, -13, -117, 112, 60, -74, 52, 116, -28, 124, -60, -55, 36, 46, -123, -118, 18, -16, -36, -105, -6, 22, 89, -70, 108, -100, 96, 86, 91, 16, 6, 100, -55, -31, -13, -69, -13, -4, 43, -9, -72, 16, 84, -56, 98, -37, 8, -20, -83, -49, -15, -8, 74, 8, -81, 1, -22, -118, 97, -56, -92, -12, 20, 33, 28, -88, 28, 57, 9, 117, 118, 52, -48, 36, 112, 110, -35, 32, -60, 89, -43, -121, 47, 27, 102, -74, 92, 53, 12, 64, -26, 52, -25, -5, 121, 79, 123, 52, 117, 33, -39, 4, 76, 20, -36, -104, -13, -6, 23, 124, -106, -31, -71, -37, -65, 89, 101, 69, 31, 89, -105, 61, 105, -42, -126, -40, -28, 55, -52, -40, 88, -1, -22, -6, 46, -28, -72, 126, -55, 109, 72, -4, -23, 7, -52, 99, 1, 13, -49, 104, 45, -48, -82, 59, -42, -37, 0, -1, 32, 25, -42, -86, -48, -4, 20, -84, -13, -30, 49, 66, -69, 95, -127, -5, 79, 72, -79, 52, 32, 46, -24, -100, 48, -125, -36, 22, -6, -26, -10, 90, -31, -37, 107, 20, 66, -60, 1, -14, 47, -124, -6, -4, -59, -70, -105, 7, -119, 69, -127, 40, 67, -49, -16, 28, -18, -21, 31, 65, 23, 21, -21, 87, 77, -30, -75, 108, -115, 52, 59, -25, -7, -73, 60, -87, 61, -125, 65, 19, -122, -7, -73, -57, -3, 42, 122, 106, -115, 111, 5, 40, -90, 125, 112, 14, -116, 74, -1, 21, -43, 36, -41, 102, -68, 49, 50, 55, -128, 50, 68, -108, -117, -87, 29, 11, -59, 96, -10, 105, -5, -69, -47, -76, 37, 109, 89, -38, 92, -46, 115, -115, -1, 3, -53, 2, 1, -61, -114, 23, 29, 121, 42, 56, -128, -46, 100, -99, -81, -46, 14, -41, 98, -118, 110, -124, -32, 4, 62, -96, 75, -44, 99, 111, -67, 69, 27, -86, 115, 115, -14, -66, -18, -4, 100, 71, 17, -82, 11, 97, 70, -91, 113, 9, -66, 75, 72, -2, 84, 79, -6, 95, 3, 62, -63, 107, 6, -52, -99, 70, 98, 39, 111, -50, -121, 91, -39, -38, -116, -68, -29, -55, -24, -127, 61, -83, 88, -28, 88, 111, 34, -7, -26, -97, -60, 32, 85, -42, 78, -16, 44, -50, 73, 114, -32, -76, 37, 79, -33, -101, 71, -91, -85, -38, -126, -102, -44, 16, -40, 112, 89, -91, -107, 96, -53, 57, 24, -46, 81, -95, -38, 62, 53, -4, 95, 108, -70, -13, 12, 125, -86, 33, 103, -90, -15, -97, -15, -64, 78, -36, -111, 1, 52, 115, -35, 35, -68, -82, 51, 51, 22, 10, -61, -118, 29, -57, -11, 72, -88, 119, 103, -9, -28, 31, -125, -54, 98, -102, -14, -42, 56, -42, 81, 96, 39, 33, -73, 59, 16, 107, -41, -109, 51, 10, 48, 36, 6, 81, -56, -12, -5, -107, -71, -116, 105, 94, 75, 110, 26, 123, -123, -12, 100, -66, -74, 71, 10, -101, -31, 65, -106, -94, -27, -98, -25, 7, -76, 58, -55, 119, -103, -25, -52, -52, 70, 51, -70, -5, -43, 64, -3, -77, -77, 107, -9, 91, 116, -52, -48, 43, 103, -41, -98, 106, 104, -105, 19, 108, -84, -116, 108, 61, -12, 124, 18, -94, 10, -33, 113, 93, -82, 92, -100, -54, 123, 104, 8, -82, 62, 123, -76, -40, 56, -92, 104, 90, -118, 92, 102, -80, 89, -44, -127, 19, 10, 56, -50, 68, 16, -13, 66, -54, -79, 109, -106, -76, -114, 59, 51, 97, 99, -101, -5, 35, 79, 107, 50, 10, 90, -95, 95, -40, 103, 58, -44, 107, 64, -9, -43, 106, 67, -90, -127, 14, 87, -57, -21, -56, -90, 51, -65, -44, -116, -125, 124, 41, 83, -6, -30, 110, -105, 39, 105, 102, 125, -98, 2, 75, -86, -32, -87, 39, -56, 81, -84, -97, 75, -89, 39, 58, -14, -120, -77, -11, -10, -36, -24, -12, 121, 54, -87, 2, 8, 52, 96, -32, -91, -92, -127, 118, -117, 127, -38, -102, -95, 108, 88, 17, -44, -5, -30, -33, -100, -126, -57, -74, 101, -9, 85, -65, -69, 49, 21, 89, 28, -62, 36, 36, 3, -61, -56, 26, 80, 22, -99, 41, 70, 102, 16, -114, -108, -116, -92, -32, -55, -104, 87, -43, -50, -32, -19, 26, -50, -110, -63, -33, -70, 76, 47, -76, -125, -24, 86, -15, 74, 9, -105, 9, 24, -50, -104, -17, -21, -101, -18, -33, -79, -69, 13, 76, 120, -8, 81, 74, 8, 33, -49, 36, -73, 61, -102, 81, 97, 103, -30, -123, -29, -32, 72, 112, -45, -68, 116, 48, 64, -97, 2, -118, 54, -25, 81, 22, 9, 101, 4, 13, 66, -27, -58, 34, -40, -38, -104, 37, -5, -124, 77, 44, -57, -34, 9, -87, -59, 29, -121, -5, -81, -102, -123, -121, -113, -126, 60, 115, -108, 44, 127, -58, -61, 87, 87, -113, -7, -99, -77, -12, -58, 77, -29, 113, -72, -98, -27, -52, -88, -11, 55, 61, -26, -11, -12, -6, 72, 56, 125, -3, -37, 47, -19, -52, 59, -20, -107, -83, -34, 107, -90, -61, -29, -8, 20, -92, -70, -109, 96, -109, -4, 21, -125, 45, -17, -103, -125, 16, 62, 14, 28, -99, -117, -5, -74, 117, 0, -15, -51, -69, 69, -57, 79, 50, -13, -128, 85, -32, 54, 39, -91, 41, 90, 52, 123, 5, 40, -107, 20, -103, -79, 96, 17, -50, -18, -25, -32, 25, 17, 44, 99, -101, -15, -93, 32, 54, 9, 23, -83, 2, -12, -44, -32, 79, 116, -118, -116, -53, 31, 113, 55, 109, -54, -23, 0, 115, 67, -100, -43, 20, 9, 3, -47, 102, -38, -95, 92, -97, -14, -50, -113, -8, -95, -91, 127, -93, -49, 69, 112, -119, 28, -66, 97, 71, -88, 80, 126, -68, 98, 37, 106, 18, -12, 22, -30, -62, 40, -87, -99, -7, 50, -33, 37, 88, -26, 9, 99, -100, -122, -58, 24, -94, 74, 2, 127, 71, 94, 52, 39, 69, -10, 34, 10, -98, 97, 7, 21, -32, -74, 58, 69, 39, 84, -68, -22, 24, -59, 1, -124, -127, -68, -88, -40, 68, -39, 24, -87, 70, -53, -96, -79, -67, -3, -58, 88, -48, 126, -5, 71, -41, -43, 96, 53, -86, 8, -11, 104, -111, 49, -38, -1, -79, 124, -19, 110, -112, 12, -120, 72, 30, 77, -70, 49, 110, -15, -23, 120, -79, 122, 50, -9, 48, 95, 123, -31, -62, -126, -116, 20, -17, -57, 78, -125, -12, 106, -37, 23, 39, -10, 34, -20, 127, 118, -111, -89, 127, -25, 28, 102, -77, -74, -106, 75, 34, -72, -116, 89, -31, 112, -103, 124, 20, -90, -124, -119, -57, -33, -45, -115, -87, 68, -100, -29, 31, 29, -51, 29, 80, -35, 119, -113, 35, -116, -10, 14, 87, -20, 67, 55, 23, -120, -8, -66, 115, 34, -12, -127, 66, 60, 0, 94, 39, -75, -51, -8, 50, -45, 56, -77, -111, 77, 9, -18, -23, 41, -56, 22, -111, -79, -2, 98, 33, 21, 105, 19, -50, 77, 72, -2, 82, 19, 4, 82, 36, 47, -109, 88, 121, 42, -109, -53, -85, -34, 41, 99, 25, -28, 31, 98, 104, -69, -73, -47, -22, 72, 60, 90, -14, 65, 121, 11, 80, -68, 21, -124, 77, 66, 109, -44, -39, 76, 118, -115, -12, 125, -4, -30, 108, -126, 97, 99, -118, 60, 13, 27, 109, 65, 117, -88, -45, 11, 126, -41, 34, -28, 50, 62, 93, 83, -72, -36, 94, 81, 37, 34, -58, -7, 116, 22, 9, -33, -22, 110, -40, -98, 121, -55, 5, 54, -6, 104, 17, -118, -1, -62, 0, 41, -12, 52, -107, -118, 30, 114, 6, 21, 112, -32, 102, -96, -70, 104, -78, 18, -10, -56, -25, 18, -76, 89, -32, -79, 49, -84, 93, -7, -96, -7, -57, 78, 114, -112, -13, -12, -42, 46, -122, 115, -33, -76, 12, -71, 39, 97, 116, 72, -125, 15, -35, 51, -62, 49, 37, 34, 70, 6, 9, -5, 76, -19, -126, 102, -93, 92, -86, 111, 52, -21, 24, -45, -50, -122, -109, -80, -29, 39, -30, -5, -74, -53, 12, 80, 16, -57, -46, 122, -128, 10, 26, -28, 3, 77, -38, -50, -112, -10, -1, -97, 125, 81, -18, 124, -27, -67, 2, -18, 89, -56, -115, 52, -80, 55, -21, -55, 97, 15, 25, -102, 117, 15, 9, -30, 35, -116, -56, 121, -4, -23, 8, -119, 78, -92, 7, -7, -121, -119, -86, 111, -6, -121, -61, 26, -122, -91, -81, -44, -17, 25, 46, -82, -65, 97, 46, 46, 84, 27, 38, 70, -26, 101, -71, 122, -34, 12, 10, -20, 70, -59, -48, -4, 101, 59, 2, 16, -104, 118, 116, -73, -100, -90, 127, -52, -105, 68, -40, -41, -74, 57, 95, 101, 15, 116, 51, -116, 31, -110, 59, -59, 26, -78, 106, -103, 28, 98, 90, 58, 36, -35, -97, 38, 75, 68, -65, 106, -42, -121, 74, -63, 118, -24, -55, -99, 24, -91, 84, -11, 26, -37, 89, -69, -35, -47, -61, -77, -121, -47, -14, 117, -30, 120, 43, 105, 70, 89, 42, 126, -101, -4, 8, -54, -107, 30, -127, 25, -125, 81, 24, -54, 46, 87, -126, -115, 12, -45, 27, -126, 76, -81, -55, 60, -65, -70, -33, 87, -128, 48, 102, 25, 58, -42, 90, -76, 94, -55, -29, 21, 30, -61, -18, 56, 97, 85, 1, -38, 93, -31, -25, -33, 4, 24, 41, -109, 4, -46, 37, 7, -13, 86, 39, 67, 31, -100, 89, 117, 123, 57, 124, -1, -104, 123, -53, 103, -119, 82, 35, -123, -20, 89, 34, -95, 56, 48, 19, -90, -33, 22, 78, -55, -44, 65, -78, 106, 117, 21, 10, -90, -128, 126, -80, -87, 115, -84, -45, 94, 5, -112, 10, 4, 9, -84, 118, 60, 3, 33, -60, -68, 82, -62, -118, -50, 48, 41, -55, 73, -85, 83, 38, 115, 120, 86, -101, -38, -104, 52, 21, -69, -31, -68, 67, -106, -65, -63, -69, -50, 53, -68, -26, -119, 86, 76, -124, 107, -87, -62, -56, -48, 14, -109, -74, 100, 53, -128, -114, -35, 11, -8, -77, 43, -82, -97, 52, 62, 98, -116, -40, 41, 64, 59, -121, -81, -10, 97, 96, -120, -87, -84, -74, 33, -88, -41, 61, -1, 40, 82, -77, -55, 21, 120, -92, 96, -33, -83, -11, 83, -98, -9, -102, 110, -115, 126, -17, 113, 73, 29, -30, 48, -109, 36, -117, -85, -41, 74, 126, -34, 54, -100, -88, -97, -120, -111, 85, -109, -39, 0, 106, -100, 102, 54, -66, 29, -101, -96, -61, -87, -65, -95, -117, -94, -39, 62, 50, 21, -39, -31, 41, -124, 20, -87, 8, -4, 26, 75, 15, 81, 113, -103, -25, -41, 88, 73, -111, 1, 108, -69, 91, 31, -114, -123, 113, 48, 96, -83, 69, 11, 12, -16, 109, -13, 12, -34, -21, 110, 112, -23, -80, -88, 2, 38, 84, 92, 19, 70, -110, 98, -9, -89, 95, 33, -57, -38, -77, -88, -79, -127, -121, -116, -63, -114, 34, -23, -100, -64, -2, 14, 92, 88, -101, 75, -91, -46, -12, 104, 39, -114, 62, 83, 45, -46, 15, -26, 17, -52, 77, -49, 93, 23, -46, -42, 1, -27, -82, -125, 119, 127, 99, 85, 101, -11, -50, 62, -89, -98, -15, -23, 66, 69, -24, -98, 122, 1, -56, -88, -83, -105, 62, -85, 117, 67, -47, -125, 83, -50, -128, -23, 19, 28, 107, 73, 73, 121, 116, -109, 11, -3, -84, -9, -47, 101, 110, -23, 68, -15, -14, 54, 24, -37, -30, -26, -4, -102, 105, 49, 108, 46, 57, 75, -91, 40, 86, 9, -1, 8, 18, 34, -72, 102, 96, 97, 68, 77, -32, -61, 90, 122, 122, -67, -87, 61, 78, 81, 122, 63, -28, -113, -14, 30, -8, 79, 3, 92, 76, 12, -47, -98, -112, -25, 83, 64, 127, 91, 28, 35, 127, 23, -51, 78, -118, -52, 91, -127, 80, 65, 85, -62, -25, -108, 16, 9, 65, 65, 10, 68, -107, 41, 85, 16, 24, -68, -86, -71, 120, 81, -73, 32, 90, 67, 125, -120, -9, 105, 27, 2, 104, -41, 109, 9, 83, 126, -57, 89, -108, 61, -56, 67, 125, 73, 96, 114, -79, 104, -51, 33, -85, 82, -64, 105, 62, -104, 9, 97, -77, -110, -80, -107, 31, 3, 13, -25, 62, -56, 110, -35, 19, 84, -81, -5, 80, 8, -20, 94, 59, -117, 43, -67, 110, 43, 112, -108, 109, 90, -109, -114, -48, -60, 64, 4, -92, 8, -53, -114, -24, 14, 31, -37, -117, 112, 99, 81, 22, 98, -82, -13, 115, -122, 18, 99, -85, -31, 19, 39, 90, -29, -66, -34, 50, -103, 125, 34, -87, -80, -81, 67, -41, -25, 19, 1, 123, 102, 50, 53, 66, -111, 78, 8, 110, 67, 39, 98, -118, 114, -62, 48, 19, -55, 4, 41, -94, 62, 64, -56, -32, 95, 53, -111, -87, -8, 3, -54, 10, 13, 103, 63, 40, 109, 31, 30, -96, 64, -21, 16, -23, 0, -65, 19, -114, -115, 112, 57, -128, -63, 74, -87, -125, -117, -94, -8, 95, 46, 37, 12, 81, -109, -9, -102, -58, -87, 8, -83, -11, -74, 11, -66, -26, 57, 64, -66, 82, 91, 40, -18, 83, -57, -9, 44, -92, -75, 85, 36, 84, 36, 44, 78, -46, -89, -2, 87, 18, 89, -101, -111, -93, 117, -103, 105, -20, -23, -8, 54, -57, 79, 97, -112, -29, 27, -53, 12, -105, -82, -100, 72, 46, 10, 92, -91, 48, -47, -52, 81, -33, 8, 76, -45, 111, -29, 48, -36, -8, 105, 51, -15, 105, -113, 71, -25, 51, -68, -91, -52, 53, 50, -72, -115, -4, -109, -32, -99, -112, 77, 102, 107, -75, -83, -28, 16, 39, -92, -25, -48, -104, 88, -83, -65, 22, -98, 31, 122, -116, 103, -63, 13, -29, -55, -46, 105, -15, 73, 101, 59, 114, -49, -50, 95, 122, -63, -116, -76, 90, 62, 6, -45, 9, 102, 65, 46, 26, 29, 124, 87, -75, 85, 69, 94, 83, -106, -5, -27, 29, -114, 118, -88, 17, -109, 99, 76, 41, 30, 91, -59, -122, -90, -99, 58, 121, 10, -86, -106, 24, 119, 48, 92, 116, -93, 49, -64, -100, -68, 31, -18, -22, -20, -57, 74, 32, 115, -62, -111, -11, -110, -49, -81, -120, 56, -50, 92, -60, 21, -127, 7, -87, 93, -31, -54, 4, 50, -96, -44, 79, -85, 1, 79, 107, -125, 44, -113, 26, -33, 23, -125, 91, 117, 15, 74, 102, -90, -97, -86, -7, 0, -114, -1, 64, -106, -44, -13, 48, -33, 90, 68, -80, -120, 32, -63, -93, 107, -12, 110, -100, -32, 47, 21, -115, -81, 97, -104, -118, 55, 51, 10, 111, 95, -69, -108, -69, 47, -47, -28, -23, -49, 50, 116, -47, 94, -78, -110, -56, 57, -36, -83, -54, 106, -79, -71, 74, -100, -92, -5, 110, 0, 0, 68, 4, 73, -3, 55, -15, 0, -78, -37, 119, 125, 77, -124, -11, 89, -80, -67, -93, -35, -54, -81, 92, 4, 32, -75, -99, -111, 102, -43, -59, 47, -84, -80, 61, 98, -69, 50, 11, -19, -127, 118, 81, 41, -34, -52, 31, -69, -30, 97, 86, -90, 57, -44, 36, -81, -126, -124, 123, 4, -110, 6, -83, -106, -121, 95, -82, 96, -69, -54, 11, 25, 125, -67, 82, -109, -6, 53, -1, 100, -78, -80, 98, -66, 6, -18, -68, 25, -19, -68, -51, 127, 89, -41, 69, 68, -88, 103, 27, 17, -93, -54, -97, -29, 56, 16, 45, 74, -112, -21, 79, -9, -109, -19, 122, 89, 115, -98, -127, 24, -49, 24, -84, -86, -70, -13, -107, 42, 91, -46, -41, -117, 111, 1, -68, 50, 105, 21, 71, 59, -115, -62, 101, 63, 29, -33, -71, -63, -102, -92, 18, -10, -88, 23, 20, -105, -32, -74, -75, -65, 55, -67, -18, -18, 70, 116, -95, 89, -105, 44, 59, 92, -24, 46, 104, 19, 60, 88, 49, 19, -39, 46, -72, 111, -94, 104, -108, 26, 99, 41, 98, -85, -64, -120, -78, -99, -71, -17, 25, 94, -38, 39, 25, -49, 59, -25, 39, -77, -29, 96, -35, -38, -92, -123, 1, -113, 121, 64, 118, -1, -128, 94, 7, 69, -92, 25, 94, 127, -29, 111, -33, -78, -95, -96, 61, 107, 118, 90, 91, 116, 120, -15, -121, -31, 62, -37, -64, -45, 61, 73, 83, 88, 0, -66, -43, -109, 35, 63, -57, 121, -63, -103, -72, -5, 110, 12, -50, 70, 41, -92, -21, -22, -60, -47, -108, 44, -8, -31, 123, 1, 66, -35, -73, -101, -3, -58, -58, 45, 72, -55, 119, 48, -81, -113, -115, -23, -22, 127, -65, 53, 70, -125, 47, 17, 94, -47, 12, -125, 43, 66, -4, -33, -26, -123, 9, 49, -117, -107, -123, 18, -97, 78, 46, -111, -36, -2, -116, -63, -91, -44, -54, 5, 26, -70, 75, -46, -59, 87, -66, -5, 107, -82, 126, -78, 21, -19, -29, 14, -8, -107, 117, 70, 97, -12, -16, -4, -25, -97, 94, 25, 45, -63, 108, 14, 20, -21, -54, 25, -45, 2, 5, -41, 28, 49, 71, -68, -40, -14, -8, 74, 67, 43, -63, -86, -22, -61, -93, 39, 46, -29, -75, -77, -79, 25, -65, -86, 107, 86, -28, -9, 55, 27, 3, -90, 37, 7, 120, -109, -110, 22, -1, 50, -30, -12, -89, -29, 18, -71, 71, 41, -126, 110, -12, 58, 12, 74, -77, -100, 111, -128, 105, -24, -93, 49, 123, -70, -104, 15, -59, -113, 116, -106, 87, -76, -10, 68, 56, -125, 99, 43, 67, 120, -24, -49, 23, 52, 113, 99, 21, -31, 54, -113, -54, 67, -92, -45, -54, 112, 88, -84, -48, -56, -98, -106, 46, -97, 29, -25, -20, -96, 67, 121, -80, 83, -81, -128, 112, -35, 5, -112, 86, 81, 5, -59, -18, 111, 53, -91, -116, -100, -70, 17, -59, 105, 94, 14, 33, -14, -105, -27, 22, -120, 108, -110, -128, 52, 86, -21, 56, 125, -14, 43, -117, -67, -13, -31, -2, -68, -112, 76, -54, -118, 114, -44, 82, -118, 91, 38, 117, -4, -86, 75, -49, 86, -107, 82, 113, -74, 97, 97, 19, -120, -46, 61, 91, 102, 94, -127, 0, 38, 45, -115, 110, 114, 80, 96, -52, 28, 3, -17, -52, 6, 10, 22, 19, -119, -128, 50, -125, 91, 10, 4, -50, -32, 64, 86, -60, 84, -1, 103, 111, -62, 61, 14, -125, -116, -103, 2, 38, 22, -106, -120, -128, -126, 67, -44, -98, -126, -106, -9, 40, -18, 70, 49, -94, -78, -85, 118, -120, -11, 30, 52, 60, 59, -81, 3, 103, 114, -31, -50, -82, 118, -82, 25, 84, 124, -41, -20, -107, 80, -125, 5, 90, -103, 98, -44, -26, -104, -113, 91, 34, 79, 100, 50, 27, -65, 86, 124, 91, 36, -43, -63, 66, -83, -1, 18, 45, -114, -86, 35, -116, -101, 20, 86, -115, 9, -84, -96, -81, 28, 83, 2, -14, -64, -15, 69, -22, -98, -55, -1, -26, -128, 81, 37, 20, -30, 103, 85, -69, -29, -30, 16, 23, -92, -53, 73, 91, 99, -75, -94, -53, -15, -73, -127, 83, 123, -110, -5, -45, -9, 15, -65, -88, -115, 61, -83, -96, 22, 39, -31, -126, -73, -83, 77, 38, 91, -124, -65, 41, 94, -78, -87, -7, -121, 60, 41, -14, 29, -123, -52, -84, -18, 6, 20, -97, -101, 116, -75, 26, -88, 49, 40, -26, 26, 49, -17, 38, 125, 62, 11, -10, -38, 76, -52, 72, 65, -83, -3, 62, 27, -21, 18, -48, 5, -32, -121, -20, -49, 48, 93, 22, 95, 95, 79, -29, -81, 87, 114, -5, 83, 35, -53, 64, -36, -117, -105, -52, -27, -109, -106, -82, 69, 69, 83, 34, 126, 10, 118, -53, -90, 55, -56, 95, -2, 59, -117, -112, -21, 5, 19, 0, 78, 38, 22, -58, 82, -117, -22, 40, 109, 18, 38, 30, -128, 17, 73, -93, 74, -78, -16, -72, -48, -12, -67, 107, -79, 47, 127, 84, -109, 67, 83, 108, 30, -81, -62, -2, -98, 97, -13, 14, 46, 9, -34, 68, -84, -81, 92, 31, -105, 125, 107, 94, 54, -62, -90, 7, 126, -48, -112, -28, 51, 41, -120, -18, -6, -102, 96, -102, 36, 5, 56, 28, 101, -122, 0, 11, -63, -114, -54, 69, -88, 62, -100, 113, -6, 40, 32, -120, 121, -86, 78, 41, -59, -103, -38, -65, 99, 25, 47, 105, -16, -98, 62, 53, 45, 42, -15, 39, -47, 77, -30, -19, -124, -82, 45, 99, 64, 1, -110, 55, 70, -60, 87, 23, 32, -35, -93, -51, -47, 84, -65, -45, -57, -88, -12, 77, -46, -112, -111, -84, -38, 36, -87, 90, -114, -70, -42, -37, -97, -78, -49, 19, 117, 107, 26, 118, 52, 38, 72, 110, 44, 100, -51, 110, 127, 83, -109, -26, 35, -8, 67, 8, -14, 41, 34, 15, -30, -60, 103, -89, 34, -81, 31, -95, 25, -105, 50, -112, -89, -53, 40, 68, 91, 4, 78, 30, -123, -111, 112, -74, -67, 75, -9, 24, -27, -9, 86, -122, 63, 88, 116, 85, 68, 75, -18, -21, 12, 13, 68, 21, -89, 105, 44, 11, 3, -17, -110, 88, 118, -54, 10, -76, 92, 36, -121, 65, -5, 15, 127, -88, 92, 22, 52, 13, -53, -60, -112, 107, 60, 13, -22, -27, 6, 11, 100, -58, 36, -112, -85, 72, -45, -52, 17, -2, -45, 89, -40, -5, -22, 43, -23, -97, -26, -49, 11, 10, -119, 45, -76, -85, -28, 119, -77, -90, -2, 80, 58, 78, 122, 29, 42, 16, -72, -104, -3, -63, -74, 38, -19, -81, 61, -18, 117, -71, 36, 10, -111, 35, 115, -86, -74, 57, -123, 81, 59, 16, 78, 67, 62, -80, 123, 12, -27, -20, 33, 100, 2, 60, 98, -9, 53, 121, 103, 28, 62, -83, -87, -91, -80, -16, -128, -104, 4, 26, 49, 19, -114, 109, -106, -69, -10, -100, 64, -8, -121, -123, 106, 90, 47, -104, 95, 52, 12, -68, -75, 126, -128, -48, -86, 63, -39, 70, -92, -27, -87, -119, 86, 116, -37, -25, 53, 10, -14, 106, -24, 8, -4, 45, -49, -36, 113, 125, -48, -12, -56, 8, -123, -71, 65, -8, 56, 127, 66, -18, 123, 64, 115, 107, 67, 1, 79, 65, -21, -54, 80, -124, -118, -107, -4, -124, -72, -10, 31, 2, -99, 54, -121, 10, 79, 75, 67, 95, -20, 121, -103, -41, -17, -15, -15, -44, 109, -60, 47, -68, -84, -7, -115, 54, 6, -91, -115, -60, 73, -111, -116, 19, -74, 73, 47, 14, -66, 40, -67, 90, 116, 50, -28, 78, 63, -13, -106, -54, -48, 0, 23, -110, 53, -63, -122, 89, -55, 92, -33, -7, 28, -2, -49, 58, 120, 69, -75, 109, 105, 76, 92, 7, -33, 26, -8, 95, 0, 21, -13, -118, -98, 7, 45, 101, 99, 61, -123, -70, -98, -53, 106, 5, 67, 16, -97, 52, -114, -94, 54, -6, 12, -127, -75, 123, 31, -22, 55, -41, 68, 57, 32, -104, -119, 104, -103, -118, -35, 12, -51, 38, -116, -57, 38, -24, 70, 19, -63, 87, -48, -106, 112, -112, -31, -40, 66, 26, -51, 52, -118, -51, -125, 75, -46, -114, -66, 38, -10, -8, 110, -123, -99, 9, 56, 0, -29, -48, 10, -32, -89, 79, -41, -58, -83, 33, 38, -111, 69, 51, -25, -10, -79, 62, 104, 36, -89, -102, -52, 73, 87, -29, -23, 45, 96, -16, 59, -87, -56, -100, 20, 48, 70, 44, -14, 25, 114, -123, 102, 49, 120, 11, -37, -45, 56, -109, -81, -12, -18, -19, 122, 111, 76, -49, 93, -95, -25, 52, -95, 40, -8, -117, -78, -110, 96, -91, 114, -59, 38, -113, -128, -55, -3, -10, -8, 11, -120, -123, 40, -77, -114, -101, -67, -100, -8, -102, 5, -64, -51, -57, 52, -42, -104, 25, -108, 126, 52, 36, 3, -126, -65, 97, 120, 94, 43, 109, 69, -111, -82, -30, 118, 36, -101, -48, 119, 110, 8, -1, -79, -35, -53, -105, -1, -85, 64, 1, -108, -68, -60, -86, -23, -6, -86, -80, -62, -121, 115, -18, 65, 107, -35, -55, -22, 61, -97, -111, -115, 18, -74, -49, 78, -47, 91, 92, 48, -47, -105, -48, 117, 16, -91, 123, 110, 108, -95, 52, 10, -96, -94, 86, 56, 66, 48, -35, 107, -6, -65, 90, -90, -45, -9, 100, 32, 124, 61, -8, -53, -5, 21, 14, -74, -107, 68, 113, -67, 36, -79, 20, -80, -67, -92, 37, 19, 5, -118, -95, 11, 74, 73, -122, 24, -114, -62, -2, -39, 36, 126, -14, 37, -12, 54, 21, -46, -37, 35, 88, 101, 28, 66, 35, 52, -116, -14, 23, 102, -21, -108, 16, -84, 14, 15, 65, -102, 125, 106, -48, 11, 34, -6, 81, -74, -128, 72, -66, 68, -43, -38, -18, -100, 26, 84, -29, -15, -10, 51, 51, 115, 54, 120, 17, 8, -115, -73, 30, 20, -90, -10, 103, -32, -74, 58, -5, -50, 14, 30, 77, -102, -61, -26, 82, -84, 101, -82, 108, 38, 127, -125, 22, -94, 56, -94, -115, -115, 36, 70, 59, -108, 46, -63, 71, -70, 71, -92, 115, -105, -94, 95, 71, -36, -67, 22, 54, -86, 127, -105, 28, -90, 18, -53, 56, 10, -10, 78, 99, 78, 0, -106, 22, 42, -92, -47, 24, 76, -67, -41, -3, -35, 60, 52, -35, -96, 41, -38, 106, -83, -14, 46, 121, 94, -26, 36, -57, 81, 98, -15, 107, 49, 12, -64, 60, 32, -10, 38, 73, -45, -64, -123, 38, -18, 87, 17, 112, 35, -14, 104, -126, -64, 85, 68, 56, -7, 103, -34, 46, 50, 122, -22, -27, -78, -55, -93, 114, 25, 87, -48, 6, -97, -92, -108, 9, 53, 36, 75, 107, -97, 32, 6, 122, -99, 114, -6, -37, -125, 50, 29, -50, 95, 111, 26, 13, -123, 51, 117, 14, 98, -70, -25, 112, -32, 117, -55, 124, 121, -112, 26, -37, -89, -81, -32, 40, -52, 100, -22, -36, 57, 33, 89, -104, 122, -46, -26, -91, 34, -110, 0, -100, 13, 67, 47, 73, -70, -78, -18, -61, -102, 77, -112, -39, 3, 90, -87, -109, -88, -87, -5, -4, -49, 55, 122, -86, -43, 17, -13, 11, -19, -65, -96, -60, 28, 120, 115, -47, 4, 18, -47, 70, -21, -73, -81, -100, -110, 41, -51, 77, 113, -118, -125, 102, -92, -87, 66, -47, 12, -112, 126, 105, -27, -38, -2, 46, 88, 43, -122, -126, 0, -125, -82, -128, -86, 83, -83, -62, -79, 34, 45, -40, 121, 65, -33, -4, 13, -90, 118, -55, -44, 13, 87, 102, -118, 50, -33, -6, -125, 72, 66, 67, -18, 35, 16, 116, -88, -87, -15, -87, -9, 101, -71, 56, 76, 99, 52, -117, 68, -23, -19, -26, -76, -96, 50, 72, 114, 57, -126, -72, 103, 104, -15, -50, -60, 0, 84, 15, -94, 34, -128, 120, -98, -22, -15, -22, -74, 93, -62, 85, 0, -107, 13, 79, 28, -70, -58, 105, -47, -65, 38, 20, -40, 124, 71, -19, -56, -83, 18, 90, 76, -41, 37, 25, -2, -58, -96, 8, 64, -98, 73, 13, 50, 97, 50, -118, -19, 46, -63, 12, -127, -23, 91, 50, 24, -16, 109, -102, 74, 30, 46, -19, -126, 78, 3, -10, 112, -107, -25, 122, 35, 32, 27, 84, 80, 1, -103, -33, -77, 20, 85, -97, -109, 44, 66, -118, -88, -123, 89, 72, -107, -76, -121, 67, 58, 22, -104, 70, -76, 87, -102, -7, -47, 39, 10, 123, 80, -119, 69, -28, 87, 57, -25, 28, 19, 80, -33, -112, 9, -30, -1, -49, 118, -19, -98, 112, 54, -82, 31, -93, 93, 53, 16, 38, 86, 14, 21, 13, 59, -109, -61, 58, -88, -89, -25, -84, 49, -117, -71, -127, -27, -90, 42, -8, 98, 85, -49, 70, -97, -98, -29, -55, 30, -105, -17, -15, 73, 115, -8, -97, -10, -8, 61, -51, 97, 88, 44, -17, -106, -23, 22, 102, -7, -71, 35, 86, -96, -81, 93, -112, -8, 79, 8, 48, 112, -60, 20, -18, -72, 124, 115, -40, 69, -90, 44, 98, -105, 96, 96, 98, -88, -100, 59, -36, 83, -2, -14, 123, 102, 33, -88, 2, -85, 39, -40, 74, 86, -75, -33, 60, -95, 84, -45, -105, -126, 29, 15, -105, 85, 75, 83, -61, 33, 76, 43, 121, 65, 66, 113, -67, 67, -26, -70, -65, 47, -83, 52, -32, -30, -26, 110, 68, 87, -44, 59, 68, 47, -25, 123, 65, -72, -90, 91, 89, -106, -33, 70, -78, -78, -117, -108, -26, 77, -21, -15, -31, -127, -18, 93, -39, 39, -30, -98, -91, 55, 116, 96, 52, 46, 120, -51, -128, 3, -16, -21, 36, -32, -44, -87, 69, 96, -16, -41, 93, -71, -88, 68, -23, -22, -88, 18, 43, -97, -73, -12, 8, -45, -37, -114, -28, 21, -93, -53, 22, 30, 72, 71, -41, 8, 115, 45, 113, 89, -34, -18, 102, -58, 51, 23, -59, -78, -117, -11, 109, 12, -102, 68, 120, -53, 2, -47, 93, -84, -56, 100, 117, -19, -37, -93, 110, -72, -18, -59, 27, 77, 115, 105, 79, -49, -4, -60, 89, -71, -116, -115, 7, 45, 9, 45, 4, -77, 38, -60, 26, -87, -116, 124, 67, 45, 52, 69, 36, 4, 64, 4, -70, 81, -94, 107, -51, 96, 17, -76, -44, 69, -34, 79, -11, 49, 109, -111, 75, -55, 57, -59, 25, 26, -47, 102, -111, -27, 47, -125, -66, 119, 96, -126, 44, 59, 119, 15, 124, -127, 32, -114, 0, 99, -122, 81, 11, -65, 62, -122, 19, 18, -53, 67, 43, 48, 99, 53, 59, 105, 108, -3, -84, 112, 50, -89, -108, -80, -47, -50, 53, 12, 13, -68, 64, 60, -75, -11, 38, 32, -90, 51, 29, 63, -122, 83, -22, -86, -11, -48, -67, 109, -113, -52, 8, 21, -71, 118, -83, 17, 49, 59, -108, 47, 49, -12, -80, 106, -64, -93, -61, -62, 78, 57, -114, 87, -47, 20, -113, 84, -91, -39, -69, 16, 0, -78, -89, 53, -81, 88, 100, -63, 56, 66, -94, 118, -65, 7, -102, 53, -8, 114, -54, 91, -25, 41, -23, -7, -111, -102, 68, 20, -119, -68, 1, -15, 44, -109, -28, -52, 113, -103, 5, 86, -121, -70, 25, 86, -51, 27, 25, -37, 106, -69, -17, -125, 3, 89, -126, -30, 20, 28, 33, 71, 25, -110, 109, -121, -108, 95, -62, -109, 22, 19, 98, 79, -51, -19, 105, 113, -43, -75, 59, -102, -74, 14, 124, -60, -88, 39, 105, 8, 90, -84, 67, -117, -68, -100, 12, -98, -23, -17, -49, 90, -77, 76, 76, 25, -19, -43, 121, 43, -40, -19, -123, 109, -24, 118, -112, 14, -115, 18, 70, 93, -6, 18, 6, -82, -49, 78, 65, 82, 127, 93, 105, -15, -94, -121, 82, -30, 84, -78, -52, -95, 78, 70, -59, -42, 117, -26, 35, -1, -28, -100, 86, -89, 67, -50, -48, 10, -9, -42, 6, -9, -107, -117, 111, 43, 32, 18, -14, -6, -11, -71, -92, -10, -49, 74, 51, 125, 42, 123, 37, -41, -63, -66, 4, 30, -90, -101, 119, -86, -123, 28, 78, -114, 118, 90, 8, 43, -1, -84, 18, 79, 7, -43, -11, 36, -21, -6, 28, -35, -97, -95, 18, 13, 71, -17, 53, 9, 34, 13, 73, 7, -11, -27, -68, -24, -28, -12, 2, 127, 47, 49, -46, -105, 19, -89, 41, -29, -106, 39, 40, -126, -111, 121, -115, -36, -124, 13, -64, 34, -109, -29, -86, 103, -98, -117, -7, -55, -89, 40, 67, -24, -122, -106, 38, -73, -95, -10, 108, 6, -97, -61, 97, 73, 63, 91, 102, -93, -84, -51, 58, 1, -110, -100, -29, -88, 66, -77, -25, 77, 65, 69, 31, 67, -47, 120, 85, -127, 119, -31, 64, -35, -111, -53, 119, 104, 118, -77, -2, 126, -8, 60, -85, 0, 100, -3, 115, -2, 78, -91, 100, 82, -75, -12, 11, -122, 123, 70, -57, -35, 80, 65, 0, -3, 26, -97, 111, -7, -43, 71, -92, -53, -108, 46, 98, 73, 112, 2, -38, 95, -127, 65, -31, -84, -109, -118, 31, 5, 70, 96, 25, 91, 88, 3, -41, -16, 109, -85, 96, 8, -124, -112, -27, 9, 36, -61, 90, 29, 8, 105, -115, -26, 76, -13, -114, 4, -11, -98, -31, 30, 40, -120, -82, -126, 61, 73, 126, 98, -62, -55, -17, -17, -71, -51, 105, 123, -76, -92, 109, 23, -89, -100, 90, 11, 64, 40, -103, -26, -14, 28, -59, -113, 54, -59, 103, 1, -121, 18, -18, -104, -43, 19, 60, -99, 28, 109, -73, 92, 115, 52, -5, -72, 118, 119, -19, 50, -106, 50, 75, 67, 117, 10, 99, -114, -42, 94, -114, 4, 18, -22, 14, -122, -111, 87, 118, 62, -69, -124, -84, -51, -88, 89, 87, 111, -53, -83, 105, -53, 82, -21, 49, 88, -96, 21, -87, 60, -29, -25, 59, -24, 6, -94, 24, 41, -84, -11, -7, -91, -8, -4, -56, 5, 65, -66, -29, 5, 18, -22, 43, 86, -53, 33, 84, -103, -40, -44, 92, -64, -41, -67, -44, 79, 54, 3, -64, 49, 15, -88, 74, -61, -97, 76, -74, -90, -65, -110, -64, -33, 120, 64, 87, -77, -125, -72, 17, -96, -72, 67, 103, 27, 72, 51, 65, -72, -30, 4, -19, -57, 32, -9, 114, -72, 26, 101, 2, 123, -91, -75, -8, 12, 36, 112, -57, -102, -16, 127, -94, 51, 16, 117, -58, 21, 79, 86, -60, 63, -86, -40, 104, 79, 71, 126, 57, -118, 36, 101, 62, -120, 28, 96, -42, 114, 20, 111, -112, -125, 23, -85, 29, -54, -99, -97, 89, -85, 25, -82, 124, -37, -56, -12, 115, -22, -107, -71, -113, 41, -126, -86, 100, 28, 12, -43, 104, -51, 113, -76, -24, 26, -95, -124, 69, 18, -20, -5, 36, 33, 11, 26, 102, 67, -113, 88, -34, 86, 48, 1, -95, -120, -21, 56, -79, 25, 24, 70, -14, 54, 62, 43, -50, -44, 89, -103, 20, -108, -90, 2, 8, -80, 84, -34, 92, -80, 115, -93, 30, 58, 53, -68, 56, -47, -65, 64, 36, 20, 59, -87, 68, -10, 47, 7, 109, 63, 122, 38, -39, 16, -117, 78, 39, 91, -73, -86, -42, 119, 73, 86, -111, 11, -117, 127, -53, -8, 44, -72, -101, -38, -9, -15, -84, 23, 55, -107, 39, 32, 37, 66, -35, -32, -100, 94, -15, 110, -100, -61, 23, 66, 45, 120, -101, 91, -75, 113, -103, -36, 101, -106, -125, 45, 121, -72, -30, -17, 31, -101, -66, 86, 113, -1, -23, 53, -89, -21, -93, 57, -20, -31, 51, 32, 5, 22, 86, -29, -107, 7, -8, 120, -38, 49, 21, 28, -98, -74, -34, -47, 54, -35, -83, 82, -97, 123, 62, 110, -6, -73, -52, 17, 52, -60, -120, -46, -90, -121, 58, 64, 103, -42, -48, 94, -57, -79, -25, -46, -6, 100, 4, -61, -96, -1, -71, 62, 1, 105, 77, -121, 61, 42, 89, -38, 66, -111, 37, 29, 20, 29, -109, -64, 16, -113, 36, 14, 79, -108, -82, -9, 3, 99, 109, -17, 62, -119, 81, -29, -32, -81, 121, 18, -41, -43, -74, 83, -49, -6, 80, 18, 69, -76, 83, 76, 3, -65, -3, 81, -42, -61, 14, 92, 58, -7, 37, 7, -99, 96, -122, 85, -74, -10, 32, -55, 40, -1, -40, -94, 114, 14, -66, -105, -74, -42, 43, 80, -88, -118, -43, -89, 7, 77, 127, 87, 73, -112, 110, 101, 67, 27, 40, 69, -4, -78, -67, -104, 104, 43, -34, 84, -23, 106, 46, -122, 97, -12, -51, -116, -82, 71, -52, -19, 22, -51, 56, -42, 85, -26, -82, 41, 17, -19, -33, -105, 108, -16, 15, -49, -64, -102, 100, 116, 40, 122, 124, 55, 67, -99, 80, -31, -90, 1, 27, 80, -105, 96, 103, -77, -84, 61, 43, 37, 80, -118, 110, 8, -106, 88, 59, -69, 46, 79, -114, -123, 56, 99, 67, -111, -45, 17, 67, 118, -61, 72, -89, -31, 64, -30, -65, 62, 57, 49, 73, -12, 35, 81, 12, -43, -89, -58, -105, 74, -45, -120, -89, 10, 107, 80, -32, -4, -3, 18, -26, -80, -46, 102, -116, 113, -36, -105, -92, 112, -48, 104, 17, 49, 116, 31, 101, 47, 20, 108, -35, 100, -86, -124, 48, 78, -118, -117, -18, -12, -41, 27, -92, 112, 124, -1, 56, -91, 21, -80, -27, -115, 40, 8, -71, -102, 50, 78, 99, -64, 72, 111, -46, 65, -75, 32, 52, 61, -6, -60, 109, 93, -99, -52, 69, 60, 39, -77, 120, 82, -81, 45, 1, -121, 31, 47, 113, 14, 126, -118, -72, -92, 11, -61, -6, 113, 18, 10, 33, -96, 13, 28, -74, -17, -74, 82, 39, 71, -116, -34, -24, -17, -51, -100, -99, -95, -111, 101, 9, -122, 64, -72, 127, 29, 105, 123, 20, 3, 20, 104, -120, 4, 108, -79, -110, 125, 90, -38, 82, 48, 4, 32, 116, 100, 50, 125, 98, -96, -84, -50, -107, 71, -46, 40, 85, 74, -45, -105, 91, -107, 40, 28, 70, 34, 73, 96, 68, 123, -112, 82, 87, 65, 115, 108, -111, -47, 67, 74, -23, 123, -13, -85, 66, -77, -13, -117, -69, 64, 39, 90, -118, -96, -95, 16, 24, 120, -101, -12, 44, 113, 91, -21, 126, 29, -60, 73, -73, -39, -110, 53, 40, 116, 49, 56, -35, 49, 102, -16, -99, 10, -3, 64, 24, 45, -103, 33, 83, -72, 23, -8, -96, -35, 115, -92, 21, 44, -22, -126, -47, 73, -37, -25, 75, -72, -95, -31, 65, -45, 109, 54, -118, -42, -107, -37, 90, 112, 82, -59, -96, -125, 72, -123, -74, 57, -112, -26, -25, -121, 31, 111, -79, -98, -111, 15, -92, 26, 0, 49, -36, -22, -116, 83, -1, -64, 110, 75, 126, 86, -91, 48, 48, 42, -35, -52, -75, 109, 22, 46, 16, 11, 50, -105, 4, 75, -95, -118, 37, 51, 108, 60, -77, 104, 12, 41, 32, -2, -64, -43, -13, 85, 62, -1, 109, -60, 92, 45, -32, -126, 7, 74, -77, 17, 68, -58, -117, -73, -57, 21, 70, -84, 65, 4, -76, -101, -7, -82, -85, 92, 40, 8, 13, -46, -12, 99, -60, 107, -45, -94, 64, -17, -110, -36, -10, 47, -57, 90, 98, -40, -79, -52, -57, 62, 4, -54, 62, -45, -17, -106, -91, -84, -50, 107, 100, -91, -46, -2, 14, 90, 79, 23, 76, -58, 107, -122, -114, 98, -79, 64, -123, -108, -6, 36, -43, -53, -116, -5, 126, 41, 47, -18, -70, 39, -118, 86, 111, 89, 75, 109, 99, -104, 71, 121, 87, 79, -88, -13, -92, 84, -75, -6, -52, 1, -72, 52, 10, 62, 68, -118, 76, -8, -30, -45, -49, -62, -53, -104, 12, -116, 39, 120, 42, -94, 0, -99, 32, -110, -10, -126, -113, 119, -33, -16, 20, -110, 57, -64, 53, -113, 64, 104, 88, 63, 36, -46, 44, 60, 43, 119, 37, 108, -37, -67, -38, -7, -31, 67, -9, -53, -24, -50, 121, 69, -71, 43, -66, -74, -51, -27, 95, 57, 31, -119, -99, 126, 103, 47, -10, 26, -125, -4, -46, 71, 69, 85, -118, -65, -18, -68, -117, 90, -26, 28, -36, 90, 111, 56, -68, 97, 51, -34, -103, 85, -65, -42, 116, 7, 30, -84, 12, -18, 21, 72, 43, 119, 26, 104, -24, -92, -98, 120, 99, -93, 30, -65, -18, 46, 70, -30, 48, -114, 124, 12, -4, 65, -115, -49, -124, 49, 25, -43, -9, 93, -6, -78, 24, -53, 71, 78, 81, -37, 32, 29, -11, 18, 21, -35, 72, -14, 26, 121, 18, -69, -97, 27, -56, -73, -88, 38, 85, -86, -38, 25, 91, -25, 99, -48, 5, -100, 51, -29, -126, 80, 68, -46, -89, 36, -20, -44, 95, -7, -118, 32, -65, -112, -62, -80, -14, -124, 47, 90, -115, -94, 53, -116, -49, -3, 70, 84, 89, 57, 0, 71, 73, 41, 20, 98, -115, -2, -118, 6, -58, 36, -104, -60, -37, 94, 15, -85, -37, -38, 73, 75, 97, -105, 97, -33, -115, 110, 81, 92, -59, -95, -56, 58, -126, 109, -85, -66, 55, 8, -101, 109, -126, 42, -95, -46, 90, -96, 69, 75, 81, 81, 14, -48, 65, 60, -98, 95, -34, 50, 15, -87, 78, 110, 125, 52, 117, 71, -121, 46, -72, -78, -66, -57, -109, 36, -68, 76, 122, 92, -30, -5, 90, 60, -39, -96, -127, -104, -61, -117, -30, -106, -117, 57, -100, 43, -113, -29, 127, -87, -117, -36, 50, -3, 58, 45, 5, 56, 37, 10, 13, 3, -93, 68, -19, -23, 94, 87, 55, -124, -36, 49, -120, 48, -56, -28, 75, 38, 118, -94, -17, 109, 103, -45, -82, 69, -103, 127, -12, -16, -47, -31, -2, -86, -21, 93, 24, 54, -64, -90, -74, -105, -91, -70, -14, -93, -2, 56, 11, 105, 111, 48, 61, 121, 90, 48, 13, 9, -89, -11, 66, -127, -30, 11, 44, -24, 7, -4, 121, 101, 21, 114, 75, 94, 72, -82, 35, 93, -2, -27, -36, -103, -113, 55, -27, -120, 68, 104, 20, 3, 63, 36, -86, 82, -42, -58, 42, -17, 47, -111, 22, 37, -93, -61, -22, 77, -80, -16, 15, -57, -54, -37, 71, -83, -99, -66, 4, 43, 27, -128, 57, 14, 68, 14, -19, 80, -5, -9, 8, 65, -100, -85, -128, -33, -81, -79, 50, -91, -107, 89, 31, -90, 35, -7, -56, -21, -37, 60, 40, 119, 86, -79, -65, -87, 46, -8, -69, 23, 42, -123, -6, -45, 19, 28, 74, 117, 45, -24, -54, -127, -51, 12, 94, 92, 79, -95, -96, 49, 36, -12, -88, -57, -38, -5, 112, 26, -48, 9, 16, 40, -24, 83, -115, -55, -86, -12, -38, -44, 16, -90, -114, -90, -25, -109, -76, -83, -50, 42, 122, -116, 17, 17, 81, 77, 111, -54, 100, 67, -7, 121, -32, 49, 56, 59, 98, -49, 58, -85, -29, -29, 13, 58, 70, -63, -54, -96, 82, 19, 76, -60, -99, 28, -101, -28, 67, 111, -40, -62, 45, -102, -123, 33, -78, 47, 16, 13, 45, 78, 15, 10, -24, -125, -108, -2, 95, 7, -103, 13, -32, 37, -35, -48, -126, -126, -97, 30, -40, -51, 24, 48, 96, -112, 101, -127, -116, -47, 1, -5, -41, -18, 26, -110, 56, 21, -111, -91, 73, 57, -113, -21, -102, 75, -76, 55, -52, -71, 74, 104, 76, 14, -41, -24, -17, 103, -86, 46, -39, 114, 5, 104, 95, 27, 108, 52, 44, 108, 35, -48, 75, 13, 68, 42, 106, -41, 58, 56, -30, -21, 103, 122, 36, -13, -76, 79, 12, -107, -9, 7, -4, 105, -71, 72, 70, 83, -116, -42, -54, -79, 88, 43, 79, -112, -4, 36, -124, 19, 113, 4, 69, -42, 102, 31, -19, -48, -29, 29, 31, -22, 115, -10, 44, -20, -54, 2, 89, -29, 75, 59, 33, 93, -117, -13, 47, -109, -61, 11, -49, -98, -107, 80, 5, 57, -12, 34, 114, -81, 127, 68, 54, 30, 78, 91, -121, 8, -93, -62, -43, -89, 1, 70, -23, -16, -98, 60, -12, -109, 4, -11, -109, 114, 84, 110, 84, -119, 64, -83, -14, 119, 34, 109, 63, -55, -122, 62, -23, 96, 61, -72, 35, 4, -89, -36, 20, -72, -62, -17, -31, -119, 8, -17, -82, 55, -7, -30, 17, 83, -98, 28, 5, -120, 81, -37, -103, -81, -96, 26, 76, -103, 74, 37, -18, -125, 120, -71, -2, -22, 2, -74, -88, 88, -1, 118, 76, 50, 14, 58, 9, 19, -12, -119, 39, 38, -120, -5, -36, -117, 110, 28, -121, -25, -23, 87, 42, 58, 83, 76, 37, 100, -23, 32, -33, -118, -103, 97, 96, 70, 10, 36, 65, 23, 5, -70, 11, -60, 93, 9, -13, 26, 71, 80, -43, 82, -48, -63, 50, 44, 47, -119, -123, -105, -52, 34, -71, 49, -17, 112, -71, 56, 106, -75, 119, -85, -127, -42, 6, -124, 4, -111, -104, -1, 124, -41, -85, 21, -6, 101, -98, 109, -119, -58, -122, 86, -16, -75, -35, 127, 79, -7, -128, 22, -83, -23, -100, -26, -50, -111, -16, -85, -22, 86, -38, 43, -10, -75, -44, -3, 109, 58, 14, -18, 23, 106, 73, -105, -14, -100, -66, 124, 67, 29, -15, 105, -11, 60, -4, -46, 86, 41, -126, -122, 34, -34, -43, 27, 93, 14, -67, 49, -89, -24, 22, -71, 124, -31, 83, 117, 32, -104, -95, -35, -57, -83, -49, -127, 30, 85, -97, -100, 120, 62, -127, -37, -112, 89, -34, -9, -71, 10, -37, -17, 115, 102, -96, 99, -27, 110, 107, -78, -3, -121, -91, -42, 75, -72, 49, 6, -122, 6, -25, -29, 51, 0, 118, -90, -41, 101, -34, -16, 73, 28, -13, -116, 118, 73, 122, -5, -21, 48, -82, 98, 77, 41, 102, 26, -98, 122, -125, -76, -6, -94, 120, -64, -85, 0, 22, -22, 73, -62, -34, -94, -39, 36, -40, 20, 90, 121, -1, -29, -72, -16, 32, 27, 48, -19, 14, -110, 32, -55, 50, 18, -57, -109, -15, -13, -69, -79, 39, -87, 0, -128, -114, -53, -77, 104, -89, 102, 47, 4, -54, -126, -120, -122, 21, -91, 80, -106, -3, 70, 94, -23, 62, -92, -69, -31, -111, -92, -99, 42, 47, -6, -81, -50, -128, 86, -127, 100, 113, -3, 29, -39, 9, -116, 110, -92, 125, -64, -35, 114, 125, 94, -106, 7, -55, -21, -7, -58, 95, 78, -122, 44, 42, 25, 79, 35, -30, -11, 127, 115, -100, 106, 45, -84, -74, -47, -118, 23, -99, 0, -108, 46, 12, -109, -122, 29, -78, 66, 84, -69, 85, 22, 48, 27, 101, -117, 1, 14, 106, 35, 125, 86, -119, -5, 64, -44, -72, 5, 127, -65, 49, 89, -14, 22, 119, -120, -47, -128, -102, 122, 73, 93, 36, 37, 107, 92, 119, 37, -44, 96, -10, -70, 53, 94, -113, 121, 66, -89, -9, -64, -20, 6, 58, -127, -26, 84, -31, -23, 38, -90, -6, -60, -127, 47, 39, 96, 58, 4, -44, 68, -31, -96, 83, 14, 127, -60, 64, -74, -40, 42, 117, -65, -117, -63, 69, 93, -74, -28, -94, 56, -12, 107, 84, 56, -6, -9, -14, 55, 123, -17, -64, 121, -56, 48, 87, -117, -73, -45, -73, 48, -70, -6, -76, -45, -15, 79, -77, -47, -88, 112, 51, -47, -99, -95, -74, -11, 72, -29, -109, -77, 70, 30, -96, -97, 53, 115, 104, -80, -67, -3, 109, 88, 8, -106, 23, 27, -49, 77, -17, -82, -86, 19, -43, -125, 53, -23, 79, 88, -75, -49, -46, 100, -102, 104, -108, 28, -18, 121, -4, 57, -45, 38, -102, -18, -102, -46, 51, -109, -91, 37, 86, -128, -74, -11, 22, 79, -72, -27, -9, -72, 41, -34, 53, -31, -53, -123, -33, -58, 8, -13, 4, -66, 32, 7, -125, 15, -93, -93, -46, 22, 14, 43, 125, 120, 75, -123, 3, -92, 96, 68, 36, -32, -114, -7, -49, 117, -28, -3, 99, -37, 67, -72, -53, 33, -77, -94, -55, -33, -17, -77, 17, 11, -57, -56, 90, -41, -110, 75, -25, 65, -10, -90, 12, 63, -19, -51, -122, -54, -71, -127, -91, -51, 72, 116, 84, -98, 8, 24, 40, -85, 57, 1, -39, 18, 18, -26, 99, -15, -96, 103, -22, -78, -12, -14, -45, -61, 83, -121, -40, -24, -83, 79, 64, -48, -44, 48, -3, -11, -82, 115, -93, -127, -13, 17, -96, 126, -39, 37, 4, -84, -19, -66, -9, 81, -77, 19, 91, -53, -3, -62, 33, -47, -123, -41, -105, -81, 65, -93, 57, 23, 20, -33, 10, -104, -122, 29, 60, 9, -1, 54, 93, 34, -19, -75, -100, -120, -32, -47, 67, 98, 62, -127, -96, -84, 33, 32, 79, -4, -24, 49, 71, 124, -11, 60, 78, 48, -8, 60, -110, -123, -126, -78, 80, 46, 25, -30, 14, -94, 91, 103, 27, -106, -110, 71, 70, -55, 116, -25, 43, 5, -88, -98, 69, 104, 124, 64, -91, -119, -44, -107, 47, -67, 73, -8, 114, -106, 113, 75, -12, 27, 33, -84, 50, 97, -128, -5, -33, 11, -33, -23, 83, -29, 90, 99, -124, -70, -89, 8, -125, 60, -55, -99, -63, 65, 109, 33, 45, -118, -41, -58, 43, -65, -47, 72, 75, -2, 123, -54, 94, 99, -65, -48, -2, -72, 107, 50, 107, -68, 103, -88, 106, -62, -56, -51, -123, -105, 101, 81, 118, -2, -49, -5, -63, -49, 71, 80, -107, -24, -11, -34, -16, -25, 107, 122, 111, 66, -86, 71, 51, 82, 101, 18, -62, -63, -38, -110, 45, 3, -30, 18, 99, -123, 83, -78, 25, -52, -19, -90, -97, 84, -15, 96, -97, 119, 69, 15, 52, -38, 38, 71, -84, 47, -31, 29, 93, -67, -123, 75, 105, -2, 76, -19, 65, -8, -39, -5, -115, 14, -116, 24, 45, 25, -113, 96, -101, -47, -7, -85, 99, 110, -31, -112, -75, 111, -75, 70, -108, 94, 20, -53, 10, 16, 67, 4, -93, 68, -99, -120, -12, 119, -122, 120, -37, -35, -2, 115, -113, 63, 47, -111, -55, 90, -118, -60, 36, 19, 6, 77, 120, 62, 3, -53, -3, 78, -68, 42, 113, -28, -119, 4, 76, -99, -71, -19, 99, -76, -33, 38, -33, -20, -85, 124, 125, 16, 61, 81, -125, -2, 50, -24, -87, 93, 66, 91, 49, -61, 57, 74, 43, 85, -29, -105, -79, -10, 124, -26, -89, -45, 84, -59, 24, -40, -110, 111, 101, 24, -91, 91, 82, -9, 72, -79, 49, 75, 5, 105, 17, 19, -105, 117, -101, -114, 25, 72, 102, 114, -21, -72, -17, 59, 97, -62, -45, 8, 37, -65, -19, -13, -35, -124, -70, -44, -26, 113, 88, -105, -64, 94, 36, -42, -17, -63, -42, 117, 30, -58, 6, 90, 28, 84, -58, 46, 54, 98, 89, 46, 66, -91, -29, -111, 8, -61, 7, -80, -14, -1, -15, 111, -115, 59, 117, 83, -127, 113, -82, -23, -23, 18, 18, 107, 51, -78, 126, 41, 126, -118, -70, -22, -41, -2, 28, -46, 16, -48, 40, 93, 97, -48, 29, 83, -38, -35, 5, 37, -97, 64, 27, -60, 79, -8, -113, 71, 103, 36, -124, 113, -70, 59, -49, 80, -97, -113, -18, -88, 3, 110, 41, 13, -11, -4, 121, -50, -9, 47, 105, -10, -15, -86, -23, 87, -52, 57, 30, 113, -111, -99, -121, -101, 105, 63, 107, 126, -40, -92, 28, 5, 0, -52, -41, -90, -56, -34, -127, 85, 121, 64, -128, 41, 28, 75, 43, -28, 48, 38, -31, 27, 81, -71, 69, -59, -97, 113, 120, -105, -107, -60, -22, 85, -66, 118, -68, -11, -99, -128, -54, 72, -20, 110, 53, -93, -16, 53, 108, 9, 99, -83, 14, -39, 99, 113, 97, -97, -10, 119, 61, 13, 106, -52, 124, 123, -57, 9, -19, -54, 74, -61, -21, -113, -44, 13, 82, -1, 32, 93, 124, 60, -94, -115, 123, 77, -119, 81, 6, -32, 70, 114, 29, 53, 76, 109, 72, 36, -9, -48, 113, 9, 66, 2, -36, 71, 88, 0, -74, 14, -55, 95, 115, 42, 76, -118, 16, 32, 56, -11, 110, 19, 44, 45, 79, -53, 119, -68, -86, -97, -84, -114, -108, -45, 11, -99, 126, 83, -1, 37, 118, 47, 123, -128, 33, -13, -7, -75, -101, -8, 108, 39, 123, -118, 114, 46, -8, 74, -55, 51, 116, 70, 73, 112, 52, -95, -41, -99, -101, -53, -106, 96, -28, -70, 81, 100, 72, 58, 51, -73, 53, -94, -13, -116, 94, -125, 99, 7, 98, -41, -78, 3, -71, -98, 112, 12, -122, 64, 40, 19, 120, 56, 76, 22, -4, 80, -19, -10, 29, 118, 49, 59, -50, 67, 52, -72, 7, 76, -92, 77, 115, 76, -22, -34, 81, -115, -29, -113, 84, 96, -57, 9, 18, 123, -127, 86, -40, 14, -53, 91, -82, 19, -122, 15, 43, 24, -72, -13, -10, -16, -26, 21, 81, -13, -118, 76, 47, 123, -79, -44, 76, -67, 106, 29, -96, -97, -62, 29, -13, 49, -21, 104, 78, -77, -94, 14, -55, -69, -105, 81, 85, 8, 114, -27, 19, 110, -76, 72, -47, -105, -103, 47, 12, -59, -92, 72, -9, -112, 58, 6, 118, -106, -85, -37, -123, 66, -47, 15, -127, 68, 80, -115, 109, 11, -34, -78, -116, -44, -19, -50, 46, -56, 18, -25, -36, 7, -62, -25, 101, -79, 5, 118, 10, -46, 84, -87, 3, 10, 42, -32, -51, -51, -55, 108, -95, -20, 124, -58, -45, 43, -124, -68, -33, -5, -100, -124, -29, 2, -3, 124, -62, 11, -18, -70, -97, -111, -80, 72, -1, 0, 93, -6, 15, 91, -47, -80, -54, -34, 92, 116, 48, -108, -87, 10, -43, 127, 48, -21, -113, 30, 70, -3, 20, -101, 120, 73, -115, 11, 125, 113, -5, 26, -69, 109, -53, 50, -58, -41, -5, 76, 49, -114, 44, -99, -108, -16, 109, 92, 109, -33, 76, 22, 96, 9, -66, 30, 90, 19, 118, -66, 126, -39, 16, -10, 103, 91, 31, 127, -7, -127, -96, 118, -113, -103, 127, -70, 44, -74, -112, -42, 94, 38, -27, -108, -104, -114, 79, -106, -41, 7, 35, 124, -86, 78, -62, -117, 0, 113, -10, -71, -5, 95, -25, -18, -120, 55, 125, 28, -104, 60, -54, -89, -88, 55, 121, 54, 16, 64, -64, -11, -80, -33, -58, -58, -60, 100, -119, -77, -50, 10, -23, 41, 0, -111, 9, 19, -101, -93, 30, 1, -39, 65, 67, 93, 88, -3, -83, -81, -79, -102, 7, -62, -37, 122, 25, -7, -34, -66, 88, -47, 93, -58, -41, 98, 72, 118, 117, 115, -31, -115, -121, -64, -106, -70, 17, -65, -80, -29, -27, -54, 23, -110, 89, 39, 77, 73, -48, 40, -123, -81, 104, 111, 56, -99, 98, -107, 93, 68, -68, 44, -25, 56, -95, 4, 79, -53, -3, -106, -42, 42, 116, 56, -81, 125, 118, -40, 41, -68, 43, -30, 111, 43, 43, 120, 120, -85, 117, -48, -53, 93, -97, 103, -49, 92, -74, 68, -27, -68, 18, -75, -7, 109, -27, -35, 41, 45, 7, -21, -78, 30, -41, -16, -14, 115, 32, 112, -30, 58, 17, -3, 111, 47, 124, -9, -24, 116, -14, -120, -103, -28, -86, 25, 29, 127, -19, 57, -65, -127, 101, -67, -110, -125, 83, 52, 127, 103, -80, 76, -101, -122, 32, 32, -86, -109, 81, -72, 4, -46, 104, 76, 0, -48, 45, -43, 99, -118, -67, 110, -18, 59, 51, 47, -63, -108, -65, -58, 121, -123, 58, -7, 99, -112, -49, 55, 81, -77, -27, 106, -52, 88, 94, -84, 109, -9, 58, -91, -127, -22, 12, -6, 84, 11, -69, 55, -77, -113, 95, 110, 5, -119, 55, -4, 28, 117, 101, 3, -59, 99, 112, -53, -33, 22, 74, 41, -97, 35, -30, 122, -118, -48, 123, 18, 122, -109, -8, 94, -117, -109, -51, -32, 110, -118, 102, 13, -39, 59, 3, 30, -51, -88, -111, -118, 34, -86, 51, 108, -74, -97, -67, -121, 60, 81, -71, -12, -121, -30, 18, -105, 49, -128, -4, 25, -83, -42, 26, -68, 108, -71, -2, -62, 55, -90, 2, 15, -105, -112, -86, 77, -112, 48, 98, -33, -4, 101, 12, -52, 66, -6, 108, 102, -53, 36, 4, 40, 36, 111, -25, -10, 42, 68, 26, 7, 91, 56, -104, -6, -29, 47, -114, -107, 100, 23, 46, -22, -71, 0, -75, -67, -22, 7, -10, -7, -63, 12, 100, -38, 30, -88, 5, 25, 30, 7, 115, 32, -24, 25, 90, 121, 19, -26, -112, -16, 62, -112, 98, -101, -121, 123, 85, -100, -27, -115, -95, -128, 35, -116, 50, 63, 66, -39, 15, 33, -7, -2, 84, 94, -23, 23, 71, -80, -27, 93, 6, -10, -2, -7, 27, 51, -114, 96, 79, -30, 70, -81, -25, 71, -119, 45, -78, -42, -73, -100, 35, 54, -19, -54, 33, -119, -109, -127, -51, 115, -20, 38, 94, 32, -120, -90, 73, -17, 11, -85, 121, 14, -93, -55, 68, 126, -90, -99, 47, 20, -93, -39, -73, 70, -21, -18, -90, 18, 43, 87, -60, -56, -5, 40, -16, 103, 8, -13, -6, 116, 69, -45, 127, -52, 6, 87, 113, 4, 43, 125, 63, -101, -36, -99, -6, 16, 0, 59, 94, 106, 41, 121, 117, 73, 70, 24, 115, -99, 65, 89, 25, 49, -28, 65, 12, 33, -125, 13, 85, -113, -48, 82, 46, -13, 51, -88, -85, -40, -40, -3, -121, -65, 75, 39, -58, 42, -127, -16, -13, -24, 21, 81, 78, 60, 83, -64, -35, 96, -71, -119, 27, 126, -15, -102, -55, -16, 95, 51, -40, -49, -114, -2, 18, -11, -104, 115, -123, 58, -53, 73, -30, 4, 94, 5, 65, -77, 104, 103, 10, -103, 35, -28, 90, 47, 19, 7, -70, -98, -63, -107, 27, -79, 80, -87, 23, -125, -19, -80, -57, -114, -101, 97, -41, 83, 12, -33, 27, 55, 45, -115, 65, -78, -108, -34, -29, 17, -28, -36, -55, 54, -36, -6, -57, 16, 65, 36, 32, 123, 15, 104, -115, 111, 78, 101, -95, -45, 126, -63, 56, -4, -20, 1, 25, 53, 38, 89, 48, 107, -44, 44, -93, 55, 124, 1, -10, -52, 116, 41, -78, -115, -60, 10, -96, 19, 12, 93, -40, -115, -77, -20, 105, 46, 108, 50, -124, 124, 81, 114, 127, -11, 52, 118, -112, -32, -39, 83, -107, -29, 83, -25, 99, -13, 47, 94, 68, 21, -25, 86, 78, -93, 91, -47, -106, -80, 119, -6, -51, 104, -12, 18, -71, 5, -23, -70, 12, -88, -115, 101, -127, -33, 125, -112, -13, 125, -1, -120, -105, 66, -92, -57, -71, -26, -109, 95, 72, 123, 12, 15, 58, 51, -103, 45, 122, 87, 51, -116, 1, -59, 58, -6, -51, 80, 36, -65, 15, -2, 122, 107, 47, 59, 71, -67, 28, 74, 15, -93, 11, -4, 13, 43, 60, 2, 52, -90, 100, -29, 26, -36, -76, -48, 89, -90, -86, -20, -69, 52, -3, 9, -53, -103, 107, -28, 80, 61, 74, 20, 23, -70, -20, -28, -8, -119, 40, -47, -79, -112, -32, -53, -73, -31, 72, -113, 23, 81, -53, -62, 62, 42, 1, -35, 21, 83, 88, -87, -49, 55, 40, 102, 120, 14, -50, 3, -119, -121, -120, 16, 82, -66, -8, -27, 99, 28, 7, -20, 76, 53, 120, 19, 67, -4, 6, 5, -19, 27, 96, -33, 54, 108, 50, -62, -113, 94, -41, 115, 119, -82, 62, 32, 118, 38, -8, 88, -120, 50, -65, 11, 58, -64, -73, -31, 36, -67, 77, -121, -93, -25, -28, 66, -71, -90, -51, -118, -36, 16, 66, -121, 54, 97, -119, 124, -2, -124, 16, 91, 2, 104, -22, 32, -16, -51, -71, -89, 123, 61, -112, 107, 107, -78, 18, -76, 65, 123, 121, -44, -91, -43, -107, -94, 102, 91, 71, -46, -63, 87, -84, -20, 112, -43, -37, -41, -67, -4, -104, 121, 4, -47, 95, -6, -4, 66, 114, 84, -68, 77, -94, -68, -37, 47, -112, -86, 102, -24, -51, -127, -34, -42, -57, 80, 31, 41, 62, 27, -22, 95, -81, -78, 9, -94, -26, -14, -13, -112, -7, -81, -33, -59, 16, 112, -18, -101, -67, 11, -33, -66, -83, -120, -60, -4, 79, -65, 37, -29, 11, -74, -59, -121, 124, -64, -68, 105, -96, -16, -70, -108, 79, -16, -24, 62, 16, -115, -83, 14, -20, 92, -37, 91, 13, 14, 20, -113, 89, -6, -90, -26, -89, -48, 79, -11, 61, 27, 81, -58, -106, -88, 114, 48, -82, -68, 74, -24, -112, 20, 104, 66, 51, 120, -119, 10, -42, 1, -93, -22, -94, 54, -65, 45, 11, -5, -93, 104, -16, 49, -125, 76, -80, 80, -109, -80, 40, 87, -64, 127, -108, 31, 56, 54, 24, -64, -72, -86, 81, -51, 99, 97, 101, 47, -98, 103, -46, -52, -6, 54, -99, -52, -86, -13, 33, -34, -82, 22, 78, 56, -58, 70, -40, -19, -116, -118, 82, 14, 16, 91, 1, 5, 22, 0, -107, -109, 54, 58, -78, 72, 23, 87, 29, -119, 122, -102, 111, 119, 90, -106, -125, -40, -80, 95, 9, -32, 80, 52, -79, 46, 109, 101, -13, 65, 87, 54, 53, 98, 100, 75, -57, -39, -5, -92, 30, 73, -63, -69, 127, 30, 104, -45, 11, 106, -45, 52, -34, 27, -31, -103, -56, 53, 92, -20, -11, 37, 15, 25, 116, 78, -1, 88, 76, -25, -108, -93, 36, 40, 35, -101, -6, 83, 92, 56, -119, 0, 19, 9, -33, -10, 63, -56, -79, 1, 60, -64, 105, -48, 113, -37, 0, 76, -89, 24, 112, 25, -125, -76, 49, 120, -52, -50, 20, 51, 21, 98, -24, 73, 119, -73, 20, -76, -41, -109, 115, 103, 34, -60, 5, 84, 36, -21, 6, -109, -82, -91, -78, -27, 123, -25, 94, -116, -67, 121, -72, 100, 122, -94, 83, -67, 7, 67, 97, -20, 42, 124, -8, 13, 69, -77, -119, -84, 41, 53, 61, 5, -101, -21, 43, -62, -93, 66, -108, -63, -110, 77, -12, 0, -27, -54, 86, 18, 112, -41, 95, 72, 38, 86, 52, -75, -97, 3, 54, 121, 32, -43, -70, -124, 90, 30, 80, 91, -12, 112, 74, 22, 122, -89, 61, -57, 31, -86, -123, -110, 79, 15, 92, -110, -96, -82, 15, -122, -67, -62, -54, -36, 25, 66, 105, 13, 91, -21, 69, 11, -69, -11, 35, 10, 72, -13, 91, -51, -37, 48, 113, -4, -49, -39, -44, -114, 92, 50, -74, -73, 21, -72, 6, 73, 117, -121, -40, -35, -42, -70, -51, 91, -106, -121, -42, -29, -114, -93, -9, 51, -95, -22, -117, 81, -35, -15, 118, -41, -39, 93, 117, -17, -80, 115, 66, -68, 100, 50, -25, -81, 119, -50, -93, 3, -53, 12, 113, -37, 16, -91, 59, 31, -32, 54, 57, -3, 2, -73, -16, -118, 73, -118, -14, 66, 2, -75, -56, 49, -70, -78, -23, 8, 31, 57, 53, 30, 28, 80, 47, -8, -31, -66, -26, 102, -52, 24, 4, -49, -52, -102, -111, -77, -116, -81, 112, 0, -88, -63, 103, -47, -22, 55, -70, -7, 117, 23, 21, 14, -47, 51, 4, -52, -11, -58, 5, 33, 59, -51, 55, 16, 2, -15, 75, -17, -85, -112, -125, 60, -97, 79, -37, 90, -79, 101, 73, -28, -51, 120, -12, 49, 54, -60, -29, -39, 65, -128, 19, -97, -3, -71, -39, -99, -21, -41, -3, 77, 108, 53, 53, -86, 84, -44, 55, -26, 33, -51, -54, -77, 24, -59, 34, -125, -68, -86, -83, 10, 73, -64, 111, 106, 45, 105, -126, -18, -10, -103, 87, -103, -106, -76, -104, -31, 63, 94, -98, 28, 36, 54, 85, -40, 125, 51, -78, 8, 74, 79, -16, 37, -6, 66, 76, -51, -31, -99, -11, 110, 82, 53, -55, -122, -100, -107, -52, 96, -16, 113, -74, -87, 96, 38, 123, -9, 28, 28, 6, 38, -99, -80, 72, -81, 18, 47, 116, -123, 92, 90, -15, 100, 10, 36, 59, 19, -97, 50, -106, 31, 50, 12, 79, 15, 57, 41, -79, 37, -74, -10, 13, -71, -27, -74, -82, 117, -53, -64, 59, -107, -67, -122, -36, -77, -72, 44, 13, 125, -23, 38, 14, 46, 51, 86, -33, -127, 27, 96, -123, 57, -43, -112, -53, 42, -102, 93, 116, 54, -69, -70, -85, -8, -88, 10, -43, 51, 1, 11, -112, -83, 30, -79, 32, 76, 119, -41, -41, -85, -95, 120, -119, 123, -115, -68, -21, 39, 45, 65, -58, -116, 100, 44, -1, 97, 102, -34, 54, -33, -29, 66, -48, -76, -16, -90, -26, 41, -68, 119, 14, -63, -53, 77, -23, -120, 63, -28, -67, 79, -109, 1, 123, -34, 50, 52, 21, 23, 122, -126, 33, -40, -79, -5, -96, 6, -95, 30, -127, -36, 82, -26, 41, 32, -81, -11, 37, 69, 95, 38, 120, 5, -81, 99, -120, 45, 123, 90, -54, 41, -16, -6, -22, 122, 23, -77, -27, -68, -82, 99, 17, -10, 32, -84, 73, -10, 114, 90, 112, -121, -65, -14, 103, 65, 29, -101, -83, 35, -128, 68, -57, 107, 111, -79, 51, -104, -99, 62, -27, -46, 7, -25, -49, -65, 110, 106, 91, 80, -119, 105, -86, 84, 113, -99, -9, 71, -114, -34, 125, 101, 65, 37, 26, -84, -25, 89, -76, -27, 43, 33, 38, -114, -106, -42, -29, 110, 77, 63, -97, 121, -101, -79, 49, -72, -74, 82, 47, 24, -23, -58, -86, 114, -46, -65, 44, 89, -77, 96, -40, 49, -108, 112, 104, 113, -78, 67, -98, -25, 67, -105, -95, 29, 65, -68, -42, -24, -81, -60, -101, 71, 50, 100, 90, 63, 39, -100, -118, 19, 9, -62, -128, -6, -51, -84, -76, 115, 53, -39, -63, -17, 86, 100, 85, 86, -69, -64, -74, -99, 120, -2, -107, 10, 115, 39, -51, 50, 124, -67, -126, -106, 62, -39, -71, 48, -92, -50, 56, -94, 14, -45, 103, 18, 102, -16, -123, -78, -58, -109, 108, -69, -110, 2, 82, -72, -100, 120, -73, 79, -3, -2, 12, 114, -85, 72, 52, -98, -82, -87, 95, 28, -37, -100, -27, 91, -57, -118, -110, -111, -125, -14, -33, -96, 79, -89, 21, -13, 99, 115, -7, 108, 29, -112, -109, 14, 104, 37, -37, -51, 60, 68, -55, -62, -127, -118, 46, 16, -57, 12, 68, -66, 7, -114, -46, 119, -49, -40, 69, 88, 111, -116, 66, 100, -43, 59, -126, -125, 96, -68, 102, 117, -105, 88, 103, -45, -120, -109, -7, 38, -118, 81, 56, -102, -64, -34, 122, 9, -39, -8, 108, -109, -114, 67, 69, -51, 116, 42, -25, 101, 21, 24, -116, 63, -112, -65, -5, 47, 96, -71, -78, 88, -79, 123, 55, 94, -108, -122, 26, 20, -11, 69, 49, 67, 46, -122, -110, 104, -107, -89, 60, -92, 3, -112, -114, 26, -65, -20, 75, 20, -40, -75, -57, -57, -114, -53, -12, 16, 116, 44, -50, 99, 66, 1, 8, -125, -104, -20, -81, 95, 106, 61, -104, -37, -95, 114, -63, -109, -46, -18, -112, 33, 125, -12, 113, -48, -12, -81, 59, 22, -98, -13, -34, 117, -117, -50, 22, 20, -91, -70, -52, 22, -55, -107, -71, 66, 82, -59, -85, -40, 95, 76, 119, 70, 24, -115, 70, -57, -84, -103, 24, 95, -121, -36, 5, 70, -119, -63, 59, -61, -13, -47, -43, 17, -128, 96, -27, 59, -44, -99, 12, -43, -51, 91, 86, -6, -93, 116, 75, 77, 95, 87, 92, 40, 117, 58, 81, 68, -91, -57, 54, -18, -72, 76, 109, 108, 42, -51, 80, 40, -74, -24, -101, -6, 30, 25, -37, -71, -44, 60, 20, 19, -78, -59, 94, -128, 24, -32, -9, 118, 27, -58, 91, 91, 9, -37, 113, -128, -107, 20, -81, 98, -100, -63, -113, 113, -53, 35, -12, 16, 87, 68, -7, -81, -75, -85, -25, 63, -95, 47, -68, -29, -68, -113, 64, 70, -67, 51, 17, -35, -6, 77, 19, -40, -12, -6, -32, 72, -1, -122, 15, 110, 77, -42, 57, -2, -99, 99, -35, -23, -93, 26, 85, -49, 62, -117, -69, 107, -66, -103, 65, 110, -19, -53, 10, 97, 39, -91, 94, 47, -116, 76, 54, 115, 31, -122, -77, 30, 38, 22, -39, -33, -118, 51, 16, -19, -126, -3, -124, 120, 76, 124, -92, 47, 5, 102, -20, -124, -33, 21, -61, -30, -7, 47, 83, 53, 61, -48, 10, -67, 122, 0, -118, 14, -85, 2, -65, -47, 46, 113, 17, -89, -53, -65, 45, 74, 123, 92, -80, -116, -101, 33, 89, 68, 105, 78, 11, 93, -82, 102, -58, -19, -75, 13, 73, 6, 8, 102, -23, 67, -78, -48, -85, 63, 124, 78, 56, 41, 69, -101, 68, -98, -41, 17, 54, -18, -99, 121, 80, -7, -51, -116, 8, -91, -73, -33, -35, -10, -46, 81, 61, -75, -103, -9, 19, 1, -95, -122, 35, 60, -98, 13, -45, -86, -95, -109, 59, 9, 107, -66, -88, 14, 49, 106, 101, 48, 104, -118, 8, -68, -9, -91, -79, -107, -128, -40, -93, 66, 115, -4, -86, 13, -114, -103, -9, -108, 50, 11, 21, 52, -46, 45, 27, 12, 125, 25, 36, 123, -12, 63, 65, 10, -6, 108, -31, 71, -25, 12, 10, -64, -56, 110, 10, -14, 57, -100, -83, 26, 16, 115, -14, -23, -12, 28, -100, -103, -88, 106, 95, -107, -126, 103, -44, 110, -51, 69, 98, -113, -83, 33, -27, 81, 125, 23, -33, -13, -95, -55, -54, 60, -111, -87, 127, -17, -33, 114, -26, -25, -59, 14, 109, 72, -74, -31, 67, -85, 125, -75, 15, -24, -56, -109, -45, 104, -71, -92, 85, 62, 12, -105, 102, 70, -103, 93, 25, 125, 44, -62, -115, 118, 11, 60, 59, -66, -85, 64, -123, 26, 0, -36, -59, -117, 123, 59, 124, 115, -71, 119, -112, -94, 72, -101, -31, -122, -8, -20, 47, 106, 115, -34, 53, -61, 69, -95, 104, -4, 101, 24, 38, 116, -73, -112, -120, -104, -62, -10, 78, -77, -42, 87, 123, -88, -26, 62, -30, 54, 25, -86, -24, -95, -92, 46, -53, -18, -34, -9, 83, 69, -97, -104, -70, -77, 44, 34, 118, -107, -67, -37, -101, -78, -18, -81, 88, 115, 12, -61, -13, -12, -89, -116, -73, 52, -97, -114, 66, 25, -11, -71, -12, -87, -115, 27, -90, -54, -123, 24, 49, -15, -37, 66, -36, 71, 1, -57, 13, 6, -92, -23, -92, 98, -35, -115, 77, 40, 39, 81, -36, -109, 108, 110, -7, -2, -4, -27, 11, 48, -108, -64, 126, -35, -67, -87, 4, -121, 98, 116, -126, 105, 18, 106, -8, 79, 44, 88, -72, 30, 9, 80, 46, -23, -74, -88, -126, 50, 23, 1, -77, -101, -79, -91, 61, -76, 66, 84, -43, -18, 6, 63, 64, 34, 117, 79, 96, -11, 24, -82, -127, -2, -106, -42, 44, -24, 56, 126, -114, 44, 78, -53, 121, -55, 10, 121, -105, 84, 25, -75, 72, -33, -122, 41, -68, 12, -35, -99, 122, 61, -24, 3, 64, -54, -75, 59, -94, -33, 59, 118, -30, -90, 55, -28, -110, -112, -62, 103, 108, -104, 89, -45, 122, 70, 54, 79, 103, -25, -20, -101, -71, -67, 91, -5, -48, -11, 104, -112, -111, 15, 38, 38, 60, -26, 89, -78, -109, 48, 80, 55, -21, -35, -57, -50, -88, 19, 70, -56, 24, 70, 29, -69, -85, -25, 100, -22, 122, 94, -6, 127, 50, -18, 64, -75, -48, -77, 105, 8, -38, 88, -84, -51, 4, -35, 85, 84, 73, 96, 3, -55, 45, -119, 111, -58, 6, -24, -53, -49, -39, -83, 105, -109, -3, -44, 79, 86, -68, 62, -110, -22, 37, -25, -101, 11, 5, 67, 25, 40, -52, -7, 10, -73, 126, 61, -103, 67, -125, -43, 109, -53, -38, 8, -59, -4, -20, -65, 11, 16, -102, 70, 43, 83, 56, 117, 31, 127, -103, -80, 121, 28, -63, 65, 0, 75, 80, -31, -98, -31, 112, 108, 90, -30, -51, -72, 15, -35, -108, 71, 79, 19, 18, -85, -42, -7, 1, 108, -16, 7, -63, 13, 67, -69, 12, 68, 112, -56, 68, -125, 78, 125, -21, -31, 45, 103, 114, -84, 74, 40, -111, -63, 0, 39, -46, -41, 117, 90, 43, 120, -17, -75, 68, 113, 97, -42, 75, -77, -45, -114, 65, -6, 110, 28, -55, 21, -75, -113, -40, 38, 35, -67, -3, -14, 50, -125, 79, -55, 65, 110, -29, 25, -9, -8, 109, 106, 105, 119, -103, 13, -35, 16, 56, -29, -57, 119, -73, 103, 123, -65, -118, -126, 12, -42, -50, -126, -122, -28, 54, 91, -109, -32, 34, -50, -40, 19, 3, -87, -44, -7, 119, -16, 48, 98, 33, 33, 1, -68, 101, 87, -39, 83, -122, -78, 8, 66, 54, 54, 99, -92, 89, -18, 113, -3, -58, -61, 33, -70, -128, 99, 27, 5, 39, -65, 53, 71, 43, 21, -4, 30, -109, 37, 84, -49, 39, 36, -99, -92, 73, 19, -13, 34, 71, 119, -66, 92, -89, -111, -68, -68, -7, 55, 58, 124, -6, -20, 41, 38, 49, -74, -90, -1, -127, 5, 89, -60, 38, 44, -17, -117, -38, 15, -112, -11, 106, 39, 14, -108, -86, -106, 75, -23, 13, 109, 76, 66, 120, -89, -40, 105, 9, 88, -18, 13, 119, -83, -70, -39, 38, -97, 41, 36, 48, -24, 104, -124, -34, -69, -53, -4, -24, 37, 45, -51, 7, 38, 48, -25, -87, 71, 73, 62, 105, -37, 27, -6, 20, 15, -7, -22, 109, -35, -11, 51, 22, -83, -92, 61, -75, 103, 53, 96, -61, 50, -84, -85, -101, -74, -92, 22, 2, -85, -23, 93, 90, -102, 8, 32, 115, -105, 124, 7, 3, -105, 123, -84, 30, 96, 50, 28, -27, -94, 75, 118, -31, -68, 53, 55, -109, -17, -124, 46, 117, 95, -95, 41, 20, 10, -58, 39, 110, -22, 21, -96, 79, 89, -19, 84, 118, -28, 63, -12, 16, 14, -84, -7, -107, 101, 117, -35, 32, -52, -38, -102, 113, 98, -22, 120, 19, -7, -116, 5, 86, -116, 116, -90, -128, -86, 9, 83, -72, -120, -119, 19, -72, 24, 58, 14, -109, -15, -122, 13, -46, 22, -60, 67, 81, -115, 106, -53, 92, -9, 120, 60, -73, -3, -63, -70, 122, 33, 61, -115, -127, 34, 60, -5, -105, -5, 67, 37, 0, -19, -5, -78, -105, 81, 17, -32, -33, -48, 60, -16, -15, -81, 90, 0, -74, 127, 68, -103, -95, -4, 23, 86, 93, -103, 33, -39, -82, -41, -98, 45, 88, -40, -12, 5, -123, -34, 23, 5, 20, 8, -53, 0, 10, -38, 65, 64, -118, -8, -37, -107, 9, 34, -127, 77, 51, -72, 17, 1, -7, 76, -63, -62, 65, 69, -49, 116, -112, 92, -16, 64, -123, -96, -103, 55, -41, 25, 56, -3, -42, 126, -104, -13, -7, 88, 112, -126, 102, -62, 96, 47, 125, 50, -124, -28, -56, -124, -77, 0, 55, -116, -86, 110, 100, -72, -114, 87, -59, 109, 31, -94, -40, -94, 54, -82, -110, 110, -61, 54, 28, -75, 77, 57, 16, -100, 24, -85, 33, -8, -98, -85, -66, -29, -128, -45, -77, 119, 15, 107, 20, -2, -28, -81, -108, 122, -13, -16, -12, -42, -37, 26, -53, 91, -120, 29, -22, 15, -70, -39, -88, -77, -50, 52, 50, 92, 92, -65, 67, 99, 119, 32, -118, -44, 5, 24, 108, -89, 95, 108, 87, 76, 112, 87, 50, -102, -108, -126, 51, -27, 114, 82, 17, 63, 44, 61, 13, -123, 15, 60, 3, -54, 49, 35, -60, -32, 13, 43, 11, -3, 12, 13, -5, 96, 102, 88, -81, -51, 117, 20, 7, -69, 102, 15, -119, 116, 109, -57, 17, 52, 12, -73, 100, -65, 100, -18, 40, 98, -48, -80, 89, 47, 93, -26, -52, -121, 44, 105, -94, -76, 49, -36, 113, -26, 78, -13, -64, -40, -40, -20, 84, -122, -56, 9, -116, 73, 29, -34, 27, 116, 47, 108, -51, -108, -33, -24, -68, -16, -29, -12, 45, 31, -68, 35, -31, 118, 41, 45, -101, -42, -91, -74, 38, -116, 6, -47, -51, -95, -85, 100, 7, -10, 79, 108, -48, 88, -114, 57, 59, 89, -43, 80, -98, 6, 78, 88, -122, -35, 14, 89, -75, 116, 104, 88, 124, -105, -82, 80, -45, -1, -44, -39, -43, -74, 86, -108, 115, -64, -85, -5, -100, 22, -121, 92, 62, -101, -98, 6, 34, -66, 90, 51, 88, -88, -85, 6, -67, -112, -19, 19, -24, -70, -24, 65, 81, 43, 31, -40, -27, -79, -68, -103, -17, -39, -92, 122, -115, 81, 98, 103, -15, -72, -112, 0, -24, 44, 74, 37, -53, 19, 121, -49, -79, 72, -122, 46, -57, -43, 98, -117, -73, 117, -95, -104, 48, -76, -100, 111, 18, 29, -82, -97, 17, 99, 53, 27, -13, 125, -76, -50, 110, -48, -51, 41, -115, -97, -38, -35, -124, -128, -12, 60, -95, 92, -35, -50, 14, 65, 72, -7, 110, 6, 104, 115, -39, -19, 16, 114, -73, 106, -77, -34, 27, 108, -101, -22, -11, 97, -26, -35, -9, -62, 26, 122, -28, 111, -114, -46, 111, 84, 121, -125, -68, -41, 0, -51, 117, -82, 39, 119, 118, 59, -50, -31, 72, -127, -22, -122, -115, -106, 11, 115, 44, 92, -83, 60, 63, -60, 91, -41, -91, -20, 56, 56, -71, -16, -54, -54, 101, -34, -70, 75, -29, 89, -11, -46, 77, 120, -110, -122, -88, 125, -25, -123, 69, 33, 124, -55, -5, 29, -123, -122, -84, -20, -87, -82, -128, 111, -94, -61, -88, -41, 123, -113, -47, 5, 67, -95, 24, -47, 30, 88, 96, 121, -109, 0, -39, -118, 106, -120, 118, -128, -77, 18, 62, -87, 103, 16, -87, -70, -103, 73, 41, -116, 30, -61, -23, 123, 44, 58, 40, 27, 50, -31, 104, -50, -116, -126, -74, -107, 55, 52, 90, 37, 69, 16, -61, -121, 93, 86, 53, 103, 54, 32, -124, -21, -19, 49, -113, -61, 71, -89, 2, -55, 114, -57, 10, -104, 69, 6, 2, -41, -106, -89, -50, 35, -45, 55, 14, 7, -117, 105, 71, 3, -50, -57, 28, -120, 90, -55, 35, 82, 20, 89, -48, 84, -16, 85, 30, -18, 127, 54, -18, 83, -63, -95, 97, -60, 27, 2, -59, -52, 7, -83, -2, -33, -103, -42, 29, -34, -10, 97, -81, 124, -39, 13, 39, -27, -82, 26, -66, 65, -1, -96, 86, -105, -45, -64, 55, 33, 64, -15, -123, 6, 105, -10, -7, 59, -55, 82, -99, -63, 19, -11, 28, 51, -72, -38, -84, 119, 0, 90, 93, 60, 39, 70, 11, -58, -10, -79, 14, -38, -14, -126, 113, 33, 35, 81, -48, 117, -56, -81, -32, -11, -66, 84, 99, 85, 14, 86, -107, -34, 57, -100, -89, -92, 5, -36, -26, 96, -14, -124, 11, -95, -37, -62, -23, -68, 73, 41, 20, 126, 101, -21, -44, 63, 12, 61, -48, -10, 20, -34, -24, -102, -89, 41, -68, -57, -59, -2, -29, 97, 84, -89, -9, -58, -121, 85, 85, 82, 2, -5, 29, 34, 90, -74, -2, 112, 42, 74, 69, 39, 24, -15, -124, 18, -97, 48, 68, 75, -76, -74, -94, 0, 1, 66, 34, -44, -89, 75, -114, 18, -105, -14, 92, -28, -99, -24, -20, -65, 56, 3, 104, 52, -58, -4, 17, -112, 127, 61, -16, -41, 104, 18, -127, 6, 67, 71, 63, 4, -119, -19, 69, -93, 1, 8, -16, -32, 77, 110, 63, 8, -12, -89, -35, 28, 12, 79, 45, 81, -69, -106, -120, 38, -118, -25, 82, 100, -103, -128, 54, 76, -115, -9, 42, -50, -70, 114, -105, -4, 28, 116, 50, 123, 126, 55, 105, -79, -105, -64, -9, 76, 5, -35, 46, -2, 119, -50, -13, -53, 101, -17, 102, 55, -120, 87, -1, -116, -70, 26, 11, -74, 17, -86, -57, -54, 9, -8, -95, 57, 31, -77, -23, 73, -28, 31, 75, 10, 50, -54, -64, -81, 104, -2, 56, 14, 95, 37, -1, 125, -27, -13, 3, -11, 50, -71, 125, 8, -93, 66, 102, -83, -11, 103, -33, 67, -12, 34, -113, -101, -108, 98, 123, -80, 9, 116, 29, 4, -33, 19, -40, 90, -53, -125, 123, 2, 111, 69, 70, 83, -13, 49, 64, 68, -114, -80, -51, -98, 73, 52, -4, 103, 56, -16, -124, -64, -39, 35, -5, -62, 126, -12, 53, -128, 118, 57, -41, -18, 4, 49, 120, 92, -6, -71, -102, 10, 88, 34, 99, 101, -110, -40, -18, -26, -124, 58, -108, -85, -106, 78, -42, 61, -63, 102, -128, -93, -97, 77, -123, 105, -95, 103, 115, 74, 87, 67, -19, -102, -123, 64, 21, -31, 126, -18, -42, -80, 60, 109, 59, -50, -90, -104, 69, 45, -123, -122, -24, -104, 34, -89, 46, -90, -86, 2, 67, 4, -77, 111, 10, -115, -70, 116, 101, 114, 19, 114, 104, -26, -14, 40, -26, 25, 27, 3, -29, -21, 110, -122, -53, 21, -85, 32, 82, -68, -112, 87, 110, 33, -52, -6, -2, 107, 54, -74, -93, 110, -39, -17, -21, 55, 116, -1, 28, 50, 113, -49 );
    signal scenario_output : scenario_type :=( -22, 12, 30, 22, -2, -34, 70, 6, -120, 28, -27, -4, 8, -7, 80, -25, -42, 26, -63, 58, -62, 55, 39, -43, -6, -70, 36, -18, 63, -2, -38, 52, -17, 35, -25, -49, 66, 11, -27, -32, -18, -11, -61, 47, -20, 8, 1, 30, 3, 17, 39, 14, 17, -25, 85, 20, -23, -38, 42, 15, -14, 20, -53, -11, -80, -40, -14, -57, 18, -1, 71, 18, -13, -34, 41, -27, 11, 18, -20, 51, -15, 36, -9, -40, 3, -17, -2, -9, -52, 5, -54, 30, -60, 117, -13, 58, -10, -7, -46, -45, 3, 3, -8, -45, 45, -42, 0, -17, -63, 1, -30, 49, 12, 60, -7, 66, -97, 35, -2, -79, 58, 32, -8, -6, -10, -14, 0, 56, -21, 15, 1, 21, 22, -15, 38, -102, 12, -10, -24, -39, -24, 40, -6, -31, 40, 27, 64, -22, -48, 29, 11, -64, 89, -18, -17, 56, -46, 55, 19, -35, 53, -97, 51, -6, 27, -54, -9, -3, 14, -73, 77, -54, 14, -21, 11, 15, -22, 28, 18, 66, 40, -1, -25, 17, 12, -48, 47, 60, -14, 9, -11, 11, 28, -46, -32, 11, -41, -13, 3, -11, 13, -93, 1, -26, -7, -45, 48, 48, 12, 38, 47, -48, 36, -51, -57, 27, -17, 25, 31, 11, -10, 32, -4, -4, 51, -29, -20, -49, 53, -20, 8, -9, -42, 63, 15, 2, -7, 28, -38, -2, 52, -38, -18, 63, -2, 75, 2, -24, 12, 3, -46, -11, 5, 59, -56, -7, 47, -32, 55, -22, -15, 2, -3, 46, -30, 2, 35, -63, 61, -48, 88, -40, 15, 2, -14, 64, -13, 36, 12, -15, -63, 23, -5, -24, -10, -7, 42, -51, 69, 28, -64, 6, -43, -45, -5, 8, 1, 13, 27, -78, -29, 34, -22, 53, 66, 37, 11, -20, 64, 11, -41, 0, -53, 9, 54, -23, 41, 65, -89, 22, -48, 1, -9, 17, 44, -64, 28, 13, -46, -18, -53, 31, 13, 37, 44, -29, 13, -1, -6, 7, -66, 79, -92, 2, 59, -14, 80, -3, -2, 26, -12, 23, -91, 40, 14, 53, 32, -4, -1, -14, -13, -2, 4, 6, -34, -22, -8, 29, -9, -45, 18, 10, 43, -58, 8, -5, 28, -15, -46, 53, -38, 54, -14, 9, 8, 49, -7, 6, -51, 76, -68, 90, -51, -61, 56, -17, 51, 3, -24, 18, -31, 0, 36, -74, -2, 23, -74, 94, 5, 2, 9, 24, -24, 17, -49, -35, 32, 19, -27, 94, -44, 41, -27, -46, -47, -75, -34, 22, -18, 36, 42, 21, 11, 20, 30, -4, -58, 7, 17, 25, 6, -9, 12, 24, -52, 43, -18, -74, -2, 10, -15, -56, 44, -26, 100, -5, 23, 6, -8, -58, 11, -9, 9, -45, 5, -11, -63, 103, -6, 46, 21, 3, 64, -39, -5, 19, 28, -68, -22, 5, 7, 87, -8, -6, -17, 21, -7, -74, -4, 18, 44, -8, 39, 46, 30, -88, -3, -45, -40, 17, -22, 75, -11, 55, -44, 15, 4, -74, 7, -14, 62, -13, 43, 37, 45, -14, -24, 36, -32, -31, 65, -58, -11, -13, 25, 10, -34, -11, 35, -15, -4, 31, 1, 39, -32, -27, 57, 27, 10, 68, -18, 22, -26, -91, 60, 24, 4, 23, -23, 70, -14, -5, -18, -63, 18, -22, 12, -55, -9, 25, -13, -19, 0, 35, 39, -29, 74, -26, -35, 66, -39, 88, -51, -11, -15, 47, 29, 5, -25, -19, -42, -40, -18, 18, -23, 19, 44, -56, 95, -45, 25, 0, -44, 24, -23, 13, 13, 6, 79, 17, -44, -2, 0, -19, -4, 36, 0, 32, -28, 63, -28, -65, 0, 3, -14, -8, 0, 60, -56, 42, 28, 34, 24, -11, 60, -94, 83, -3, -17, 8, -20, -12, 8, -15, 59, 22, 27, -38, -37, 2, 24, 10, -18, 7, 15, 15, -44, -46, -17, -23, 4, -39, 49, -57, -4, -7, -31, -68, 26, -15, 17, 4, 10, 22, -36, 36, -6, 61, 7, -17, 29, 42, -61, 61, -79, -30, 48, -31, 89, -38, -30, -3, 21, 29, -9, 8, 5, 62, -28, 29, -49, -31, 17, 37, 2, -35, 78, -106, 15, -49, -38, 62, -66, 90, -86, 9, -2, -83, 59, 2, -9, 58, -75, 5, -74, -38, -7, -3, 39, 58, 2, 72, -55, 11, -25, -100, -2, 29, -51, 77, 9, 6, 30, -57, -22, -26, 39, -55, 15, -80, 46, 38, -28, 25, -29, 10, 45, -64, 39, 17, 30, -6, -19, 12, -51, -31, 34, -9, 32, 11, -18, 55, -71, 49, -24, -51, 54, -56, -49, 51, 0, 40, 13, 5, 19, 44, -96, 70, -37, -21, -25, 22, 11, 30, -43, -39, 10, -4, -22, 38, 18, -19, 6, 58, -62, -10, 20, 0, 38, -35, 18, -68, 17, -6, 0, 32, 36, 57, -20, 59, -103, 29, -2, -58, 15, -13, 41, -23, 39, 9, -11, 68, -2, -54, 60, -20, -6, -14, -90, 45, -2, 11, 40, 40, 15, -75, 45, 6, -40, 41, 1, 26, 17, 8, -6, -18, -14, 7, -61, 68, -56, -8, 97, 23, 29, -1, -13, -28, -41, 12, -45, -4, 25, 55, -37, -10, 46, 43, -7, 0, 47, -54, -46, 28, 45, -14, -3, 0, -6, -40, -29, -31, 0, 63, -38, -7, 71, -25, 1, 25, -65, 39, 10, -74, 48, -53, -19, -44, 17, 69, -35, 29, -46, 45, 9, -68, 65, -52, 12, -7, 15, 52, -39, 37, -29, -27, -4, -8, -56, 17, -14, 38, -9, 13, -17, 47, -29, -103, 3, -14, 41, 4, -66, 8, -43, -23, 15, -40, 52, 56, -42, -6, -61, -23, -9, 25, -35, -12, 21, -8, 3, -47, 31, 17, -86, 99, -18, 51, -22, -30, 2, -38, -25, -76, 66, 25, -32, -4, 39, 9, -19, -113, -1, 11, -26, -11, 17, 3, 96, 4, 46, 21, 31, 32, -56, 52, -81, 13, -26, -70, 34, -71, 71, -43, 102, -5, -29, 4, -37, 3, -61, -21, 24, -49, 108, -46, 11, 12, 5, 26, -15, -12, 25, 19, -57, 99, -65, -60, 25, -3, 54, -4, 9, 26, -1, -12, -30, -66, 32, -10, -66, 61, -73, 68, -48, -41, 79, -13, -21, 69, -25, 34, 26, -82, 68, 14, -80, 59, -110, 21, 13, -68, 53, -70, -24, 42, -54, 71, -11, 5, 27, -4, 3, -37, 87, -65, 69, -24, 12, 70, -43, 5, 41, -47, -21, 28, -57, -21, 29, -85, 69, -56, -30, 71, -32, 19, 110, -8, -44, 66, -52, 43, -8, -74, 41, -20, -42, 22, 0, -34, -44, -20, 7, 34, 0, 2, 22, -59, -11, -5, 8, -86, 69, -91, 37, 32, 1, 55, -42, 58, 12, -82, 3, -44, 12, 64, -42, -36, 34, -28, 64, -20, -29, 54, -66, 58, 10, -52, 37, -64, 23, -32, 8, -19, 79, 6, -29, 9, -36, -39, -48, -66, 48, -31, 38, -27, -14, 28, -80, 25, 8, -24, 46, 35, -15, 36, 37, -17, -27, -14, -28, 19, -23, 23, 26, -93, 10, 38, -19, 85, -1, 0, 13, -47, -64, -57, -34, -11, 59, -14, 27, -72, 32, -12, 22, 27, -5, -13, 2, -7, 28, 14, -52, -24, -1, -27, 0, -10, 68, 27, -8, 8, -3, 23, -68, 77, 22, 56, -38, 1, 38, -52, 27, -110, 57, 1, -51, 77, -4, 75, -40, -23, -3, -32, 22, -7, 21, 69, -23, 8, 54, -17, 15, -72, -6, -12, 20, -27, 35, 15, 19, -27, -25, 44, -30, -18, 46, -26, -21, -1, 4, 31, -40, 41, -14, 127, -38, 6, -12, 28, 9, -30, -6, -17, -48, 3, 4, 3, -24, 0, 20, -49, 29, -90, 82, 22, 2, -23, 17, -22, 9, -13, -99, 9, -34, 41, 24, 20, -3, -5, -1, -52, -20, -48, -18, 55, -40, 61, 21, -59, 15, -13, 1, -14, 0, 81, 40, 14, 15, -75, 4, -34, 6, -29, -8, 106, -37, -29, 10, -39, 81, 2, 37, 37, 10, 83, -56, -51, -27, -34, 20, -36, 1, 21, -19, 72, -54, 0, -69, 8, 13, -30, 31, 71, -19, -64, 45, 8, -23, 68, -31, 3, 15, -87, 6, 17, -46, 27, -1, -57, 0, 19, 13, 3, 78, 17, -41, 28, -54, 12, -4, -27, 36, -1, -5, 85, -23, 68, -25, 25, -5, -34, -21, -44, -24, -2, -36, 96, -24, 10, 12, -27, 30, -66, 56, -90, 14, 5, 4, -10, 19, -14, 54, -15, -28, 35, 39, 6, 11, -56, 37, -61, 36, -64, 11, 62, -19, 9, 70, -35, 81, -36, 0, -45, 2, -39, 23, -27, 14, 89, -27, -31, 49, -3, -95, 74, -21, 21, 30, -2, 43, -54, 19, 5, -99, 109, -43, 57, -35, -26, 61, 13, -10, -11, 37, -26, -32, 1, -40, 8, 29, 25, -14, -10, -11, -14, 22, -73, 28, -17, 0, 23, 54, -11, -63, 57, -42, -34, 17, -30, 70, -8, 21, 85, 27, -36, -6, -27, 2, 6, -55, 34, -19, 77, -55, 0, -7, -20, 0, -35, 3, 38, -61, 10, 63, -36, -3, -40, 86, -61, 7, 1, 39, 44, 10, 25, 31, 58, -34, 18, -29, 29, -77, -11, 1, -28, 74, -1, -1, 15, -9, -79, 90, 11, 4, -14, 21, 11, -80, 4, 26, -29, 47, -54, 17, 6, -20, 25, 36, -72, 42, -13, -28, -51, -81, -24, 44, -46, 77, 32, 29, 37, -43, 63, -26, -25, 0, 48, -14, 36, -34, 45, 3, -83, 31, -54, 15, -18, 11, 8, 5, 38, -41, -18, 37, -26, 2, -74, 18, 29, -20, 8, 55, -23, 3, 4, -17, 45, -53, -11, 0, -29, 61, -58, -6, 85, -34, 38, 4, 11, 9, 23, -32, 24, 37, -45, -28, 81, -30, -11, 73, -42, 44, -30, 5, -12, 7, 0, -80, -28, 26, 8, -37, 7, 3, 22, 4, 22, 10, 2, 123, -20, 35, 3, -15, -60, -74, -57, -4, 1, 8, 28, 14, -20, -2, 34, -57, -29, 49, -13, 9, -20, -1, 52, 22, 47, 87, -65, 0, -26, 5, 20, -60, -17, 21, 18, -38, 14, 29, -12, 7, -61, -4, -31, 0, 9, -43, 83, -109, 26, -42, -18, 2, -90, 11, 9, 38, 36, 57, 14, -2, -52, -9, 9, -20, 58, -20, 5, 6, -13, 6, -42, 57, -24, -8, 86, 6, 62, -46, -7, 0, -3, -19, 0, 34, 23, -35, -20, 51, -38, 49, -74, 47, -34, -7, 26, -70, 65, -4, 8, 6, -61, 39, 15, 23, 3, 45, -61, 2, -1, -3, -49, 7, 93, -48, -9, 8, -31, 1, -37, -5, 99, -11, -29, 17, 7, -2, -64, -18, 83, -23, 21, -9, -29, 47, -47, 76, -5, 15, 38, -8, -37, 72, 3, -54, -17, -35, 14, -34, 0, 64, -19, 77, -37, 29, -76, -2, -40, 41, -76, 34, -6, -45, 94, -38, 47, -92, 34, -12, -15, 3, -17, 14, -21, 28, 14, 51, -25, 49, -57, 62, -18, 8, 20, -17, -42, -27, 22, 6, 8, 3, -40, -11, 0, -48, -6, 30, -39, 78, -62, 35, -3, -2, 34, -5, 38, -87, 21, -6, -48, -22, 14, 14, 12, -75, 7, -11, -5, 5, 28, 20, -11, 26, -23, -25, 76, -4, 27, 22, 83, -69, -6, 6, -32, -19, -30, -11, -30, 2, 22, 0, 48, -7, 26, -52, 116, -19, -10, 28, -41, 22, -17, 17, 13, 3, -6, 9, -8, -58, 20, -37, -46, 63, 6, -23, 9, 0, 39, -75, 57, -22, 90, -2, -42, 65, -85, -2, -32, -53, 51, -73, 22, 71, 1, -19, 4, 4, -63, 43, -39, 40, 11, 10, 10, 18, -23, 18, -54, 46, 31, 27, 10, 17, -7, 13, -10, -53, 20, -17, 10, 10, -11, -11, 27, -55, 11, 28, 12, 64, -8, 25, 23, 40, -5, -36, 56, -25, 23, -34, 7, -43, 7, -37, 85, -21, 58, -25, 39, -9, -73, 7, -51, 22, -21, -24, 49, -61, 42, -21, -62, 109, -44, 93, 8, -25, 74, -61, 5, 65, -78, 7, 4, -63, 76, -41, 12, -19, -10, 42, -32, 9, 58, 52, -13, 76, -66, 15, -36, -36, 18, -4, -85, 37, 15, 21, 27, -47, 25, -35, -9, -12, -24, 76, -24, 1, 24, -40, 45, -56, 59, -59, 90, -40, 17, 54, -88, 45, -43, 32, 40, -30, 38, 1, -6, 37, -57, 93, -36, 6, -27, -20, -29, -12, 25, -113, 75, -58, -5, -32, -24, 107, -46, 18, -32, 21, 17, -68, 60, -39, 4, 22, -23, 72, -53, -8, -4, -73, 30, 30, -11, 49, 17, -41, -44, -49, 39, -8, 23, 43, 21, 21, 40, -49, 48, -29, -52, 23, 42, -28, 10, 15, 8, 1, 54, 0, -36, 72, -65, -30, -24, -43, 53, -8, 48, -8, 85, -80, 39, -11, -63, -38, -74, -11, 31, -18, 43, -52, -22, 21, 30, -17, 34, 17, 3, -34, -35, 5, -64, 54, 9, 5, -9, 24, -19, 24, -3, -44, -11, 46, -42, 9, 19, -68, 36, 1, 27, 40, 23, 5, 78, 2, -57, 19, -37, -51, 12, -39, -41, 76, 28, -6, -24, 40, -25, -64, 24, -94, 98, -51, 29, 59, 12, 15, -64, 0, 24, -5, 27, 31, 36, 17, 8, -17, -14, 20, 55, -11, -3, 11, -25, -30, -27, 24, -39, 14, 17, -40, -39, 12, -35, -5, -62, 34, -6, 29, 45, 12, 68, -21, -72, 3, 9, -3, -13, -7, -6, 30, -62, 41, -8, 38, -21, -6, -4, 31, -37, -39, 15, 15, -88, 6, 45, -15, 34, 14, 75, -11, -19, -26, -12, -5, 18, -20, 62, -73, -10, 47, 1, 10, -28, -6, -20, 47, -88, 62, -46, -15, 90, -19, 6, 31, -24, 0, 15, -23, 61, -43, 29, 5, 31, 9, -8, -17, 40, -8, 48, -55, 21, -87, 19, 13, -45, -15, -41, 91, -31, 17, 46, 32, 68, -8, -10, 19, -52, 5, -30, 31, 54, -63, -2, 3, -15, -49, 36, -94, 12, 8, -31, 31, -41, -38, 6, -2, -34, 125, -14, -13, 43, -34, -38, -29, -49, 54, 34, -28, 9, -42, -39, 10, -38, 43, 36, 34, -2, 45, -18, 79, 44, -5, -54, 9, -34, 22, -36, 13, 34, -71, 63, -113, 92, -15, -27, 62, -15, 65, 23, -42, -2, 3, -79, 20, -2, -30, 89, -36, 35, -4, 32, -25, -20, 10, -68, 28, -56, 86, -38, 69, -22, 46, -64, -27, 19, -23, 20, -19, -14, 31, 8, -23, 29, -58, 13, -53, 23, 13, -24, 74, -11, 80, -58, -9, 64, -10, 6, -51, 30, 2, 5, -5, -1, 20, -26, -40, 5, -4, 58, -14, -14, 59, -8, -19, -36, -8, -44, -37, -42, -51, 18, -31, 25, 23, -39, 23, 52, 24, -40, 18, 39, -32, 28, -34, -17, -25, -74, 1, -34, 4, 19, -29, 39, 0, -25, 40, 13, -53, 19, 11, 77, -74, -34, -35, -36, -23, -5, 15, 29, 30, -45, 28, 69, -31, 21, -2, 18, 7, -10, 90, -80, -8, -3, 4, -25, -2, -71, 43, -39, 32, -22, 38, 69, -20, 71, -27, 44, -36, -44, 5, 7, -51, -19, -88, 0, 25, -13, 44, 9, -15, 15, -82, 27, 17, -7, 14, 2, 57, -5, 26, 37, 45, 13, 8, -9, -28, 19, -94, 82, -66, 65, -4, 18, 11, -15, 56, -13, 34, -21, 24, -41, -26, 0, -10, -86, -21, 23, 68, -44, -57, 3, -39, 36, -22, -3, -30, 81, 2, -1, 27, -23, 21, 62, -39, -56, 68, -10, -7, 19, -89, 11, -38, 23, 0, 11, 31, -10, 54, 2, 15, -14, 42, -6, 11, -42, 26, -8, -56, -32, -20, -28, -71, 1, -28, 39, 4, -27, 62, 27, 55, 14, -47, 8, -60, -53, -31, -34, 44, 14, 21, -37, 52, 28, -71, 37, -37, 66, -34, 14, 48, 18, -35, -35, -38, -38, -25, 48, -26, 19, -14, -28, -22, 40, -13, 43, -3, -17, -18, 29, 1, -79, 52, -81, 26, 1, -7, 19, -63, -18, 27, -14, -13, -13, 72, 28, 40, -9, -4, -8, -22, 10, 4, -41, 8, -27, 26, -104, 69, -8, -41, 92, -35, 49, -106, 18, 10, 7, -4, -25, 21, 37, 10, -43, -23, -38, -5, -18, -34, -6, 22, 75, -24, -7, 42, 3, -11, -61, 4, -65, 15, 0, -74, 22, -51, -26, -18, 26, 15, 49, 10, 44, -44, 53, -12, -55, 51, 20, -52, 20, 39, 17, -46, 9, 63, -8, -8, 0, -32, -8, 5, -74, 38, -34, -41, 17, 45, -44, -11, 61, -42, -8, 43, -18, 37, 41, -10, 48, -111, 19, -5, 1, -61, -29, -17, 52, -47, 48, 31, 31, 4, 7, 85, -81, 48, -47, -3, -11, -14, -34, 63, -66, -29, 61, -11, 12, -53, -1, 13, 47, -31, 13, 2, -66, -36, 10, 2, -6, 44, 52, -2, -22, 23, -20, -44, -42, -29, -38, 42, -48, 36, 70, 10, -9, 11, -30, -37, -31, -60, 36, -23, 24, -10, -89, 49, -7, -22, -36, 10, 80, -58, 21, -9, -60, 31, 18, -34, 28, 4, -15, 22, 41, 2, -35, 76, -92, 41, -61, -42, 106, -49, 27, -4, -63, 77, -12, -3, 1, -21, 111, 42, 21, -39, 23, -26, -30, -32, -49, 127, 13, 5, -34, 18, -45, 24, -25, -22, 18, -15, 3, -6, 22, -20, 114, -105, 25, -24, -43, 38, -78, 60, 38, -11, 30, -42, 23, 2, -71, 31, -23, -17, 26, 32, -63, -49, -17, -29, 45, -35, 30, 51, -41, -21, -51, -42, 25, 9, -8, -4, -14, 40, 26, 28, -38, -11, 13, -31, 34, -7, -44, 56, -8, -24, -57, 4, -35, 18, -24, -83, 11, -42, 14, -62, 3, 42, -7, 45, 35, -1, -43, 32, -18, 27, 40, 1, 11, 22, -5, -74, -25, -45, 25, 9, -48, -47, 3, -9, 6, 85, -2, -19, 39, -46, 51, -49, -31, -9, -69, 56, -31, 23, 42, 31, 4, -55, 13, -58, 46, -46, 34, 13, 65, 55, 51, 34, -59, -25, 0, 40, -10, 46, -14, 63, 44, -89, -30, -81, -23, 32, 8, 29, -15, 11, -22, 62, 4, -11, 68, -17, 3, -23, -89, -14, -13, 0, -42, 20, 17, 44, -2, 19, -4, 13, -2, -41, 35, -57, 95, -51, 51, -44, 23, 9, -42, 12, -74, -44, -4, 30, -17, -3, -24, -27, 9, -14, 63, -69, 12, -27, -3, 13, -7, 42, -55, 0, -6, -64, 37, 11, -85, 39, 5, 5, 56, -23, 0, 15, -43, 8, -44, -45, -24, -49, 4, -83, 127, 0, 30, -22, -20, -2, 1, -8, -47, 19, -3, -19, 53, -51, -38, 100, -26, 14, 17, -2, 69, -75, 14, 60, -75, 27, -15, -52, 69, 31, 14, 28, -22, -56, -6, 38, -8, 1, -29, 19, -4, -44, 65, -31, 38, -51, -12, 31, 30, 3, 15, 12, 4, -83, -38, -36, 43, -3, 13, 72, -12, 48, 56, -110, 35, -54, 49, 11, -48, 20, 1, 23, -40, -73, 10, -5, 0, 12, -31, 40, 24, -1, 28, 0, -13, 76, -11, -59, 42, -54, 51, 13, 12, -3, 9, -44, -52, -2, -46, -34, 79, 3, 52, -42, -10, -28, -17, 1, -10, 46, -18, 39, 19, -106, 32, -8, -58, 89, -49, 34, 14, -18, 43, -58, 2, 11, -68, 28, 56, -11, 11, -68, 35, 30, -10, 36, 5, 53, -52, 64, -61, -21, -14, -21, 44, -14, 31, 6, -32, 6, -10, -38, 27, -51, 41, -105, -20, 45, 26, 12, 9, -27, 65, 53, -66, -13, 43, -31, 31, -105, 24, 32, -20, 35, -42, -26, -48, -34, 35, 36, 74, 14, -7, 14, 20, 15, -98, 56, -38, -4, -38, -89, 8, 37, -13, 24, 63, -1, -1, -26, -31, -2, -5, 5, 18, -29, -40, 27, 6, -29, 26, 61, 47, -13, 2, 25, -39, -92, 7, -39, 28, 32, 24, 22, 15, 7, 43, -104, 68, -10, 46, -78, -37, -7, 24, 19, 15, 58, -30, 20, -12, -7, -49, -71, -8, -51, 18, -37, 18, 69, 0, 6, 90, -82, 17, -9, -24, -72, 62, -30, -2, 70, -42, 55, -44, 73, -57, 7, -51, 52, -5, 14, -48, -5, -5, 24, -43, 13, -75, 46, 22, 25, 31, 13, 0, -24, -11, 44, -7, 8, -49, 29, -21, -35, 34, -49, 10, -14, 28, -6, 65, -83, 41, -36, -85, 26, -28, 47, 24, -47, 23, -97, -10, 4, 7, 12, 8, 62, -42, 109, -34, -14, 20, -97, -2, 53, -30, 62, -26, 30, 59, 10, 28, -31, 27, -46, -35, 17, -18, -71, -18, -34, 21, 28, -11, 0, 15, -1, -46, 45, 8, -9, 79, -61, -12, -13, -34, 26, -85, -15, 44, -13, 47, -7, 62, -46, 54, -63, -7, 40, -47, -14, 26, 59, 14, 21, 65, -52, 39, -5, -5, -44, -3, -35, -31, -27, -22, 78, -44, -30, 74, -45, -32, 23, -30, 80, -7, -64, 39, -37, -77, 59, -13, 58, -23, -17, 39, 28, -64, 18, 91, 2, -23, 0, 34, -19, 1, -46, 14, -34, 80, -35, 45, -37, -21, 40, -20, -18, 15, -25, 44, -40, 47, 7, 8, 51, -10, 38, 6, 61, -29, 15, 61, -18, -47, -22, -25, 6, -53, 2, -12, 26, -2, -4, 89, -23, -44, 28, -2, -29, -44, 38, 43, 35, 42, -26, 43, -90, -1, -6, 2, -46, -28, 54, 56, -37, -18, -21, 5, -15, 4, 12, 41, 18, 83, -7, -58, 19, -6, -6, 39, -11, 6, 23, 10, 1, 4, 40, -5, 25, 53, -75, 4, -28, -97, -2, -25, 0, 20, 31, 70, 69, 49, 38, -37, 41, -47, 6, -55, 64, -11, -72, -3, 1, 13, -52, 62, -24, 32, 52, -83, -39, 8, 5, 14, 43, -31, -9, 34, 45, -4, -5, -3, -2, -53, 10, 0, -57, 23, 35, 2, -18, -3, -36, -35, -1, -9, -37, -22, 105, -71, 70, 37, -46, 46, -128, 31, 1, -46, 20, -23, 32, 35, 65, 35, 28, -19, 57, 42, -45, 5, -1, -29, -25, 4, 47, -10, -57, -2, -30, -28, 66, 19, 12, -27, -9, 3, -6, -55, -27, 2, 56, -11, -3, 10, -6, 35, -9, -36, 74, -34, -10, 14, -24, -38, -13, -52, -58, -39, 66, -25, 25, 11, 43, 41, -31, -3, 43, -26, -23, -21, -9, 5, -55, 15, -58, 43, -12, 48, 12, 80, -17, -1, -10, -48, -7, 21, -20, -22, 45, -80, 31, -51, 40, -30, -39, 63, -79, 117, -42, 29, -9, -12, 64, 10, -58, 27, -31, 2, -35, -4, 32, -108, 45, -37, 0, -65, -30, 30, -4, -5, 18, 28, 8, 20, 44, 17, 32, 58, -3, 6, -9, 20, -19, -71, 44, -42, -62, 42, -48, 56, 41, 37, 0, 18, -63, 18, 49, -49, 4, 23, -102, 38, -19, 31, -18, 11, 54, 19, -10, -35, -8, 35, -55, 6, 35, -38, 51, -46, 89, -66, 13, 77, -21, -65, -10, 21, 18, 22, 56, 37, -26, 36, -85, 41, -1, 45, -17, -36, 49, 6, -53, 30, -61, 20, 36, -68, 22, -14, 29, -44, 6, 19, 13, 14, -45, 8, -27, 8, -26, -5, -10, 116, -12, 10, 63, -51, -19, -23, -54, 44, 0, -30, 39, 18, -59, -24, 10, -14, -7, -22, 11, -37, 6, 5, 37, 25, 62, -1, -42, 65, -60, 95, -70, -58, 49, 3, 34, 10, -32, 35, -38, -1, 29, -20, 15, 51, -14, -9, -63, -1, -45, 68, 0, 22, 1, -7, -12, -19, -6, 45, -4, 4, 14, -56, 34, 18, 54, -3, 7, 30, 0, 13, -51, -11, -4, -41, -79, 54, -9, -15, 7, 0, 56, -21, -2, 52, -2, -12, 53, -5, -69, 68, -59, 8, 14, -13, 63, -105, 51, -24, -35, 43, -69, 60, -24, 43, -56, 18, 20, -108, 36, -4, -61, 98, -83, 6, 76, -30, 38, -22, -13, -12, 24, -44, 85, -40, 41, -74, 12, -8, -69, -9, 83, -18, 45, -59, 28, -1, -71, 41, -6, 46, 13, 39, -19, 14, -36, -24, -37, 22, -39, 3, 15, -29, 62, 30, -9, 6, 44, -72, -5, 2, -58, 24, -6, -30, 20, -2, -46, 66, -76, 26, 55, -65, 47, -91, 28, 38, -29, -35, 38, 14, -2, -41, -23, 42, 0, -13, -4, 3, 59, -44, 48, -39, 55, 15, 1, 59, -94, 32, -48, 0, -56, 40, 55, -39, -3, 23, -41, 10, -31, -95, 58, 0, 40, 66, 20, -28, 21, -24, -5, 5, -23, 13, 18, 37, -51, 36, 20, -64, 14, -25, -15, 70, -15, -23, 18, 29, 7, -22, -9, -3, -35, 18, -30, -29, 52, 13, -7, -15, -29, 22, -24, 26, -31, 15, 8, 77, -109, 6, -24, -37, 70, -44, 27, 1, 17, 3, -13, 14, -85, 44, -32, -25, 27, -64, 60, -1, 62, 3, -25, 54, -30, -34, 1, -117, -7, 11, -3, 65, 13, 35, -4, 12, 17, -88, -5, -58, 37, 8, 19, 36, -5, 39, -104, 15, -22, -79, 70, -2, 85, -25, -39, 0, -29, 21, -53, 102, 19, -3, 52, -108, 59, -2, -6, -3, 46, 34, -72, 42, -54, -8, -2, -45, 13, 63, -75, 31, -38, -2, 24, -43, -56, 35, -17, 7, 25, 61, 29, 56, -15, 15, 31, -71, 12, -26, 34, -35, 14, 29, 8, 25, 1, -24, -12, -46, -40, -5, -64, 32, -43, 6, 88, -9, -15, 54, -26, -13, -7, -79, 0, -26, -24, 28, 12, 80, 51, -7, 5, -19, -20, 13, -13, 9, 25, -18, -30, 80, -42, -8, 5, 51, 54, 4, -6, -8, -36, -39, 2, -27, 70, 7, 0, -66, -21, -65, 22, -47, 57, 72, 47, 14, -8, -3, 11, 0, -10, 44, -39, 10, 35, 28, -12, 31, 23, 34, -117, -1, 2, -7, 2, 55, -29, 93, -87, 6, 26, -76, 88, -3, -31, 35, -11, -10, 26, -17, 46, -49, -1, 72, -35, 46, -56, -21, 28, 34, -62, -21, 10, 75, 0, 23, -19, 71, -35, 14, 17, -83, 27, -53, -18, -39, 15, 19, 2, 75, -4, 49, -4, -29, 49, -79, 108, -27, -24, -21, 37, -11, -11, 2, 18, 48, -12, 34, -68, -4, -48, 0, -30, 29, -27, 18, -41, 12, 23, -54, 26, -6, 48, 29, -37, -4, -1, -56, 2, -1, -49, 39, -36, 94, -58, 52, -90, 87, -6, -40, 2, -23, 62, 14, -27, 18, 54, 34, 1, -48, 22, -18, -55, -49, -47, -27, 0, -31, 75, 41, -5, 24, 3, 42, -65, -52, 102, 3, 5, 8, -10, 37, -62, -9, 54, -19, 15, -82, 31, 3, -17, 48, -23, 10, 107, -48, 10, -6, -25, -7, -15, 0, 22, -5, 21, -34, 73, -61, 59, -88, 38, 3, -15, -36, 22, 6, -2, 21, 6, 64, 23, -5, -29, 35, 7, -63, 27, -43, 20, 11, 83, -4, -2, -32, -25, -19, -4, -28, 64, 0, 12, 6, 17, 44, -24, 24, -79, 37, 51, -14, -8, -9, 81, 21, 34, -13, 34, 20, -14, -39, -36, -32, -65, -11, 12, -55, 66, -61, -12, 37, -64, -24, -8, -62, 96, -39, 26, 44, -43, 38, -39, 52, -69, 45, -69, 21, 71, -20, 4, 71, -57, 38, -13, -34, 11, -20, 31, 32, -85, 4, -8, 51, -6, 0, -21, 18, -40, -14, 29, -91, 62, -34, 79, -53, -13, 51, 0, 22, -78, 13, -54, -37, 21, -37, 24, 43, -27, 25, 13, 22, 17, 1, -13, 30, -30, -22, -27, 44, 0, 30, 56, 58, -46, 11, -56, -64, 39, 6, 12, 18, -23, 26, 3, -10, 51, 51, 74, 29, 2, 38, -18, 37, -18, -61, 3, -68, -14, 29, 17, 35, 0, -3, 21, -66, -11, -54, 17, 49, -17, 0, 70, -74, 18, 22, -63, 38, 10, -31, 17, 1, -14, 22, -68, 37, -39, -21, -64, -21, 20, -22, 15, 12, 7, 22, 71, -66, 19, -56, -52, 10, 14, -47, 3, -79, 52, 9, -54, 19, 32, 64, -42, -37, 23, -9, -40, -29, 53, -9, 47, 12, 6, 26, 59, 53, 37, -8, 5, -20, -45, 1, -92, 107, -44, 34, 48, 1, 44, -98, 47, -32, -37, 109, -34, 42, -20, 44, 6, -81, 3, -36, -86, 49, -2, 20, -1, 9, -4, 51, -57, 69, -10, 56, -60, -1, 21, -52, 98, -8, 31, -48, 54, -29, 15, 9, -8, 72, -24, -62, -4, -4, 27, -40, 77, -70, 8, 0, -57, 45, 10, -30, 32, -23, -45, 51, -44, 24, 31, 45, 14, -28, 20, -59, -93, -36, -4, 20, -1, 59, -7, -36, 42, -48, 14, -8, -26, 66, -15, -72, -18, 29, -7, 55, 7, 11, -27, 0, 44, -30, 73, -25, 14, 35, -2, 7, -38, -10, -14, -38, -51, -1, -54, 39, 1, -35, -9, -53, -4, 25, -30, -58, 5, 11, 23, 12, 19, -46, 27, -35, 8, 8, -76, 62, -49, -10, 1, 14, 27, 17, -4, -47, 85, -32, -4, 25, -39, 58, 3, -32, 13, 41, -73, 82, -49, 29, 14, -32, 82, -58, -1, 87, -17, -10, 8, -26, 28, 42, -38, 15, 18, 27, 38, -45, -9, -3, -25, 9, 82, 28, 12, 12, 11, -31, -47, -28, -37, -5, -15, 25, -11, -4, 28, -91, -4, -5, -28, -53, 60, -23, 97, 4, 14, 0, -20, 38, -26, 42, 10, -17, -22, 2, 6, -51, -4, 53, 30, -19, -53, 24, 46, 24, 18, -9, -41, -18, -11, 12, -61, 59, 21, 0, -1, -77, -3, -11, 13, 25, 34, -31, 2, 41, -5, 2, -36, 58, -34, 41, -32, 30, 48, -54, 36, -59, 24, 15, -24, -22, 73, 3, -25, 78, 29, -89, 41, -40, -62, -35, -19, 57, 7, -28, -38, 17, 0, -10, 28, -18, 27, 26, -73, 54, 7, -14, 43, -30, 0, -3, 0, -57, 65, -53, -12, 64, -7, 44, 43, -30, 31, -26, 30, -124, 79, 21, -35, 49, -72, 8, -3, -44, -10, -59, 51, 3, 10, 60, 34, -14, 58, -32, 18, -32, -26, -26, -12, -26, 26, 32, -5, -51, 36, -13, -31, 0, -72, 81, 58, -30, 8, -10, 6, -10, -57, -21, 28, -1, -24, 22, -37, 49, -23, -19, 28, -11, -68, 8, -59, 7, 60, -9, -9, 30, -62, 27, 4, -34, 58, -5, 49, -29, -11, -10, 11, -8, 83, -30, -37, 8, 21, -71, 90, -14, 7, 69, -64, 7, -62, 5, -46, 71, -17, -18, 61, -39, 18, 0, -56, 0, 46, -24, -47, -15, 51, 14, -35, -5, 19, 8, -56, 54, -13, -18, 35, -41, 89, -42, -15, 83, -73, 103, -22, 0, 94, -82, 15, -46, -29, -21, 11, 58, 34, 8, 14, 42, -44, -35, -60, 60, -3, 7, 28, -55, 59, 6, -85, 69, -47, -17, -20, -49, 71, -25, 57, -22, -31, 77, -62, 72, -4, 4, 70, -37, 70, -32, -11, 2, 58, -29, -26, -19, -9, -8, -6, 38, -54, 62, 0, -57, 65, -64, 75, -31, -43, 27, -5, 5, -57, -34, -12, -21, -22, 31, -3, 11, 25, 38, -39, 22, -11, -26, -49, -58, -7, -11, -17, 26, -10, 25, -68, -4, 5, -38, 59, 36, 36, -25, 36, 1, 12, -45, -32, 22, 66, -6, -22, 28, -6, -32, 0, 0, 32, -39, -56, -18, -18, -43, -11, 52, 43, 10, -38, 17, -40, 64, -7, 29, 41, 64, -20, -32, -53, 8, 34, -6, -2, 15, -52, -28, -22, 53, 4, 1, 4, 30, -22, -57, 1, 14, -10, -43, 42, -37, 73, -23, 26, -62, 28, 55, -8, 18, 64, -58, 12, -43, -61, 26, 3, -12, 77, -38, 24, -1, -61, -24, 63, 8, -15, -10, -52, -10, 13, -69, 79, -20, 28, 76, -13, -5, 25, -3, -14, -2, -53, -23, -4, -3, -34, 77, -9, -79, 31, -37, 13, 29, -22, -4, 58, 52, -8, 9, 22, -52, 28, -5, -77, 12, -5, 15, -29, 3, 19, 17, 35, -42, -17, 28, -25, 23, 25, -31, 58, -21, -13, 28, -41, -11, -7, 24, -52, -48, 51, -47, -4, 20, 19, 37, 5, -5, 91, -48, -14, 78, -38, 47, -26, -29, 28, 21, 0, 39, 1, -19, 40, -10, -35, 23, 46, -6, 39, -46, -36, 7, -30, -5, 23, -3, 35, 20, -58, 43, 20, 32, 22, 42, 83, -42, -25, 4, -30, -20, -71, 2, 27, 14, -20, -1, 20, -8, 65, -46, -20, -39, -64, -19, 10, -3, 48, 0, -8, 0, 7, 18, -17, 43, 26, -60, 25, 15, 12, 11, -14, 69, -5, -60, 39, -30, -21, 39, -48, 45, 12, -12, 39, -3, 18, 23, 69, -42, 45, -36, -48, -61, -42, -22, 20, -13, 31, 74, -59, 1, 17, -6, -100, 36, -20, -18, -13, 60, -22, 78, -41, -14, -19, 4, -2, 45, 11, -20, 15, -8, -59, -27, -78, 34, 44, 18, -10, -27, 8, -49, 25, -31, 3, 73, 11, -19, 61, -51, -18, -58, -81, -10, 18, -21, 4, -21, 58, -44, 37, -22, -41, 39, -48, 59, -51, 43, -32, 20, 34, 19, 17, -26, 58, -24, -23, -30, 14, -52, -40, -42, 15, -17, 62, 75, 70, 11, 6, 7, -47, -23, -66, -8, 32, -82, 77, -21, 25, -5, 3, 48, -78, -30, -21, 0, 30, -52, -3, 47, -77, 85, -37, 37, 27, -21, 58, -56, 46, 45, -3, 61, -45, -20, 5, -11, -11, 49, 21, 1, 20, -11, -18, -3, 13, 44, -47, -41, 22, -15, 74, -45, -14, -2, -58, 63, -57, 70, 11, 34, 5, -35, 74, -20, 20, -28, 77, -4, 69, -39, 6, -17, -20, -28, 23, -52, -18, 12, 35, -40, 44, -6, 22, -29, -10, -63, 11, -30, 39, -24, -42, 61, 12, -15, -60, 19, -28, 29, -64, 9, 21, -55, 83, -30, 27, 3, 65, -13, 45, -20, 11, -36, -12, -32, -40, 30, -52, 1, 59, 42, 26, 37, -64, 52, 5, -32, -17, -32, -27, 30, -40, -21, 72, 11, 37, -8, 25, -22, 57, -10, -30, -17, -1, 23, -54, -10, 2, 76, -17, -47, 62, -86, 49, -12, -76, 48, -126, 90, 21, 45, 53, -12, 6, 1, -37, 19, -5, 36, -19, -25, -29, -68, 29, 11, 3, 0, 19, 12, -76, -2, 42, -13, -9, 40, -31, -43, 31, -4, 11, 15, -44, 66, 36, -12, -8, -25, 20, -38, -52, 2, -13, 72, -32, -14, -23, 14, 34, -10, 31, -25, 65, -17, -41, 68, -15, -37, -22, -61, 9, 25, -47, 13, 9, -24, 99, -44, 23, 57, -29, -24, -47, -42, 38, -9, 18, 68, 5, 49, -49, -21, -12, 0, -52, -29, -5, 15, -10, 25, 35, 2, -4, -47, 80, 8, 14, 23, -37, 5, -46, 55, -77, 63, -29, 0, 37, -62, 53, 5, -20, 36, 71, 3, -63, 15, -56, -9, 20, -44, 20, 41, 35, -17, 31, -57, 57, -22, -18, -21, 14, -20, -41, -8, -3, 61, -19, 57, -46, 41, -19, -88, 20, -24, -15, 4, -10, 21, 100, -28, 9, 26, -53, -74, -7, 5, -19, 0, 1, 5, 40, -70, -15, 28, 11, 76, 7, -2, 47, -11, -43, -44, -55, -49, -1, 14, 10, 29, -12, -1, -55, 34, -62, 76, -29, -40, 36, -78, 79, -27, 34, 4, 45, -25, 8, 35, -64, 40, 9, 23, 3, -5, -40, 85, 0, 17, 26, 27, 55, -57, -28, -27, 10, -3, 5, -23, 19, 15, -5, -13, -20, -34, 0, -51, 37, -49, 51, -46, 22, 4, -14, 110, -29, 0, 18, -51, -40, 7, 35, 0, 8, -29, 62, -11, -92, 38, -49, 75, -30, -26, 35, 57, -46, 4, -88, 40, 3, -51, 55, 19, 59, 11, -6, 51, -30, -12, 30, -15, 34, -2, -77, -53, -29, 43, -28, 40, 17, -24, 51, -65, 48, -11, 28, 55, -68, -2, 25, 49, -17, -28, 5, 10, 56, -49, 1, 61, -30, -12, -45, 39, 22, -65, 47, -44, 1, -7, 2, 26, -44, 36, -30, -36, -14, -27, 48, 38, 25, 0, 0, 27, -60, -40, -23, -6, 6, -53, 9, 92, -22, 14, 41, 57, -77, 55, -19, -18, 45, -43, 22, -28, -38, -20, -6, -1, -27, 0, -54, -74, 0, 44, -2, 21, -30, -1, -18, -9, 11, -62, -9, 42, -4, 27, -81, 24, -23, -59, 54, -8, 0, 56, -74, 27, -10, -78, 40, 25, 37, 20, -11, -4, -39, 59, -8, 20, 17, -53, 8, 8, 34, -23, -2, 9, -22, -12, -34, 6, 14, 12, 34, -2, 43, 20, -2, -77, 3, -11, 17, -40, 41, 8, 62, -36, -58, 8, -31, 6, -2, -54, 36, -107, 34, -1, -54, 58, -12, 81, 28, 11, -15, 3, -53, -35, -26, 15, -18, 25, 15, 56, -13, 2, 23, 37, -49, -17, -19, 3, 24, -37, -15, -49, -23, -12, 35, -13, 40, 14, 19, 46, -14, -14, 26, -43, -21, -22, -39, -39, 66, -45, -38, 68, -69, 74, -44, 1, 14, -20, 31, 3, 14, 1, -20, -17, -29, 81, -21, -8, 47, -96, 24, 37, -9, 62, -9, -39, -25, -3, 18, -30, 49, -46, 15, -4, 2, -39, -71, 87, -9, 14, -15, 28, 57, -73, 55, -89, 45, 21, -52, -23, -4, 35, -9, 12, 37, -36, 39, -35, 60, -69, -35, 0, 12, 36, -31, -32, 54, -47, -17, -17, -72, 56, 17, 14, 0, 14, -52, 85, -8, 31, 42, 29, -9, -22, 42, -57, 32, -75, 56, 1, -103, 43, -46, 72, -43, 13, 39, 44, 25, -29, -11, -36, -38, -24, 10, 11, -3, 22, 80, -81, 38, 18, -85, 48, -12, -22, 21, -52, 4, 6, -78, 18, -53, 81, -8, -15, -17, 56, -53, 25, 18, -35, 88, -78, 26, -23, 34, 28, -63, -3, -77, -42, 37, -10, 0, 21, -17, 63, -10, -13, -17, 42, -49, 96, -44, 15, -32, 1, -47, -8, 80, -26, -26, 39, -32, 44, 15, -28, 21, -42, 25, 27, -95, 8, -40, 6, -11, -14, -2, 61, -6, -23, 66, 14, -62, 72, -53, -45, 29, -17, -11, -45, 63, -22, 38, -46, 87, -62, -9, 29, -48, 15, 41, -45, 14, -35, 34, 10, -25, 0, 46, -53, 29, -5, -31, -52, 5, -7, -100, 108, -31, 15, 79, -63, 52, 6, -23, 93, -109, 45, -36, 49, 22, -74, 54, -71, 0, 13, -77, 54, 15, 4, 44, -57, -20, -45, -11, -36, 2, -68, 24, 60, -11, 27, 55, -85, -1, -58, -27, 48, 28, 4, -13, 43, -1, -29, -70, -2, -27, -38, 3, -18, 4, -4, -10, 18, -11, 12, -4, -19, 78, -15, 14, -29, 7, -73, 0, -52, -28, 48, -1, 51, -6, 73, -40, -9, 10, -13, 20, -69, 2, -25, -2, 8, -20, -11, -3, -30, -14, -26, 11, -55, 81, -54, 8, 4, -43, 6, 45, -14, -10, 62, -81, -8, 29, -24, -15, 80, -107, 38, -40, -73, 48, -66, 93, 15, 68, -11, -8, 14, 11, 44, -58, -5, 9, -10, -42, -32, 0, -32, -22, -10, 41, -29, 27, 87, -7, 10, -44, -10, 31, 0, 48, 26, 0, -29, 80, 10, -13, 29, -1, 46, -12, -54, -2, -24, -14, -56, -3, -12, 104, -53, -25, 8, -25, 30, -23, 1, -5, 42, -28, -9, 25, -26, 66, -19, 31, -10, 58, 6, 59, -66, 36, -56, -44, -29, -14, 47, -15, 20, -25, -42, -29, -60, 9, 11, 6, 15, 80, -40, 71, -51, -13, 47, -55, 87, -55, -39, 87, -77, 89, -13, 7, 55, -73, 6, 49, 34, 0, 9, -26, 9, -9, -46, 8, 6, 24, -43, 49, -64, 18, 34, -4, 64, -15, 20, 40, -43, 48, -99, 9, 43, -30, -12, 38, -19, 114, -18, 42, 6, -53, 37, -38, 55, -23, -21, 20, -32, -30, 24, -11, -20, 34, 69, -13, 8, -58, 2, -37, 38, 17, 25, 25, 22, 32, -57, 7, -38, 8, -36, -1, -1, -43, 23, 6, 9, 100, -9, -19, 0, -11, 48, -9, -9, 65, -32, 20, 8, -92, 14, 29, -31, 15, 6, 24, 24, 14, 10, -35, 38, -48, 53, -36, 24, 52, -62, -41, -47, -61, 3, -8, -29, 35, -43, 73, 36, -6, 20, 34, 37, -25, -22, -14, -41, 24, -59, 9, -21, 26, -1, 13, 71, -41, 12, 43, -6, 8, -25, 45, 5, -36, 47, 44, -13, -1, -79, 32, -39, 7, 29, 80, 41, 3, 1, -1, 38, -56, 23, 56, -1, -36, 64, 21, -53, 30, -59, 51, 9, 5, 6, -21, 17, -28, 2, -9, -59, 28, 64, -43, 19, 56, -6, 35, -52, 39, -55, -7, 82, -66, 27, -23, 20, 37, -36, -28, -26, -46, 38, 34, 10, 37, -25, 15, -32, -62, 34, -30, -4, 77, 5, 25, 28, -9, 3, -76, -56, -57, 2, -14, -27, 48, -58, 60, -56, 62, -41, -5, 74, 1, 64, 15, -44, 22, -32, -22, -3, 8, 4, 40, 10, -34, 6, 97, -36, 37, -18, -4, 40, -41, 91, -43, 13, 58, 4, 36, -56, 46, 4, -39, 10, -64, 30, 0, -37, 70, -69, 40, -93, 3, 26, 0, 73, 53, -10, 26, -9, -62, 15, -40, 35, -11, 0, 49, -72, -17, 13, -51, 74, -5, 62, -24, 29, 62, -49, 48, -46, -27, -27, -47, -42, -2, 54, -17, 21, 29, -5, 3, 20, 13, -41, 32, -9, -20, -20, 51, -78, 62, -91, 64, 9, -52, 25, -48, 43, 10, -41, 7, -3, -19, -23, 27, 34, 27, 1, -54, 10, -42, -24, 32, -62, 60, -51, 57, 12, -2, 42, 28, 10, -11, 5, 21, -9, -127, 3, -34, -20, -17, 57, 87, 30, -22, -26, 34, -5, -27, -23, -14, 77, -48, -27, 6, -4, 34, 3, 43, 17, 64, -1, 14, 63, -25, 55, -45, -38, 13, -48, -40, 90, 6, 37, -4, 0, 10, -14, 25, 43, -10, -55, 35, 32, -4, -41, 12, 42, -11, -49, -7, 40, -11, 52, -30, 10, -6, -28, -45, -44, 21, -63, -15, 7, 18, 37, 9, 43, 11, 70, -19, -17, 41, -113, 61, -19, -20, 54, -7, 17, -25, 42, -44, 99, -28, 2, 30, -41, 70, 5, -20, 42, -10, -29, -14, -24, 12, -19, -44, 69, 21, 1, 37, -9, -22, 14, -18, -31, 38, -60, -22, -37, 11, 8, -38, 40, -46, 87, -26, -13, 61, -58, 14, 120, -27, -24, 35, -49, 12, -42, -27, 76, 0, 19, -52, -24, -42, 15, -23, 23, 19, -54, 52, 17, -35, 14, 2, -22, -11, 30, -69, 59, -57, 34, 41, 10, -7, 11, -10, -32, -66, 37, -4, 6, 43, 64, 22, -6, -29, 6, -73, 28, 28, 17, 58, -19, 54, -37, 6, -23, -64, 8, 20, -36, 1, -27, 48, -25, -13, 63, -6, -31, 52, -20, 1, -6, 70, 48, 20, -57, 22, -48, -23, 17, -72, 70, -28, -2, -9, 15, 12, -38, 57, -63, 10, -48, 74, -34, 44, -59, 36, -1, -65, -41, 37, -31, 45, -25, 18, 32, -44, -28, -30, 29, -61, 36, -31, 20, 49, -34, -8, -7, 21, -17, -39, 7, 20, -76, 69, -26, 23, 73, -46, 32, -20, -18, -5, -22, 28, 56, 1, 7, 92, -116, 53, -29, -32, 5, -63, 43, -5, 15, -39, 30, 66, -48, 19, -5, -62, 32, 18, 28, -17, -13, -42, 8, -18, -40, 88, -18, 51, 7, -13, 86, -80, 1, 39, -40, 73, 1, 46, -27, 36, -5, -70, 38, -1, -28, 65, -89, 31, 44, -11, -34, 0, 41, -12, -18, -37, -23, -36, -1, 19, -31, 56, -27, 27, 21, -14, 17, 8, 23, -34, 22, -20, -5, 6, -71, 69, 3, -87, 44, -28, 10, 54, -24, 13, 51, -68, 42, -25, 0, -41, -28, -48, 22, -2, -46, 59, -90, -9, 19, -11, 47, -7, -3, 30, -32, 40, -17, 73, -5, 14, 4, -24, 11, -85, 94, -25, 57, -23, 1, 11, -13, -72, 35, -14, 29, 59, -12, 7, 35, -59, -20, -4, -28, 8, -108, 26, -30, 80, -6, 43, -19, -24, -15, -77, 63, -44, 29, 32, 18, 15, 24, 9, 14, 41, -10, 61, -37, 79, -25, 8, 56, -65, 92, -43, 2, -2, -4, 35, -20, -59, -3, -45, 6, -38, 61, -24, 14, 4, -1, -7, 0, 0, 36, -59, -2, 4, -12, 47, -8, 10, 9, -25, -7, -69, 60, -27, 31, 51, -46, 4, 41, -17, -55, 38, -74, 8, -36, -27, 68, -41, 51, -23, 31, 47, -24, 7, 0, 10, -59, 0, -6, 10, -19, 22, 40, 64, 62, 21, -25, 8, 0, -19, 17, -21, 18, 45, -40, 68, -51, -58, 15, -8, -43, 94, 2, 18, 32, 18, -37, -37, 35, 41, -17, -54, 19, -29, -30, -15, 0, 64, 0, 24, 24, -53, 92, -95, 66, -9, -1, 104, -64, -7, 14, 9, -66, 10, -41, -36, 103, -47, 34, -56, 20, 56, 4, 22, 32, -26, 7, -47, -45, 20, -8, 37, 52, 17, 19, -1, -26, 0, -4, -93, 54, 24, -43, 13, 65, -10, 22, -2, -45, 18, 7, -25, -35, 1, 4, -54, -63, 27, -17, 35, -48, -13, 49, -17, 41, -18, 22, -6, 61, 54, -28, -26, -8, -48, 24, 21, 15, 5, -43, 46, -15, -49, 57, -39, 57, -58, 49, 49, -29, -25, 23, -8, -83, 41, -37, 30, 0, 73, 41, -3, -6, -59, -9, -28, 51, -62, 0, 22, -14, 46, -20, -2, 9, -4, -5, -39, 48, 30, -61, 83, -115, 14, -37, -90, 82, -42, 38, 42, 56, 4, -19, -5, 37, 32, 41, 49, 5, -14, 27, -10, -35, 39, -83, 17, -11, 30, -64, 2, -1, 8, 19, -7, -4, -4, -39, -10, 43, -14, 37, 9, 2, -99, 22, -14, -11, -8, -17, 63, -43, 45, 15, -51, -13, 0, -21, -18, 71, 28, -24, -10, 31, 10, -44, 2, 75, -49, 51, 31, -74, -37, -12, 21, -5, 59, 4, -32, 18, -37, 30, -2, -13, -65, 72, 6, 15, -35, -8, 31, 14, 62, -2, -57, 53, -55, -2, 9, -47, 72, -57, 13, 24, -13, -66, 95, -45, 23, 32, -56, 14, -10, 25, -23, 15, -49, 69, -26, 6, 28, -14, 40, -15, -41, 87, -34, -31, 62, -8, -8, -17, 15, -57, 83, -68, 42, -2, -60, 70, -14, 47, -59, 10, 9, 12, 15, -22, 35, -36, 69, -18, -64, 44, -31, 5, 25, 19, -22, -27, 13, -30, -1, -4, -15, 5, 2, 2, -55, -19, -23, 22, 18, 57, 37, -45, -4, -53, 2, 3, 2, 18, 47, 1, 18, 6, -8, 17, -3, 31, -2, 24, 0, -36, 40, -43, 20, 46, 32, 79, 49, -5, 31, -62, 0, 14, -32, 1, 5, 88, -13, -37, -6, -31, -5, -4, -41, 49, -29, 24, 68, -9, 36, -73, 28, -9, -29, 72, 11, 8, -38, 55, -60, 81, 4, 25, 45, 3, 27, -100, -6, 34, -10, 29, 52, 3, 2, -32, -55, 9, 24, -52, -31, 55, -56, 94, 0, 22, -29, 57, -2, 9, 14, -14, 22, 11, -69, 22, -21, 15, -29, -23, -8, -44, 2, -26, -13, 45, 62, 54, 24, -26, 21, -49, 34, -6, -21, 20, -51, -2, -9, 3, 4, -76, 71, 32, -40, 60, -49, -3, -19, -47, -6, 22, 2, -4, 117, -57, -27, 12, -31, -17, 26, -58, 25, 31, 27, -53, -15, -21, 5, 20, -2, 10, 43, 53, -27, -6, 28, -30, -63, -12, -3, -10, -7, 26, -73, 25, -65, -11, 11, -107, 35, -30, 32, -14, 23, 12, 81, 1, 54, 11, -29, 63, -44, 13, -77, 42, -20, 57, -30, -18, 56, -48, 56, -41, 102, -10, -26, 26, -52, -34, -5, -31, 12, 85, -69, 19, -9, 2, 11, -57, 38, -65, -57, -13, -1, 30, 2, -7, -34, 19, -36, 54, -26, -32, 21, -17, -73, -28, 7, 2, 36, 7, 20, 76, -13, 14, 19, -29, -3, -58, -17, -87, -2, 11, -59, 79, -58, -34, 55, -9, 1, 9, -7, 65, -23, -7, 74, -34, 0, 79, -12, 28, -3, -91, -2, -30, 6, -47, -30, 97, 2, 30, 54, -54, 76, -8, -9, -18, -60, -62, -56, -28, -6, 17, 51, 32, 0, -7, 25, -7, -10, 38, -57, 52, -12, 55, -24, 1, -7, 1, -28, -4, 7, 5, -22, 32, -9, 75, 11, -4, 7, 11, -58, -20, 45, -39, 49, -88, -8, -11, -46, 69, 0, 27, -36, 29, 19, 11, 44, -24, -7, 24, -34, -13, -9, -6, 37, -22, 20, 48, 48, -35, 2, -17, 0, -6, -13, 6, 0, 43, -44, -7, 24, -91, 59, -11, 41, -5, -6, 116, -69, 36, -4, -56, -17, -37, 47, 2, 5, 8, 75, -29, 47, -14, 24, 41, -45, -4, 49, -2, -39, 60, -14, -52, 27, 4, -1, -49, 53, 2, -92, -31, 14, 7, -21, 31, -62, 24, -43, 24, -20, 6, 17, -13, 74, 3, -13, 11, 0, 63, -42, -3, 3, 32, -55, 25, -9, 6, 37, -85, -23, -44, -57, 54, -30, 28, 24, 5, 76, -53, -23, 63, -54, -14, 76, -5, 61, -11, 26, 55, -85, -1, -20, -23, 13, 0, -76, 78, -60, 6, 9, -39, 99, -19, 3, 27, 0, -24, 45, -22, 3, 29, -10, 18, -21, -59, 43, 26, -23, -35, 24, -7, 13, -37, 0, 29, -69, 63, -93, 41, -10, 36, -21, 54, 52, 14, 46, -66, 18, 2, -44, -46, 35, -12, 57, -13, 4, 54, 31, 46, -63, -20, -15, -31, -21, 11, -28, 31, -5, 59, -5, 89, 4, -65, 1, -35, 34, 3, 41, -32, -3, -22, 27, -26, -15, 18, -70, 22, -42, 42, -32, 7, -31, 21, 17, -17, 53, -56, 75, -78, 11, 5, -44, 34, -3, 62, 27, 68, 13, 22, -45, 6, 7, 44, -96, 20, -38, -12, -13, -46, -69, 32, 2, -38, 81, -8, -2, 66, -24, 23, 30, 17, -28, 10, -23, -55, -18, 21, -28, 31, 39, 23, -24, 88, -81, 23, 23, -7, 4, 44, -9, -11, -10, -42, -24, -8, -30, 37, -22, 49, -24, 14, 5, -21, -29, -56, 0, -20, -14, 45, -15, 29, 38, -46, 6, -6, -3, -89, 30, -85, 42, -36, 32, 54, 36, 37, 5, 25, -52, -54, -82, -4, 39, -45, 19, -34, 38, 19, -4, 64, 36, -39, 19, -21, 31, -37, 9, 38, -27, -70, 44, -1, 4, 39, -30, 100, -69, 32, 52, -116, 10, 5, -42, 43, -31, 56, 24, -3, -27, -21, -41, 0, 15, 26, 19, 20, 80, -58, 21, -29, 10, 7, -79, -35, -57, -37, 4, 13, 54, 20, 8, 4, 34, -47, -11, 28, -34, 24, -55, 23, 32, -81, 21, 61, 5, 4, -45, 78, -72, 81, -18, 9, 36, -34, 45, -47, 26, 12, -47, 60, -64, 32, 3, -38, -35, 63, 10, 3, 81, -94, 0, -89, -24, 4, -4, 18, 42, 23, -6, 71, -38, -41, 48, -23, 7, 45, -17, 29, 29, 32, -34, 3, 47, -112, 17, -5, -8, 88, -15, -6, 46, -44, 22, -37, 1, 12, 47, -3, 2, -9, 6, 31, 12, -81, 19, -43, -6, 52, -70, 12, -43, 24, 2, 9, 59, -31, 21, 47, -74, 35, -53, 37, 26, -68, 76, -49, 9, -10, -105, 8, -38, 13, -52, 21, 63, 53, 6, 2, 45, -24, -66, -42, -17, 18, -34, -11, 81, -29, 57, -21, -22, 40, -42, 61, -10, 71, -18, 31, -30, 27, -24, -72, 13, -26, 28, -30, 30, 37, -30, 26, 64, -47, 23, -34, -35, -14, -28, -39, -29, 0, -7, 35, -57, 10, 49, -22, 41, 11, -21, -18, -1, -74, 82, -44, 56, 13, -20, 20, -57, 14, 19, -25, 12, -96, 29, -2, 3, 18, 37, 22, 34, 61, -4, 9, 0, 25, -5, 24, -46, 9, -55, 12, 7, -5, 68, -15, 20, -43, -55, -29, 17, 18, -62, 8, -62, -19, 40, -30, 71, 29, 12, 25, -18, -24, 14, -69, 3, 24, -51, 24, -58, 56, -73, 31, -6, 25, 80, 13, 11, -3, 10, 108, -6, 22, -17, -23, -11, 5, -42, 14, 3, 35, -13, -39, -30, -49, -8, -69, 18, 20, 3, 19, 72, 47, 73, 29, -51, 12, -35, -30, -28, 20, -37, 42, 7, -8, 25, -44, -1, 57, 0, -26, 20, 0, 37, -45, 19, -25, 21, -31, 27, -62, 42, -62, 52, -3, -39, -47, 52, -26, 22, 52, 31, 19, -5, -14, -56, 21, 27, 15, 20, -19, 8, -5, -3, -29, 105, -65, 29, -80, 1, 9, -56, 43, 10, -7, 114, -52, -3, 30, -75, 66, -29, 60, 31, 12, 46, -62, 6, -7, -40, -58, 47, -106, 79, -48, 29, 102, 17, 39, 0, 52, -18, -52, -32, -25, -56, -35, 78, -22, 11, -40, 45, 31, -38, -11, 14, 28, -30, 61, 65, 28, -22, -36, 6, 20, -22, -39, 9, 26, 13, -48, 13, -20, 70, -18, 80, -30, -13, -12, -53, 13, 3, 35, 29, -10, -5, 14, -102, 78, -1, 9, 11, 54, -45, 24, 6, 0, 42, -2, -55, 98, -106, 102, -38, 29, 109, -49, -5, 38, -11, -25, 0, -23, -35, -79, -26, 48, 1, -9, 6, -5, 32, -19, -7, 62, 19, 17, -54, 8, -44, -32, 12, -104, 48, 14, -18, 34, 32, -23, -24, 19, -40, 14, -85, 102, -9, 49, 43, -51, 46, -68, -39, -20, 24, 14, -81, -2, 1, 29, -31, -42, -13, 40, -4, 27, 73, 21, 29, 3, 2, 32, -45, 27, -15, -85, 8, 29, -13, 82, -30, 17, 9, -38, 21, -90, 40, -41, 60, 40, 23, -7, 32, -4, -100, -25, -21, 41, 32, 54, -7, -4, 14, 11, -2, -31, 56, -10, -19, 22, 11, -45, -42, -14, -8, 42, -6, 68, -44, 57, -64, -21, 41, -24, 15, -24, 25, -32, 19, -12, -13, 61, -46, -9, -46, 54, 29, -18, 0, 99, -61, -4, -36, -56, 21, -52, 57, -69, -36, 38, 23, 0, 20, 53, -45, 49, -20, -14, -32, -9, 22, -42, 80, -39, 41, 79, -93, -4, -23, -23, 34, -13, -68, -7, -49, 45, -24, 48, 13, 26, 54, -105, 5, -35, -32, 14, -29, 7, 37, 29, -11, 34, 53, 9, 56, 2, 40, -69, 42, -2, -73, 37, -42, -25, -23, -25, 39, -63, -15, 75, 0, -2, 59, -42, 74, 15, -26, -41, 40, -1, -53, -32, -15, -4, 2, -11, -35, 35, -72, 93, -40, 42, 15, 47, 37, -35, 40, -31, -26, 21, -12, -7, -18, -19, 35, -15, -10, 78, -36, 48, -27, -35, -5, -6, 0, 24, -6, -10, 29, -31, -2, 38, -98, 11, 19, -19, -5, -12, -40, 17, -39, 17, 58, -8, -11, 15, 46, 31, -7, 10, 68, -23, 38, -94, 23, 13, -41, 15, -37, 86, -42, 32, 27, -34, 15, -60, 20, 6, -6, 62, 26, 48, -15, 24, 54, 18, -11, -8, -39, 23, -21, 40, 21, -38, 35, -73, -32, -30, 20, 8, 17, 17, 23, -6, 103, -15, -43, 13, 10, -44, -2, -40, 35, 7, -35, 36, -9, 8, -54, 3, 26, -51, 94, -15, -3, 15, -6, 0, 22, -52, 31, 15, 44, -28, 5, 17, 14, -64, 12, 1, 10, 27, -1, -21, 4, 0, -4, -29, -44, 27, -42, 48, -10, -14, 26, -71, 64, -14, -25, -3, 80, -26, 43, -9, 3, 11, -78, 43, -43, -20, 5, -2, 4, -56, 51, 30, -18, 29, -2, 40, -10, 9, -32, 70, -42, 0, -28, -2, -15, -68, 36, -80, 71, -38, -13, 29, -21, -28, 5, 19, -10, -14, 17, 23, 29, 6, -17, 18, 20, -73, 102, -46, 10, 3, 7, 9, -55, 59, -60, 90, -55, -10, 17, -92, -27, 8, -8, 34, -17, 14, 72, -83, 20, 4, 75, -28, -6, 21, 46, -45, 4, -1, 10, -28, 23, -27, 65, -24, 14, 2, 99, -49, -46, 14, -41, -8, -64, 1, 52, -17, 80, -42, -9, -31, -25, 9, 12, -20, 36, 58, -26, 64, -72, 68, -32, 10, 17, -29, -58, -26, 1, 3, 52, -13, 41, -22, 69, -17, -69, 10, -2, -36, 7, 31, -47, 60, -88, 46, -13, -28, -53, 61, -60, 71, -5, -21, 49, -51, 20, 85, -24, -22, 2, -3, 9, 32, -21, -10, 10, 22, 1, -6, -4, 60, -71, 9, 29, -26, -2, 53, -17, 29, 32, -19, 43, 6, 57, -73, -8, -27, 43, 4, 14, 52, -39, 56, 52, -64, 26, -35, 21, -42, -14, -36, -32, 7, -91, 44, -46, 79, 23, 26, 22, -24, -26, -11, 4, -21, -1, 42, -55, 31, -5, 60, -23, -22, 49, 21, 0, -11, 32, 48, -59, 35, -35, -58, -35, -46, -13, 9, 46, -21, -36, 31, 19, -78, 79, -22, 5, 13, -70, 28, -23, -8, 22, 59, -30, -5, 44, -17, 24, -40, 109, -13, -23, 25, -47, 26, -26, 19, -91, 4, 13, 6, 30, -19, 35, -58, 9, 29, 2, 12, 18, -24, -20, 22, -83, 7, -17, -24, 88, -8, 22, 20, 10, -53, 53, -25, -63, 31, -54, 0, -38, 76, -11, 13, -3, -3, 66, -21, 36, -59, 13, 23, -56, 39, 4, 23, 44, -14, 66, -45, -61, -34, -61, 34, -57, 64, 49, 7, 52, -41, 74, -23, -39, 51, 8, -35, 10, 42, 0, -57, 21, -17, -61, 20, -58, -4, 34, -21, 62, -88, 38, -40, 3, 32, -41, -9, 39, -4, 10, -42, -30, -12, 21, -31, 74, -23, -17, 62, 6, -27, -24, 31, 35, -36, 7, 68, -36, -63, 15, 28, -37, 37, 68, -64, -9, 35, -42, 73, -13, -11, 35, -94, 71, 19, -43, 11, 27, 51, -4, -54, 37, 1, -51, 60, -41, -22, 105, -22, 1, 71, -91, 15, 10, -40, 10, -26, 58, -14, 8, 36, -29, 60, 10, -102, 1, -63, 38, -21, 43, -12, -45, 43, -19, 6, 41, -2, 44, 2, -44, 74, -71, 60, -34, 30, 48, -42, 21, 55, 52, -49, -17, 17, 31, -9, -38, 42, -30, 18, 39, -80, -5, -81, -4, 35, -69, 68, -19, 18, -7, -92, 97, -1, 20, 40, -13, 98, -27, -32, 9, -22, 32, -47, 52, -80, 22, 1, -45, 87, -14, -17, -11, 9, -20, -53, -29, 7, 10, 36, -43, -17, 40, -2, 49, 42, -42, 23, -54, -18, 32, -57, 82, -114, 0, 8, 34, -24, 19, 35, 41, -4, 3, -61, -28, -47, -22, 38, -43, 43, -71, 22, 19, -20, 31, -20, 21, 53, -19, -20, -22, 20, 8, -12, -44, -9, 71, 17, 57, 12, -1, 3, -30, -45, -24, -42, -1, 30, -77, 30, 9, 9, 6, -24, -27, -21, -29, 6, 46, -52, -25, -18, 6, 2, -19, 51, -27, 18, 44, -28, -9, 0, 11, -32, -10, 11, -62, -56, -13, -13, -6, 7, -3, 81, -7, 29, 13, 6, 8, -55, 2, -56, 104, 0, 37, -30, -19, 8, -19, 15, -18, -44, 61, 41, -2, 23, -19, 10, -62, 35, -68, 42, -26, 24, 34, -7, 42, 19, -19, 41, 7, -40, 19, -34, 13, -56, 0, 57, -38, 9, 20, 3, -39, 32, 0, -26, 59, -42, 7, -53, -73, -45, -43, 2, -38, -19, 82, -40, -25, 57, 55, -14, -13, 54, -85, 3, -48, -15, 45, -15, 66, -49, 32, -21, -66, -20, 10, 0, -2, -18, 7, -39, 0, 27, 5, 44, -8, 30, 20, -15, 37, 32, -69, -2, 5, 3, 0, -73, 54, -5, 15, -26, -21, -2, -27, 36, -92, 65, -27, -2, 53, -80, -32, -19, 27, 0, 7, 27, -64, -1, -17, -28, 63, -63, 37, -35, -11, 7, -18, 55, -20, -20, -10, 59, -68, 39, -42, -39, 51, -20, 42, 49, 17, 54, -44, 23, -73, 30, 20, -44, 8, 5, -32, -26, 22, 0, 53, 4, -47, 34, -56, 48, -19, 7, 18, -14, 13, -63, 2, 35, 51, -15, -73, 10, -47, 3, 15, 15, 22, -45, 55, 15, 34, -26, -12, 46, -32, -11, 14, -6, 51, -60, 45, 45, -73, 65, -35, -40, 9, -63, 7, -12, -77, 58, 31, -38, -48, 74, -62, 35, -35, -17, 75, -51, -18, 88, -25, 58, 1, 26, 27, -3, 12, -3, -63, 0, -15, -22, -21, 27, 13, 10, 73, 2, -46, 5, -14, -60, -59, 24, -46, 54, -14, 54, 10, 35, 41, -15, 32, -30, 2, 70, -58, 17, -35, -17, 41, -9, 23, 36, -26, 69, 11, -4, 28, -56, -21, -34, -59, 15, -17, -26, 44, -8, 60, -68, 12, -38, -22, -44, -26, 10, -29, 81, -53, 41, -24, 37, 35, -57, 13, 30, -8, 15, -34, 47, -58, -10, 2, 48, -18, 48, -66, 29, -52, 47, -59, 22, -18, 49, 1, -42, 38, 15, -51, 77, -75, 28, 55, 57, 51, -9, 19, -34, -28, 11, -49, -8, 12, -78, 61, -15, -43, 58, -34, -28, 32, 20, 49, -21, -38, 40, 24, -47, 97, -6, -54, 27, 1, 17, -49, -43, 27, 0, -58, 63, -18, 127, -51, 6, -8, -12, -6, -45, -20, -34, 0, -19, -68, 39, -28, -14, -29, 59, -12, 22, 56, -63, 41, -78, 24, -31, 3, 8, 65, 11, -22, -30, 22, -12, 42, -54, 2, -29, 41, -31, 32, 56, -31, 0, 5, 6, 14, -25, 28, -64, 24, 17, -45, 11, 29, 22, -21, 0, -76, 4, -25, -4, -7, 31, 19, -26, 9, 41, -21, 2, 37, -28, 53, 18, -26, -2, 0, 97, 3, 6, -10, -5, -61, 1, 0, -10, -35, 28, 52, 39, 11, -34, 9, -43, -10, 2, -22, 20, -15, 77, 8, 31, 38, -43, 2, -47, 74, -38, 5, -7, 52, 11, -22, -34, 62, 18, -56, 29, 30, -64, 105, -64, -38, 60, -76, 48, 45, 19, 12, -35, 41, 8, 0, -46, 32, -44, 47, 15, 23, -10, -28, 38, 29, -4, 4, 7, -19, 45, 22, -43, 32, 10, 3, 25, -61, 28, 32, -97, 54, 12, 7, 65, -37, -6, 25, -65, 39, 14, -2, -5, -70, 8, -4, -14, -36, 73, 36, -27, 70, -74, 57, 11, -58, 56, -25, -24, 10, -4, -23, 60, -82, 23, 25, -40, 75, -79, -18, 24, -28, 56, -14, -40, 82, -61, 0, 12, -37, 87, -93, 8, -27, -63, 63, 10, 40, -4, 0, 44, -54, 7, -49, 44, -21, 26, 7, -2, 46, -3, 38, -60, 26, 17, -90, 65, -64, 96, -34, 49, 51, -6, 0, -54, -21, -37, -2, 0, -24, -6, -43, 11, 14, -17, 0, 0, 23, 9, -77, 63, -38, 0, 53, 13, -30, 24, -51, -10, -53, -36, 68, -32, 38, 65, -70, 37, 27, -15, 37, -68, 24, 21, -79, 42, -62, 41, 14, -39, 12, -5, 60, -35, 47, -17, 0, -56, 42, 30, -62, 54, -10, -24, 62, -52, 76, -65, -46, 3, 1, 11, -49, 20, 40, -20, -63, 0, -55, -10, -1, -9, -23, -48, 11, 9, -38, 28, 29, -13, 51, -9, 6, 40, -35, 80, -74, 61, -4, 11, 0, -62, 17, 1, 40, -28, -3, 11, 6, 105, -60, -17, 35, -10, 22, -82, 55, 13, -87, -15, -24, 6, -13, 40, 25, 92, -34, 11, 32, -49, 25, -44, 25, -47, 17, -94, 69, 1, 37, 28, 5, -31, 7, 12, -5, 24, 0, 73, -99, 25, 34, -34, 69, -44, 2, -15, -7, -43, 34, -39, 39, 6, 46, -37, 59, -17, -18, -59, -39, -36, -27, -11, -43, 59, -27, 37, 31, 48, 32, 47, -20, 68, -10, -32, 19, -12, -77, 36, -76, 45, -43, 39, 53, -12, -60, 56, -25, -31, 15, -49, 59, -74, 51, -20, -38, 6, -18, -22, -75, 92, -40, 17, 18, 4, 46, -42, 59, -57, 45, -8, -37, -42, 20, 18, 1, 19, 8, 40, 30, -51, 17, 6, 7, 12, -14, -31, 35, -60, 11, -42, 8, 49, -19, 15, -43, -19, 44, -12, 57, 22, 66, -48, 52, 36, -70, 82, -53, 77, -78, -2, 42, -15, -41, 19, 66, -28, -17, -10, 31, -12, 9, -52, 10, -14, -42, 103, 10, -2, 36, -21, -5, 37, -97, 41, 8, -66, 63, 10, -55, 17, 12, -52, -14, -13, 74, -24, 18, 28, -8, 37, 6, -85, 10, -9, 6, -40, -6, 6, -76, 45, -9, 75, 54, 11, -17, 38, -34, 46, -60, 8, 21, -3, 27, -61, 15, -32, -24, 18, -15, -66, 27, -52, 71, -45, 9, 85, -97, 54, -14, -29, -31, -39, 54, 32, -51, -28, 28, -25, -10, -5, -10, 3, -96, 31, 29, -15, -2, -56, 75, 11, 11, -20, -60, 42, 11, 40, 1, -36, 43, -39, -29, -14, -71, 12, 6, -10, 43, -22, -23, 15, 15, 9, -25, 69, -59, 20, 42, -32, -30, 10, -39, 8, -92, 82, -54, 77, 9, 19, 40, 35, -28, 24, -115, 9, -29, 38, 17, 19, 80, -32, -2, -32, -42, -12, -25, -77, 25, -22, 6, -41, 115, -30, 26, 49, -49, 24, -8, -21, -12, -62, -54, -41, -10, 9, -17, 30, -2, 34, -10, -46, 30, -83, 21, -46, -4, 26, 11, 72, -14, -48, 65, -22, 18, -23, -36, 59, 0, -2, 69, -64, -51, 32, 17, -44, 32, -17, 51, -41, 14, 19, 40, -53, 9, -23, 36, 61, -1, -13, -9, -34, -9, -24, 44, 2, 20, 42, -39, 66, -69, 34, 68, -29, 24, 35, -9, 4, -21, -30, -42, -44, -24, -28, 19, -66, -37, -22, -2, -15, 51, 1, 0, 41, -95, 49, -13, 5, -51, 7, 68, -18, 2, 15, 12, -14, -9, -22, 36, -25, 69, -32, 23, 37, -22, -60, -62, -29, 26, -27, 53, 45, 53, 13, 42, 20, -81, -1, -12, -6, 9, -11, -8, 40, 71, -42, 7, -3, -55, -42, 4, -29, 73, -36, 15, 25, 30, -99, -20, -8, -48, -18, 6, 24, 54, 58, 24, -9, 79, -69, -44, 5, -38, 52, -12, 0, 51, -25, 37, 23, -13, 18, -9, -23, -46, -35, 41, -49, 70, 3, 34, 0, -20, 69, -19, -13, 38, -9, -13, -30, -27, 47, -8, 56, 23, 3, -46, 34, 62, 2, 5, -42, 11, 5, -12, 61, 56, 7, 1, -20, 14, -47, -21, 23, -1, 81, 28, 21, -15, -42, -55, -24, -12, -4, 30, 5, 36, 37, 58, -7, 22, 45, -87, 41, -43, -55, 97, -6, 26, -18, 6, -56, 15, -43, 46, 0, 2, 11, -43, 83, 0, 20, 2, -51, -1, -7, 15, -61, -25, 81, 5, 7, 18, -46, 62, -2, -44, 38, 8, -48, 76, -44, 93, -2, 5, 49, -86, 40, -81, 40, 14, 4, 73, 10, 14, 63, -48, 22, -49, 58, -47, 63, -36, 14, 87, 6, -55, 10, -38, -36, -2, -30, -11, 3, 12, -38, 69, -49, 48, -10, -35, 40, -18, -4, 27, 56, -51, -19, 21, -36, 45, -40, 52, 0, 124, -37, -39, 17, -12, -28, 29, -23, 8, 20, -69, -11, 29, -38, -29, -54, -6, 37, -17, 40, 12, 54, -41, 49, 0, -55, 88, -38, -65, 47, 1, 19, 9, -7, -6, -4, -3, -12, 103, -75, 5, 4, -21, 4, -82, 2, -21, -10, 36, 21, 24, 43, -20, -35, 56, -60, 79, -20, 55, 10, -29, 90, -75, 61, -19, -11, 13, -15, -17, 46, -52, 1, 61, 31, -34, -12, 21, -18, -55, -34, 4, -26, 23, -9, 61, 35, 2, 17, -8, 47, -37, 26, 6, 28, -34, -8, -54, 37, 21, -54, 5, 76, 8, -70, -19, -56, -51, -8, -14, 8, 36, 45, 30, -22, 40, -49, 0, -22, -5, -39, 17, -49, -6, -40, 6, -10, -30, -3, 55, -4, 13, 21, 46, -24, 35, -27, -70, 17, 2, -42, 49, 24, 47, 0, -37, -7, 34, 20, 22, 17, -41, -7, -10, 3, -68, 79, -59, 17, -15, 14, -10, 66, -19, -31, 77, -8, -1, 2, -70, -12, -49, 36, -44, 38, 34, -47, 62, -64, 10, 18, -66, 49, -10, -5, 62, -61, 36, -35, 15, 42, -28, 38, 20, -38, 97, -36, 27, -62, 11, 18, 12, -2, -19, 27, 14, -76, -17, -99, 1, 46, -1, 18, -31, 43, 0, 3, 6, -42, 37, -38, -8, 41, -89, 12, -3, -66, 69, -27, -27, 98, -65, 31, -40, -26, -14, 0, -62, 74, 20, 15, 13, -25, 72, 61, -26, -46, 6, 7, 13, -48, -8, -6, 20, 10, -24, 8, 27, 18, 30, -34, -10, 93, -9, 57, 1, 3, 29, -21, -6, -4, 40, -104, 34, -57, 48, -27, 53, 61, 48, -49, -24, -37, -22, 53, -9, -41, -17, -24, -6, 6, -3, 81, 30, 4, 64, -70, 0, -3, 2, -48, -2, -40, 0, 53, -1, 63, -35, 44, 17, -72, 9, -80, -9, 5, -26, 49, -30, 17, -53, 36, -49, 35, -51, 36, 1, -5, -41, 27, -37, -39, 53, 32, -9, -17, 57, -53, 31, -72, -7, -55, 55, -20, 36, 94, 8, -35, 40, -23, -21, -25, -20, 45, -43, -45, 15, -37, 5, 13, 59, -11, -5, 0, 2, -103, 31, 36, -47, 46, -41, 80, -20, -14, -6, 26, -15, -102, 10, -7, -31, 45, 78, -11, -11, 15, 0, -1, -57, -7, -19, -28, 46, 17, 8, 58, -69, 28, 10, -27, -41, 11, 1, 20, -54, 55, -22, -87, 20, -8, -4, -45, 42, 5, -4, 39, 6, 47, -37, -19, -56, 43, 39, -9, 21, 2, 90, -12, -41, 37, -52, -19, -57, 6, 48, -13, 14, -34, -2, -19, 30, -63, 29, -19, -58, 13, 20, -24, 10, 47, -52, -25, -5, 78, -45, 38, 7, -2, -21, -37, 23, 31, -30, 10, 87, -15, 12, -65, -2, -5, 41, -61, 43, 8, -59, -41, -6, 18, -68, 62, -103, 42, -19, 24, 24, -34, 60, -93, 71, -4, -12, 43, -58, 51, 24, -68, 52, -24, 5, -5, -65, -12, 1, 21, -19, 0, 60, -34, 13, 90, -19, 29, -34, -4, -58, -9, 8, -4, 26, -4, -15, 68, -31, -68, -34, 47, 40, 8, 46, -46, 48, 18, -36, 22, -32, -6, -43, -26, -34, 73, -43, -28, 22, -25, 23, -87, 6, 29, 12, 22, 43, -27, -42, 48, 27, -7, 45, 19, -5, -20, -30, -17, -9, -30, 0, 46, -25, -10, 7, -44, -15, -7, -15, -80, 38, -28, 53, -12, -27, 46, -76, 64, -38, 9, -19, 42, -4, -5, 63, 13, 26, -3, 23, -2, -7, 44, -77, 57, -106, 93, 3, 39, 59, -14, 40, -44, -27, -76, -20, -24, -4, 13, -28, 58, -30, 15, 40, -46, 27, -36, 59, 31, -39, 42, -62, -37, -46, -60, 91, -44, 53, -44, 34, 54, -70, 3, -38, 41, 8, 27, 31, 99, -61, -10, -61, -45, -1, -30, 5, 36, 78, 68, 23, -7, 19, 39, -28, -60, -15, -22, 9, 11, 48, 52, -4, -5, -3, -57, 39, -17, 20, 64, -99, 9, -8, -12, -1, -19, 37, 48, -22, -1, 53, -41, -21, -14, -52, 15, -70, 29, 51, -5, 60, -20, 10, -24, -22, -49, -18, 3, -9, 24, 107, -32, -1, -34, -24, -29, -32, 41, -53, 80, -55, -21, 65, -8, 26, -39, 23, -40, 62, -7, -2, 3, 2, -9, 64, -41, -32, -11, -51, 2, -47, 62, -30, -1, 57, -29, -35, 0, -56, -5, -44, 11, -10, -24, 48, -60, 13, 23, -83, 71, -8, -25, 82, -76, 64, -19, -10, -12, -57, -8, 65, -28, 51, 13, 17, -10, -38, 2, 24, -47, 19, 0, 72, -42, 43, -12, 1, 13, -39, 10, -37, 1, 35, 9, 8, -39, 10, -31, 6, 45, 13, 25, 4, 2, -22, -49, 3, 39, -10, -14, 5, -3, -37, -27, -64, 17, 30, -43, 1, 57, 8, -8, -26, 5, 57, -13, 28, -82, 43, 0, -14, 26, -21, 21, -45, 3, -7, -39, 48, -63, -8, 54, -52, 77, -18, 46, -68, 37, 25, -82, 69, -81, 43, 51, -6, -23, 17, 15, -86, 21, 25, -91, 61, -58, 39, -5, -42, -38, 78, -37, 56, 15, -46, 8, 4, 9, 28, 39, 27, 20, 28, -49, 57, -37, -86, 32, -5, 57, -10, 12, 27, -24, -45, -8, -3, -46, 35, -72, 3, -35, 66, -1, -29, 75, -90, 53, 17, -95, 22, -20, 70, -55, -13, 18, 53, 51, -9, -13, 7, -56, -51, -30, -37, 62, 1, 30, 34, 0, -32, 37, -12, -29, 32, -116, 23, -4, -40, -12, 88, 27, 0, 47, -53, 38, -4, -34, 3, -20, -17, 24, -105, 44, 20, -74, 24, -58, 99, -44, 59, -46, 46, 18, -70, 49, -72, 71, -47, 12, 110, -25, -24, -37, 5, 18, 11, 35, 0, -3, 49, -48, -39, -39, 92, -28, 42, 37, 3, 54, -25, -8, -12, 31, 17, 8, 11, -61, 6, -17, -64, 81, -70, 1, -9, -1, 19, -35, -29, 69, -38, 68, 15, 27, 100, -41, -37, -15, -20, 21, 12, 15, -41, -7, -38, 0, 29, -73, -14, -37, -44, -24, -10, 10, 66, -40, -4, 9, -18, -2, -106, 53, -9, 12, 3, -21, -18, 62, 36, -15, 3, 14, -17, -6, -75, 79, 30, 4, 7, 31, -38, 38, -105, 79, -29, -9, 103, -82, 12, -72, -23, 4, -49, 66, 10, -7, -8, -9, 70, 17, 18, 36, 2, 14, -3, -39, 65, -13, 13, -23, 29, -38, -64, 17, 24, -9, -20, 47, -91, -19, -21, 21, -4, -23, 14, 3, 34, 3, -35, 20, -6, -29, -52, -11, 29, -70, 24, 20, 63, -23, -13, 48, -6, -3, -41, -58, 34, 34, 20, 24, -10, 47, -25, -56, -38, -5, 60, -41, -34, 72, -27, 38, -21, -19, 1, -17, -2, -86, 43, 29, -6, -37, -31, -32, -14, 38, -23, 2, -42, 68, 7, 8, -48, 19, -24, -56, 73, -29, 32, 14, -48, 9, -34, 23, -32, -3, -48, 39, 5, -85, 52, -52, 39, -34, -4, 7, -24, -11, 47, 35, -12, 35, -4, -6, 28, -31, 57, -38, -13, 46, 2, -10, 18, 37, -11, 28, -49, -44, -3, -63, 7, -23, 10, 79, 7, 0, -14, 4, 39, -12, 0, 71, 1, 41, 55, -48, 7, 8, -4, -51, -69, -43, -34, -14, -22, 4, 34, 70, -4, 73, -71, 34, -3, -23, 82, -20, 34, -65, 13, -31, -38, -11, 17, 18, 14, 20, 0, 2, -83, 43, -14, 36, -1, 35, 0, -38, 71, -36, -7, 69, -64, 43, -64, 10, -34, -39, 4, -48, 75, -7, -37, -11, 95, 0, 40, 18, -15, 13, -31, -40, 42, -53, 32, 20, 8, 2, 8, -45, 14, -2, -85, -5, 91, -4, 52, -4, -8, 30, 35, -9, -68, 39, 20, -4, -7, -41, 56, -57, -15, 20, -87, 43, -13, 31, 11, 31, -22, 83, -54, -20, -28, 22, -38, -49, 34, -61, 94, -75, 69, -36, -17, 65, -58, 103, -27, -29, -11, -27, -51, 29, -14, 47, 11, -42, 9, 42, -35, 32, 0, 9, 23, 10, 63, -45, -9, -69, 2, 25, -7, -5, 6, -15, 45, -49, 2, 83, -13, 40, -36, -2, 0, -2, 28, -51, 11, -31, -3, 40, 12, -36, -11, -11, -52, 0, -4, -14, 52, -69, 54, -20, -35, -63, -43, -37, -19, 8, -4, 18, 40, -17, 21, 46, 7, -5, 17, 5, 100, 0, 10, -24, 47, -21, -17, 23, -24, 26, 35, -19, 19, -14, 28, 14, -43, 51, -31, 19, -31, 45, -39, 27, -104, -9, -29, -13, -5, 41, 39, 41, -14, -17, 18, 5, -100, 53, 12, -55, 48, -26, 8, -30, -72, 66, -36, 39, 35, 45, 25, -18, 17, 18, -12, 10, -27, 6, 65, -19, 14, -13, -15, -13, 78, -49, -21, 62, -34, 53, -60, -26, 69, -73, 39, 0, -41, 99, -23, 66, -23, -22, -23, -13, 51, -44, 19, -13, 9, -4, 29, 38, -37, 47, -59, 28, -2, -56, 7, 6, -28, 12, 20, -44, 53, 0, 25, -37, -9, 24, -40, 24, -14, -10, 13, -72, 24, 12, -13, -88, 12, -21, -13, -6, 44, 47, 32, 54, 8, -6, -6, -3, -45, -6, 7, -75, 13, 19, -29, 64, -49, 45, -36, 0, 52, -3, -62, 36, -21, -77, 61, -60, 38, 23, 6, 13, 8, 70, -78, 20, -4, -2, 6, -17, 36, -17, -12, 48, 43, 38, 56, 54, -30, 32, -13, -20, -35, -82, -7, 7, -37, 29, 0, 6, 70, -110, 43, -12, -6, 25, -88, -44, 25, 15, -47, 1, 15, 92, -61, 32, -3, 43, 3, -89, 34, -27, 23, -22, 63, -66, 2, -65, -2, 31, -39, -12, 27, 8, -24, 27, 22, -27, 49, -23, -20, -30, 35, 54, -11, 17, 61, -31, -5, -76, -3, -27, -37, 30, 8, -27, 9, 45, -8, 53, 13, 27, 40, 39, 17, 23, 55, 19, -59, 29, -30, -35, -79, 26, -26, 11, -22, -20, 2, -95, 37, -12, -11, 54, 39, 20, 58, -65, 61, -48, -7, -22, 15, 43, -42, 78, -66, 8, -4, -21, 61, -71, -4, 10, 0, -2, -95, 12, -21, -40, 45, -13, -8, -24, 2, -36, 55, -21, 6, 49, 70, 1, -4, -14, 21, -39, 10, 0, -36, 49, -103, 17, 24, -66, 61, -41, 31, -26, -38, 12, 24, -11, -26, -6, 77, -9, 39, 42, -19, 19, 8, -3, 58, 2, 42, -31, -57, -25, -26, 10, 49, 52, 24, -40, 12, -74, -3, 25, -38, 76, -2, -1, 27, -92, 53, 19, -60, -5, -51, 22, 19, -63, 21, 12, -4, 82, -21, 20, -8, 36, 9, -98, 18, 9, -18, -22, 13, -79, 25, -8, -38, 46, -8, 0, 57, -62, 42, 12, -104, 57, -38, 43, -15, 40, 9, -58, 36, -27, 26, -87, -2, -19, 6, -12, 36, 1, -79, 45, 5, -18, -7, 22, -13, 6, -28, 20, 25, -74, 27, -25, 5, -41, -15, 82, -52, -18, -5, -4, 71, 9, -17, -31, -1, -3, 4, -37, -10, 22, 37, 17, 20, 40, -58, -5, -52, 17, -20, -3, 25, -5, 30, -28, -46, 105, -24, 46, 3, 39, 19, 4, -64, 0, -48, -55, 15, 28, 19, 31, 12, 64, -73, 57, -3, -18, 79, -71, -9, -31, -24, 4, -44, 105, -46, 53, -73, 0, -21, -7, 8, 2, 1, -29, 35, 11, -61, -3, -9, -40, -28, -1, -41, 8, -51, 15, -13, 27, -78, -8, -10, -54, 99, -28, 26, -36, -59, 11, -8, -20, 47, 62, 73, -29, -34, 38, 6, 0, -70, -13, 38, 41, -3, 28, 46, -15, 22, -55, -26, 14, -28, 56, -37, -6, 5, -28, -12, 12, -6, -55, -8, -58, -49, 36, -54, 83, -7, -5, 51, 36, -4, -46, 9, -42, -6, -87, 1, -14, -29, 96, 9, -4, -15, 5, -4, -13, -85, 38, 66, -15, 44, 14, 64, -68, -42, 0, 24, -48, 36, 19, 2, 66, -38, 39, 6, -85, 8, -25, 12, 7, 71, -6, 11, 20, 36, -13, -36, -26, -2, 53, -32, 0, 68, -24, 23, -64, -7, -5, 37, -26, -20, -58, 25, -2, 21, 3, -14, 53, -90, -5, -32, -35, 38, -1, -23, 59, 0, 28, -36, -29, 0, -1, 5, 6, 40, 55, 9, -10, -35, 64, -10, 32, -38, 11, -2, -42, 9, -41, 2, -22, 89, -44, -12, 65, 15, 0, 36, -73, 28, 23, -60, 73, -55, 5, -23, -28, 41, -30, -34, 2, -18, -11, 3, 36, 42, 78, -4, 17, -21, 21, -25, -38, -7, 34, -3, -39, 30, 17, -64, 24, 32, 10, -9, -31, 11, 0, -24, -45, 31, -40, 85, -3, 34, -29, 90, -30, 32, -98, -21, -10, 4, -5, -18, 0, 36, -36, 18, -27, 65, -58, 44, -99, 65, 24, -51, 7, -4, 35, -29, 9, 56, -71, 53, -65, 27, -55, 11, -53, 17, 59, 15, 15, 12, 12, 38, -57, -25, 36, 3, -2, -44, 18, -14, 5, 28, -8, -37, 19, 20, -41, 12, -89, 55, -2, 40, -7, -6, 34, -43, 46, -23, 24, 62, -23, 14, -2, 24, -24, 26, 62, 0, -21, -17, -32, -8, -54, 39, -26, 79, 0, 29, 7, -90, 57, -14, -13, 13, 10, 13, -32, 63, 25, 46, 0, 10, -36, -40, -14, 37, -18, 70, 3, 34, -63, -24, -54, -19, -6, 5, 44, -18, -8, 46, -21, 29, -10, 91, -72, 17, -35, 10, -66, 2, 86, -10, -8, 4, -43, 74, -14, -11, 52, -66, 65, -17, -55, 79, -39, 112, -14, 6, 81, -70, -7, -35, -10, -10, -27, 40, -74, 52, 0, 2, 21, 0, 78, -57, 35, -4, 8, -77, 9, -79, 46, 4, 20, 35, -8, 9, 3, -41, -1, -7, -75, 65, 11, 22, -52, 12, -27, -45, -34, -26, 3, 44, -6, -42, 56, -1, 2, 27, -20, -45, -54, -9, 5, 19, 10, -12, 55, -5, 14, 59, -19, -2, -12, -60, -48, 12, -21, 53, -5, -34, 42, 13, -106, 65, -18, -78, 15, -23, 83, -52, -15, 15, 25, 42, 27, 14, -9, 44, -1, -94, 5, -54, 14, -11, -88, 24, -51, -2, -28, 7, 64, -12, -4, 38, -11, -8, 32, -105, 58, 1, 27, -6, 5, 62, -73, -13, -32, 48, -36, -2, 15, 55, 17, 45, -53, 18, -14, -60, 13, -35, -56, 94, -11, 38, 0, 5, 77, -40, 15, -34, -61, -26, 40, 9, 24, -30, -25, 53, 32, -19, -17, 8, 6, 7, 30, -48, 21, 23, -47, 65, -85, 41, -23, -37, -6, 44, -47, 55, -66, 10, 55, -28, -11, 3, 23, 7, -61, 10, -5, -35, 24, 79, -25, -5, -19, -9, 11, -2, -4, 15, 70, -10, -12, -4, -21, 12, -43, -49, 49, -21, 56, 20, 0, -14, 74, -20, -44, 1, -71, 42, -25, 1, 7, 15, 11, -47, 109, -45, 25, -25, -23, 61, -55, 19, 4, -75, 66, -10, -44, 37, 40, 48, 29, -5, -21, 19, -19, 25, -34, -37, 51, 48, -55, -60, 23, -18, 66, -63, -38, 2, -20, 21, -22, -17, 14, 43, -45, 44, -76, 18, -60, 36, -13, 60, -41, -14, 69, -56, 56, -37, 13, 56, 6, 29, -37, 17, -5, -47, 19, -21, 26, -55, 29, 75, -72, -5, 23, -55, 45, -45, 19, 31, 7, 15, 47, 6, 19, -27, 51, 2, -75, 37, -7, -5, 21, -57, 4, -56, -32, -74, 25, -41, 71, 9, 22, 59, -75, 38, -15, -27, -15, -81, 22, -7, 41, 10, -31, 20, -1, -42, -8, -18, 91, 0, 19, -22, -17, 28, -10, -3, -15, 39, 25, -3, -42, 32, -8, -93, 42, -7, -17, 57, 25, -44, 27, -41, -4, 77, -36, -6, 66, -64, 51, -57, -13, 119, -22, 27, -46, 34, 5, -68, 23, -49, 54, 53, 15, 7, 10, 6, -65, 34, -29, 46, -2, -35, 55, 5, -6, 62, -79, 10, -29, -8, -82, -3, 58, -38, 8, -35, 41, -21, -6, 61, -2, 61, 37, 3, 63, -39, -6, 4, -1, -39, 25, -71, -10, 8, 23, -19, 21, -1, 40, -22, 18, 41, 52, -51, 5, 37, 26, -30, -7, 87, 9, -45, -5, -52, -27, 0, 14, -24, 8, -26, -42, 35, 0, -9, 42, -68, -45, -20, 6, -26, 24, 58, 56, 37, -41, 12, 18, -41, 24, -3, -49, -8, -6, 23, -11, 6, 31, 22, -64, 54, 13, -61, 25, -4, 35, -35, -31, 26, 9, -12, -22, 5, -25, 12, -43, -62, 0, -4, -5, 7, -9, -31, 27, 20, 4, 51, 11, -6, 42, 20, -21, 93, -23, -32, -22, -15, 7, -28, -40, 13, 75, -42, -6, 58, -30, -1, -74, 55, 51, -30, 5, 23, 9, 26, -94, 12, -59, 2, 12, 36, 49, 10, 12, 52, 12, 34, -82, -4, -35, -4, -12, -3, 37, -21, 17, 47, -62, 5, -82, 3, 24, -56, 39, 20, 21, 21, 11, 44, -42, 21, 5, -58, 81, -44, 66, -42, -14, 22, -12, -52, 64, -39, 69, -13, -18, 71, -65, 52, -62, 62, -18, 0, 54, -56, 44, -58, -46, 40, 10, -72, -21, 54, 0, 28, 37, 54, -70, 82, -93, 51, -19, -54, 109, -66, 14, 26, -77, 47, -61, -25, 25, -32, 12, 7, 5, 63, 28, 8, 5, 55, 80, -38, 0, -7, -34, -40, -7, 2, -37, 17, -3, 42, -41, 0, 34, -11, -32, 8, 38, -20, 23, -18, 82, -63, -7, 22, -36, 10, 9, -73, 30, -5, -26, -10, 28, -55, 64, -18, -8, -4, 48, -25, 6, 31, 52, -93, 3, -5, -34, 32, -45, 17, 51, -51, 38, -19, 44, -86, 44, -13, 4, -21, -43, -17, 2, -61, 61, -18, -24, 82, -32, 15, 60, -74, 17, -36, 21, -29, 30, -27, 72, -17, 69, -29, -2, -29, 26, 15, -57, -31, 38, -14, -4, -19, -31, 26, -39, 37, -54, 79, -45, -56, 37, -7, -8, -42, 61, -19, 36, 41, -72, 48, -41, 40, -42, -66, 38, -34, 14, 1, 45, 6, -4, 57, -89, 54, 1, -112, 0, 18, -18, 21, -30, -3, 62, 25, 10, 1, 40, -18, -72, 43, 5, -23, -62, 15, 39, -21, 24, 60, -4, 55, -62, 26, -38, 2, -79, 31, -52, -19, 7, -46, 89, -41, -2, 8, 23, 69, -53, 19, -24, -7, 47, -29, 58, -75, 30, -73, 41, -11, 27, 13, 27, -31, -46, -9, -11, -35, 44, 63, 64, 37, -6, -22, 10, 27, -31, 36, -73, 24, -17, 18, -40, -22, 43, 22, -23, 42, -4, -21, 2, 34, -65, 63, -57, 24, 0, -5, 23, -4, -43, -53, 2, 29, -48, 39, 23, 23, 14, -3, -43, -23, -40, -45, 5, -17, 53, 28, 86, -7, 6, 11, 8, -13, -13, -20, 26, 1, -86, 11, 1, -53, -34, 96, -26, 25, 24, -26, 0, 40, -14, -14, 11, 10, 0, 0, 44, 1, -32, -37, -9, -13, -25, 9, -13, 26, -15, 25, 13, 43, -4, 24, -7, -17, -26, -41, -20, 18, 57, -7, 56, -28, 8, 23, -58, 27, -41, 25, 18, -31, -37, 62, 5, -86, 36, -37, 22, -34, -2, -45, 42, -25, 39, -76, 24, -25, -64, 15, 52, -23, -11, 1, 8, -31, -83, 19, 28, -11, -59, -19, 0, -6, -4, 61, 64, 4, -32, 46, 9, 13, -24, -32, 11, -25, -51, 2, -89, 34, -5, 4, 8, 1, 42, -20, 82, -56, 7, 108, -53, 41, -76, -39, 25, 23, -23, 28, -30, 90, 8, -41, 42, -65, 49, -21, 5, 45, -36, 53, -25, 88, -20, -27, 27, -32, -12, 64, -76, -2, 38, 14, 3, -7, 23, -1, -27, 76, -55, 64, 10, -81, -4, -68, 27, -6, 9, 65, -18, 47, 31, -32, 107, -75, -7, -51, -49, -9, -57, 18, 5, 24, 68, -9, 14, -3, 19, 27, -11, 98, -64, -25, 9, -35, -30, -15, -30, 72, -25, 29, 17, -36, 72, -7, -27, 9, 22, -64, -5, 37, 21, -27, -57, -27, -71, 34, -7, 57, 14, 7, 44, -29, -56, -22, 31, 20, -28, -15, 74, 19, -68, -23, 4, 37, -34, 57, -20, -8, 54, -29, 5, -62, -1, 34, -47, 65, -41, 18, 34, -75, -7, 8, -28, -9, -48, 42, -40, -28, 108, -27, -11, 6, 3, 83, -30, -1, 22, -68, 57, -41, 49, 51, -2, 64, -55, 63, -15, -69, 87, -9, -13, -26, -80, 24, 53, 6, 23, 9, -19, -40, -75, -22, 56, -26, 37, -41, 44, 10, -74, 79, -38, 77, -18, -22, 49, -60, 42, -56, 47, 7, -34, 26, -25, 42, -19, -19, 34, -28, -24, 5, -27, -8, 25, -14, -32, 22, -28, -4, -8, 18, 11, -5, 76, -32, -32, 44, -4, 25, -71, 11, -40, 13, 10, -22, 19, -3, 43, -22, -7, 51, -58, 44, 40, -63, 23, -55, -69, -40, -2, 54, 11, 39, -18, 22, -17, -54, -76, 1, 4, -26, 23, 61, 17, 21, -10, 28, -15, -47, 4, 9, -30, 25, -74, 89, 11, 10, 52, -72, 17, -6, 4, 30, -4, -32, 11, 18, -35, -48, 75, -36, 12, -30, 57, 24, 10, -17, 27, -85, 15, 0, 8, 48, 31, -28, 19, 71, -27, -11, -32, 63, -54, 6, 102, -14, 64, -71, 46, 8, -39, 18, -47, -21, 11, -19, -69, 53, -30, 35, -76, 52, 35, 40, -54, 30, 5, -53, -10, -100, 43, -8, -37, 0, 21, 39, -38, 83, -39, 48, -28, -57, 10, 13, -63, 6, 7, -12, -19, 25, 15, 40, -34, -11, 62, -38, 95, -6, -3, -13, -13, -2, -46, -39, 35, -29, 5, 0, 59, -8, 23, -11, 52, 24, -53, 44, -64, -2, -6, -59, 2, 17, -26, 43, -47, 52, -65, 68, -5, 12, -10, 34, -65, 8, 36, -36, 27, -1, -23, 34, -59, 7, -11, 53, 7, 81, -14, 14, -12, -27, 78, -19, 10, -60, -5, 19, 24, 14, 7, -15, 41, -57, 70, -62, 74, -7, -42, 17, -9, -37, -8, -22, 25, -44, -44, 61, -24, 46, 0, -15, -17, -1, 49, -41, 36, -80, 20, 9, -18, 34, 5, -10, 86, -73, 80, -58, 69, -36, -76, 38, 32, -35, -19, 63, -26, -36, -57, 30, 12, 2, 3, 61, 0, -42, 25, -47, 20, -58, 17, 0, -12, 32, 32, 19, -60, 9, 5, -26, 21, -17, 83, -1, 17, -43, 13, -12, -30, 26, -72, 1, -11, -61, 104, -14, 55, -28, 19, 29, 18, 7, -10, -8, -26, -95, -14, 32, -36, 31, -6, 56, 26, -61, 2, -18, -24, 38, 20, -17, -6, -9, -29, -61, 49, -30, 52, -44, -5, 63, -10, 23, -11, 32, -60, 82, -18, 18, 19, -40, 21, -49, -31, 63, -21, 14, -75, 3, -22, -24, 59, -8, 15, 43, -21, 47, -78, 15, 4, 61, -69, 25, -5, -23, 10, -75, 60, -5, -23, 21, -8, 78, -38, 3, 18, 29, -22, -57, 18, 9, 5, 13, 5, 54, -38, 12, 36, -79, 82, -88, 47, -14, 0, 18, -39, -2, 24, 63, -49, -2, -34, -9, 3, 26, 6, -41, -1, -53, -76, -1, 23, 10, 5, 1, -13, 83, -43, 28, 42, 53, 42, -29, -17, -13, -37, 38, -76, 12, 59, -37, 70, -31, 31, 92, -80, 13, -29, 0, 2, -70, 41, -30, -13, 42, -31, 44, -52, 25, 47, -49, 0, -19, 0, 55, -38, 23, -56, -31, -42, 15, -42, 12, 93, 10, 39, 46, -7, 60, -91, 26, 0, -31, 5, -6, 88, -51, -38, 20, 36, -44, 27, 25, -34, 73, -72, 11, 44, -34, 29, 59, -47, -72, 45, 34, -14, -17, -46, 43, -25, 31, 19, -20, 63, -53, 38, -21, -58, 1, 27, -22, 12, 15, 5, 68, 27, 14, -7, -8, 0, -6, 25, -102, -30, -7, 0, 9, -9, 10, 48, 5, -14, -4, -35, 19, 12, -29, 72, -83, -17, 0, -3, -80, 64, -55, 44, 19, -12, 64, -20, 56, 59, -14, 43, -59, 55, 39, -42, -42, 18, 1, -61, -36, -9, -42, 94, -26, 31, 51, -7, 32, -59, 14, -20, 28, -71, -47, 5, 11, -34, 14, -19, 97, -21, -14, 38, -49, 65, -27, -8, 2, 34, 47, -49, -34, 62, -13, -31, 14, 0, 76, -22, 4, 52, -80, -22, 15, -1, 45, 35, 54, -53, 41, -63, -15, -56, 25, 30, -22, 37, 10, -21, 59, -49, -34, -6, -8, 49, -12, 24, -28, 62, -11, 9, -1, -45, -35, -29, -29, 39, -100, -1, 12, -87, 62, -37, 75, -2, 27, 40, 8, 15, -27, 64, -43, -63, 26, 35, -55, 12, 42, -45, 2, 9, 11, 25, 63, 85, 23, -27, 35, -47, -49, 1, -56, 78, -2, 24, -23, 17, 2, -90, 52, -51, 8, -19, 61, 13, 18, 10, -54, 73, -11, 51, 52, -10, -25, 35, 0, -2, 7, 75, -49, 57, 42, -72, 10, -85, 32, 22, 11, 22, -57, -5, -24, 2, -15, -7, -75, 63, -28, 17, 13, 14, 86, -29, 55, 28, -70, -10, -52, 17, -19, 35, -14, 31, 17, 58, 4, -40, 4, 8, -8, 21, -18, 20, -28, 63, -11, -12, 31, -31, -24, 22, -4, -36, 89, -35, -22, -15, 9, -4, -26, 51, -4, -53, -8, -12, 3, -9, 96, -30, -26, -5, -87, 20, 32, 38, 9, 11, 15, -21, 21, -93, 53, 2, -71, 15, -45, -9, 75, -23, -30, 12, -26, -24, -56, 39, -4, 5, -24, 11, -43, 24, -100, 1, 64, -17, 54, -9, 6, 81, -4, -5, -18, -15, -8, 28, -49, 62, 4, 9, 14, -9, 56, -37, -85, 3, 23, -37, 31, -17, 6, 65, -29, 58, 8, -19, -27, -3, -24, 26, -27, 17, 41, -4, 88, -45, 3, -10, 21, -27, -9, 79, -1, -42, -17, -5, -43, 4, -5, 0, 70, -34, 6, -18, -23, -72, 4, 31, -34, 6, 14, -36, 32, 22, -35, 72, -51, 43, 29, -75, 0, -5, -44, -5, -2, 83, -4, -24, 11, -6, -28, 21, -37, 37, 47, -22, 27, -68, -39, -31, 3, 32, -30, -38, 22, -28, -15, 38, -13, 47, 56, -20, 63, -107, 73, 27, -62, 46, -83, 32, 17, -22, -51, -22, -47, 27, 14, -18, 64, -25, -14, -21, -74, 53, -44, 47, 38, 29, -17, -28, 106, -2, 49, 13, -2, 32, -24, 31, -55, 29, -38, -13, -45, 51, -36, 42, -7, -5, 83, -47, 27, 10, -15, -1, -31, -54, -21, -48, 63, 12, -21, 27, 28, -23, 45, -85, 20, -82, 12, 34, -83, 59, -26, -8, 29, -79, 6, -74, 64, -6, 20, 21, 3, -21, 28, -30, 28, 57, 22, 58, -26, 9, -6, -9, -1, 34, -57, -10, 2, -13, 59, -22, 26, 52, -78, -11, -32, 14, 47, -28, -14, -53, 28, 27, -5, 32, 37, -5, -58, 8, -24, 55, 8, 27, -11, 27, -32, -59, 0, 8, -89, 18, -4, 40, -8, 7, 39, 57, -25, 3, -7, 21, -88, 64, 21, -29, 27, -40, 18, -60, 11, -10, 15, 63, 31, 40, -59, 10, 2, 54, -43, -10, 38, -56, 17, 26, -23, -7, 22, -46, 98, -52, 77, 2, -58, 23, -47, 13, -55, 9, 29, 23, -51, -1, -6, -34, 43, -8, 19, -3, 43, -8, -9, 20, -13, -22, 21, -20, 74, 24, -13, 19, 24, 0, -79, 1, -8, 20, -46, -37, 21, 6, 0, 14, 49, -38, 55, -44, 22, -69, 20, 51, -44, -6, 0, 10, -28, 19, 43, -32, 26, 47, -72, 14, -24, -60, -5, -26, 49, -22, -37, 47, -29, -102, 8, -35, 9, 1, 15, 6, 17, 26, 24, 21, 60, 21, -32, 38, -46, 37, -36, -4, -71, 28, -4, 28, -55, -17, -13, -4, 9, 8, 36, -27, 60, -110, 29, 77, -11, 25, -1, -5, 12, -6, -54, 63, -82, 30, 26, -54, 26, 49, -99, 79, -95, 23, -31, -75, 73, -10, 26, 13, 17, 4, 47, -41, -8, 78, -69, 31, -64, -18, 32, -21, 55, 30, 86, 6, 14, 72, -55, 2, -14, -53, -56, -19, -54, 65, -11, -1, 10, 69, 55, 15, 11, 14, -24, -9, -20, -56, 5, -81, 17, 3, -92, 49, -54, 69, -13, -81, 13, -12, -21, -28, 28, -7, 12, 31, 15, 4, 17, -9, -27, 18, -74, 54, 48, -3, 27, -27, 59, -29, -59, 39, -97, 44, 18, -17, 6, -43, 89, 8, 7, -35, 32, 7, -41, 89, -66, 52, -8, -15, -29, -49, 38, 23, 5, 56, -9, 20, -24, -30, -26, -40, -35, -68, -1, -31, -13, 30, -11, 10, 51, 41, 37, 38, 12, 23, -12, 35, -36, -55, 44, -23, -28, -38, 8, -19, 28, -27, 15, 78, 6, 37, 2, 0, 75, 10, 11, 15, -11, -20, -13, -14, -87, -1, 40, -36, 14, 25, 35, -6, -2, 52, -78, 48, 8, -31, 29, -27, 64, -58, -22, 20, -8, 4, -36, 55, -37, -17, 20, 15, 3, -73, 0, 2, -13, -8, -37, -24, 58, -57, 32, -11, 24, 15, -11, 45, 44, 12, -29, 25, -54, 0, -42, -12, -13, -64, 20, 26, -52, 9, 51, -57, -13, -26, -38, 30, 14, 77, -7, -9, 29, -26, 3, -30, 7, 39, -37, -40, 19, -75, 1, -2, 46, 57, 21, 17, -29, -58, -21, 0, 39, 14, 8, -28, 47, 26, -22, -3, -37, -12, -21, 5, 20, -38, 21, 8, 10, 19, 24, 31, -56, 39, -47, 12, -14, 22, 2, -32, 5, -4, -21, -66, -38, -30, -12, 13, -28, -63, 47, -23, 12, 5, 23, -26, 87, -38, 20, 35, -57, 72, -10, 47, 29, 0, 46, -68, 10, -19, 21, 36, -10, -27, -8, -12, 49, -34, 55, -32, 8, -26, -70, 46, 3, 17, 2, 39, 15, -82, 9, -10, -72, 26, -39, 15, 28, 41, 28, 30, -37, -45, 10, 1, 0, -43, 9, 36, -11, 48, -6, -7, -41, -21, -31, -24, -79, 25, -4, 27, 30, -3, 73, -110, 35, -19, -29, -1, -18, 4, 0, -9, 46, -73, -11, 28, 38, -58, -7, 15, -37, 41, -73, 27, -86, 12, 40, 3, 26, -5, 19, -2, 10, -10, -52, 37, -57, 41, -49, 61, -9, 8, 46, 6, 36, 35, -26, 12, 19, -19, 32, 1, 35, -10, 49, -45, -22, 31, 55, -5, 7, 34, 12, 39, -56, -26, 38, -45, -4, -1, -18, 93, 5, 30, -45, 26, -74, 8, 35, -27, 45, -34, 38, -52, -57, 69, -35, -20, 46, -2, 73, -36, 6, 0, -20, 0, -23, 14, 54, -28, 32, -25, -10, 5, -10, -39, 82, -2, 27, 38, -28, 68, -27, -31, 55, -31, -52, -40, -8, 7, -69, 47, -35, 29, -11, -29, 82, -55, 60, 29, 65, 12, -12, 70, -70, -7, -38, -30, 39, -20, -22, 29, -14, 38, -44, -22, 3, -86, -31, 81, -35, 75, 9, -26, 48, -106, 36, 15, 15, 64, -1, -31, -4, 32, -52, 60, -9, 13, 47, -29, -2, 25, -15, -19, 10, -10, -24, -34, 20, -53, -7, 11, -31, 10, 22, 15, -46, 66, -36, 10, 73, -82, -15, -6, -46, 7, -34, -1, 58, -32, -7, 7, 46, -74, 74, -38, -6, -66, -11, 2, -41, 57, -6, 28, 25, 53, -5, 13, -1, -10, 52, -30, -43, 27, -45, 2, 59, -91, -18, 12, -47, 5, -23, 21, 30, 14, 38, 62, 12, 31, -61, -48, -2, 15, -37, 19, 18, 52, 15, 15, -8, -14, 11, -31, 28, -62, 30, 6, 26, 17, 0, 42, -69, 48, 47, 15, 19, -46, 10, -51, -19, -45, -27, 27, -44, 46, -66, 98, 4, 7, 77, -70, 25, 19, -22, -38, -3, -85, 15, 8, -4, -74, 45, -7, 1, 34, -5, 59, -96, 44, -32, 9, -97, 0, 45, 30, -3, 8, 20, 32, -58, 31, -41, 23, -46, -40, -1, -68, 23, 7, -19, 53, -56, -26, -5, 2, 19, -31, 2, 27, 36, 51, 3, -30, 13, -80, 20, 4, -32, 14, 24, 46, -39, 41, -5, 49, 42, -35, -23, 14, -25, -72, 21, 12, 22, -12, 15, 34, -82, 37, -46, -39, 38, -34, 110, 19, 7, 9, 21, 1, -47, -40, -15, -22, 20, -56, -32, 55, 61, -76, -8, 25, -32, 35, -59, 29, -46, -12, -27, 6, 40, -44, -23, 86, -45, 111, 4, 5, 25, -58, -9, -18, 11, -39, 64, -45, -24, 27, -77, 20, 20, -19, 37, -57, 53, -6, -51, 71, 0, -34, -35, -7, 66, -38, 66, -27, 25, -10, -49, 61, -9, 19, 68, -2, 28, 68, -126, 59, -21, -23, 41, -87, 18, 11, -18, 21, 36, -48, 23, -45, -9, -46, -38, 41, 39, 23, -7, 14, -26, 8, -10, 22, 11, 6, 0, -38, 40, -27, 49, -26, -4, 8, 0, -27, -28, 25, 22, -38, 37, -94, 8, -58, -40, 8, -49, 117, -9, 48, -11, -14, -47, -20, -13, -68, 12, -80, 47, 13, 19, 14, 64, -31, 47, -38, -65, -23, -18, 25, 0, -20, 12, -29, -58, 10, -91, 109, -38, 31, 23, 0, -19, -19, 53, -90, 53, -112, 76, 37, 21, 22, -4, 63, -70, -8, -5, -11, 42, -48, -31, 61, -34, 24, 9, -35, 17, 14, 31, -8, 20, 113, -31, -6, 30, -35, -15, 1, -72, 35, -24, 44, -41, -44, -13, -2, -74, 52, -43, -12, 47, -12, 41, 18, -3, -59, 34, -43, 44, 9, 63, -8, 2, 70, -49, -32, 2, 5, -4, -45, 59, 4, 4, 88, 30, -75, 20, -103, -6, 13, -55, 26, -14, 30, 47, 9, 47, 14, 25, 27, -35, 1, 26, -17, -12, 116, -55, 0, 20, -24, 18, -17, -8, -45, 51, -1, -36, 49, 20, -42, 18, -85, -30, 22, -22, 27, 8, 29, 5, 21, -81, 22, 23, -15, 57, -37, 38, -55, 57, 34, -8, -69, 22, 6, 30, -29, -21, 4, -55, 7, -36, 62, 3, 18, -14, 10, 13, 12, 18, -37, 27, 51, -41, 95, -5, -52, 45, -40, -7, 18, -47, 6, -36, 12, 15, -18, -64, 22, 0, 69, -27, 5, -22, -24, -9, 15, -12, -52, 5, 29, 3, -71, -52, 22, 37, 6, -13, -41, 26, 23, 20, -6, 7, -10, 40, -25, 20, 41, -41, 21, -7, -1, -79, -28, 35, -38, 71, -30, -5, 8, 9, 2, -45, 45, -88, 51, -22, 37, -8, 56, 2, 39, -58, 38, -41, 14, -40, -49, 43, 19, -36, -70, 47, -17, 1, 15, -39, 42, -40, -14, 30, -6, 45, -22, -4, -29, -4, -32, 0, -24, 20, -14, 48, -23, -4, 24, -86, -12, -43, -42, -35, 49, 47, 47, -1, -25, 28, -48, 81, -22, 32, -31, -9, 6, -49, 39, -68, 71, 23, -26, 63, -34, 48, 0, -53, 13, -20, -28, -14, -10, 6, -29, 0, 7, 17, -81, 21, 45, -48, 36, -39, 10, 58, 0, -3, 24, -6, 6, -73, -72, -47, -10, 19, 6, -6, 6, 48, -22, 0, -17, 45, -43, -7, 15, 0, -5, 38, -38, 32, 48, -64, 31, -4, -10, -9, 12, 22, -89, 28, -44, -8, 37, -37, -7, 44, -10, -12, 27, 8, 34, -80, 4, 4, -57, -15, 72, -59, 78, -27, -26, 18, -44, 3, -4, -40, 78, -17, -20, 58, -11, 42, -36, -21, 6, -78, -3, -18, -54, 61, -13, 42, 0, -6, -64, -1, 1, -51, -15, 24, 45, 39, 31, 21, -3, -41, -57, -38, -14, 56, 28, -3, -36, -4, -39, 4, -23, 7, -42, 21, 12, 0, 13, -4, 57, 27, 39, 55, 42, -72, -13, -60, -14, 3, -10, 3, -18, -7, -7, 93, -26, -17, -11, -5, 22, -54, 6, 79, -23, 49, -51, -56, -13, 39, 22, 56, 34, -19, 20, -40, -48, -9, -38, 28, -42, 35, -48, 97, -30, 12, 20, 4, -9, 70, -34, -35, 62, -61, 6, -44, -4, 28, -5, 98, -18, -10, 25, -34, 2, -36, 34, -108, -15, -13, 36, 8, 26, 17, -24, 35, -46, -13, -59, 1, 24, -34, 0, 54, -21, 98, -8, -35, 22, -47, -11, 31, -6, 20, -2, 76, -40, 103, -51, 17, -55, -85, -6, 29, -17, 58, 2, 15, -17, -23, 18, 28, -20, -22, 52, -56, -44, -34, -20, 57, 1, 32, -3, -17, 58, -11, 62, 38, 23, 0, 0, -26, -36, 7, -31, -4, 42, -9, -26, 78, -57, 70, -57, 4, -71, 17, -7, -58, 31, -49, 102, -47, 19, 38, -19, 53, -21, -38, 59, -18, 38, -23, -56, 7, 43, -45, 8, 58, -11, 70, -26, 38, -10, -45, 5, -48, 31, -9, -2, 0, 64, -110, 19, -38, -1, 82, -42, -7, -9, 34, -14, -66, 63, -56, 75, -75, 8, 40, -13, 36, 2, 18, 8, -72, -7, 17, -18, -44, 74, -68, 28, 4, 20, -34, 77, -36, -12, 41, -20, -83, 31, -39, -43, 11, 51, 26, 0, 26, -2, 2, -7, -10, 76, -18, -23, 29, 42, -51, -43, 35, -8, 1, -51, 66, -30, -59, -10, -26, 45, -4, 26, 59, -4, -15, 51, -45, -56, -2, 54, -30, 29, -10, -10, 57, 10, 45, 41, -51, -4, 8, 14, -5, -44, 11, 22, 18, -62, 20, -65, 18, 43, -51, 0, 0, 78, -40, 3, 29, -57, 58, -25, 34, 35, 0, 43, -5, 36, -128, 6, 6, 1, 41, 17, -31, 26, 23, 12, -9, -15, 42, 3, -8, 0, 42, -8, -20, -58, -27, -25, 12, 22, -38, -18, 56, 25, -28, -9, -1, -25, 17, 8, -53, -3, 45, -1, -10, 12, -43, 45, -19, 54, 31, 58, 26, -13, 21, -32, 17, -49, 10, -65, 36, -35, -13, -8, -36, 79, 5, -1, 9, 74, -98, 25, -40, 14, -13, 25, -49, 36, 91, -14, 58, -56, 44, -25, -29, 15, -18, -36, -7, -23, 35, -2, 10, 4, 65, -12, -8, 19, -2, -8, -37, 56, -28, 2, 23, -72, 27, 41, -9, -22, 18, 46, -61, 87, -25, 60, -74, -1, -35, -63, 32, 5, -36, 31, 6, 15, 0, -49, 56, 31, 20, -28, 26, -37, 15, -32, -18, 82, 25, 54, -73, 5, -87, -45, 20, -10, 65, 22, -21, 41, 27, -13, 17, -5, 17, -47, -35, -64, -12, 56, -24, -21, -15, 69, -43, 23, 0, 8, 22, -6, -9, 49, 13, -35, 27, -59, 51, 72, -32, -49, 38, -49, -3, 0, -5, 95, -49, 30, -62, -43, -19, 0, -18, 58, -57, -11, 20, 13, 9, 17, 28, -66, 22, -14, 60, -12, -1, -23, 46, 14, -40, 13, 38, -20, 104, -11, -13, 64, -28, 29, 31, -52, 1, -55, 2, -30, -26, -31, 60, 59, 12, -14, 0, 18, 39, -62, -9, 52, -76, 10, 26, -20, -11, 41, 29, 46, 2, 20, -11, 13, 44, -43, 32, -24, 34, 42, 6, -25, -13, -3, -48, 78, -4, 21, 17, -35, 40, -35, -2, -1, 32, -13, 25, 27, 32, 24, 85, -47, 48, -21, -39, -36, -55, -40, -44, -35, 47, -58, -4, 72, 24, 18, 41, -27, 103, -45, -15, -49, -41, 29, -17, -11, 36, -47, 114, -65, 10, 6, -49, 40, -7, 29, 68, 66, 22, 11, 41, -74, -19, -24, -45, 7, -98, 13, 28, 3, 20, 56, 17, 21, 22, -39, 3, -46, 7, -76, 103, -44, 66, -21, 6, -8, -39, 2, 24, -82, -13, 39, -64, 23, 45, -12, 48, 4, 25, 1, -43, 13, 26, 14, -9, 44, -1, 43, -14, -21, 24, -42, -31, 90, -21, 32, 17, 60, -4, -85, 34, -49, 52, -66, 8, 36, 9, 8, -34, 73, -58, 30, 8, 31, -63, 29, -49, 52, -23, -5, -6, 18, -41, -11, 18, 9, -3, -62, 18, 60, -37, 44, -62, 51, 8, -11, 94, -54, -8, -10, -17, -31, -43, 29, 12, 64, -9, -3, 47, -14, -76, -23, -42, 36, -37, 2, 60, -43, 73, 24, -3, 65, -72, 1, 10, -2, -49, 3, 0, 20, -92, 19, 59, -17, 61, -73, 46, -44, -14, 20, -81, 35, -60, 62, -52, 4, 113, -49, 22, -12, -35, 0, -41, -9, 17, -38, 42, -26, -12, 4, -34, 4, -6, -48, 57, 19, -30, 37, 14, -54, 61, -6, 19, -39, 15, -13, -22, 17, -64, 68, 21, -40, 63, -9, -46, 51, -18, -24, -53, -38, -3, -36, 11, 39, -22, 86, -13, -30, -30, -42, -32, -1, -49, 19, 27, -6, 65, 23, -56, -13, -32, 6, 53, 9, 8, -38, 6, -20, -1, 55, -47, 3, -9, 58, -45, -22, 28, -12, 52, -89, -15, 64, 21, -17, 22, 23, 0, 55, -51, 40, -64, 36, -3, 36, 0, 1, 23, -113, -21, 3, -5, 1, 13, -1, 76, -11, 28, -32, -10, 46, -27, 13, 40, -19, 62, -83, 39, -34, 42, 21, 63, 40, -22, 18, 4, 6, -115, 73, 35, -60, 46, -80, -2, 27, 30, 0, -7, -3, -14, -23, -6, -117, 52, -32, 23, 37, -22, 55, -85, 20, 29, -26, -40, 21, 52, -4, -57, 1, -11, 48, -4, -2, 39, 39, -100, -21, -20, 9, 5, 7, 58, 31, -12, 37, -27, -15, -21, -2, 11, 7, -81, 26, -32, 6, -14, 19, -14, 7, 34, -46, -35, 0, -17, -66, -14, 29, 15, 62, 43, 22, 2, 1, -32, -53, -17, -60, 31, 39, -49, 34, -27, 9, 28, -57, 38, -90, 17, -4, -4, 83, 73, 58, 12, 18, -19, -25, -43, 0, -12, -43, -4, 8, -46, -22, -25, -58, 66, -44, 74, 26, -11, 3, -90, 51, 6, 4, -8, -3, 59, -78, 98, -61, 19, 48, -43, 27, -45, 77, -5, -35, 0, -69, 29, -18, -11, -13, 10, 102, -38, 12, 27, -47, 22, -52, 25, -12, 31, 59, 11, -8, 100, -96, 58, -11, -39, 61, -52, 72, -47, 78, -54, -4, 1, -42, 32, -7, -46, 41, 32, -9, 9, 0, -3, -6, -57, -13, 2, 19, -12, 53, -38, 47, -51, 24, 43, -19, 54, 0, 80, 45, -36, -4, -9, -61, -48, 7, 2, 58, -29, 64, -34, 48, 20, -111, -27, -43, 30, -43, 81, 27, 9, 55, -75, 46, 2, -38, -36, 25, -8, -93, 30, -13, 44, -12, -10, 38, 32, -38, 34, -94, 47, -9, -36, 87, 20, 27, -45, 12, -28, -13, -13, -55, 96, -46, 12, -54, 61, -14, -13, -44, 32, 10, -56, 83, -41, 14, 107, -34, 42, -58, -11, -8, -23, -6, 43, -5, 4, 0, -82, 40, 38, -28, -19, -11, 18, -59, 52, 20, -17, 6, 37, 57, -36, -26, 59, 3, 15, -38, 11, 53, -47, 25, -107, 90, 10, -38, 71, -29, 98, -13, -91, 42, -47, -19, 5, -63, 92, -74, 37, 48, 5, 51, -29, 1, -48, -48, -3, -42, 82, 6, -46, 3, -27, -35, 62, -30, -18, 43, -61, 46, -37, -35, 41, -69, 49, -32, -54, 31, -19, -7, 35, -51, 45, -30, 35, -30, 69, -48, -25, -17, -36, -11, -70, 61, -35, -10, 43, 18, -54, 1, 35, -26, 65, -18, -7, 31, -21, 25, 9, 13, -32, 41, -3, -7, 19, 35, 48, -28, 8, 63, -43, -5, -80, 30, 31, -42, 53, -2, 11, 1, -51, 0, 0, -14, -30, -4, -23, 47, 0, -28, 29, -45, 11, -30, 3, 14, 24, -49, 13, 36, 49, 29, -6, 30, -35, 42, -7, -49, 40, -94, 51, 69, -37, 22, 30, -44, -29, -54, -25, -71, 59, -29, 11, -3, 23, -30, -7, 18, 19, 10, 8, 38, -10, -36, 49, 7, -36, 14, 21, -14, 0, -12, -34, 95, -38, 4, 60, -57, 63, -8, -30, 77, -76, 2, -48, -6, 13, -6, 10, 47, 18, -89, -6, -63, -20, -13, -25, 89, 7, -17, -25, 43, -20, -56, 31, 2, 51, -94, 12, 42, 18, -18, -30, 56, 29, -61, -15, 10, -9, 21, -56, -9, -17, 38, -3, 3, -29, 6, -7, -9, 1, 23, -49, 28, -3, 43, -21, 11, 32, -68, 56, -5, -8, 20, 76, 57, -7, -5, 20, -63, -7, -54, -12, 5, -4, 5, 11, 63, 0, 53, 30, 11, 21, -51, 95, -34, 8, 22, 20, 44, -29, 25, -22, 47, -49, -56, 44, 18, -6, 35, 30, -48, 35, -5, -36, -30, -46, 15, 26, -29, 12, 25, -68, 22, -64, -23, -2, 26, 23, 20, 32, 1, 51, -19, -75, 38, 47, -5, -57, -3, 5, 0, 44, -12, 1, -1, -10, -2, -11, -31, 9, 20, -82, 74, -75, 41, -58, 58, -4, -34, 24, -2, 80, -14, -21, -3, 24, -40, 61, 6, 43, 29, -26, 2, -43, -24, -1, -24, 45, -44, 51, -41, 48, -76, -11, -75, -7, 9, -59, 54, -47, 38, 18, 19, 12, 0, 59, -91, 12, -4, -18, -9, -20, -3, 5, 9, -53, 5, -32, -1, -9, -21, 56, 18, -17, 19, -23, 113, -48, 37, -42, 63, 5, -53, 66, -49, 3, -12, -7, -12, 20, 28, 36, 30, -39, 35, -43, 80, -30, -25, 39, 30, 65, -41, 10, -5, -11, -54, -41, 55, 2, 32, -63, -14, -35, -24, 31, -24, 40, -46, -24, 83, -46, 43, 44, 18, 89, -14, -27, 60, -38, 6, -87, 57, -21, -42, 38, -39, 63, 2, -5, 27, 7, 55, -2, 20, 49, -82, 7, -10, 13, -71, 56, 38, -36, 45, -24, 40, -13, -20, 23, -56, -8, 24, -97, 54, -22, -53, 110, -4, -35, 7, 30, 0, -58, 6, -54, -55, -42, 46, -34, 34, 13, 44, 0, -36, -31, 90, 3, 30, 6, -13, 45, -58, 19, -34, 18, 38, -61, -24, 12, -24, 35, 11, 29, 36, 2, 3, 60, -3, -21, -10, 15, -37, 1, 30, -6, 10, 11, -13, 77, -43, 28, -21, 8, 18, 13, -80, 25, -26, -23, 46, -48, 15, -49, -9, 11, -65, 64, 9, 40, 19, 18, 4, 12, -14, -2, -4, 44, -57, 5, -18, -24, -34, -22, -9, -8, -41, 62, -38, -39, 38, 18, -40, -17, 17, 37, 11, -11, -48, 14, -7, 1, 54, 46, 29, 57, 6, -79, -10, -36, 13, -49, -42, 30, -9, 19, -38, -4, 1, 17, 3, 42, 1, 55, -14, 5, -3, -11, 4, -9, -8, 93, 0, 2, -32, -11, 32, -65, 82, -49, -18, 76, -34, 69, -15, 54, 19, -58, 71, -52, 56, -21, -25, -1, 15, 4, -11, 40, -97, 38, -8, -4, 34, -42, 9, -44, -32, -1, -34, 0, -56, 78, -24, -15, 78, -94, -11, 46, -28, 0, 63, -8, 69, -44, -24, -9, -21, 17, -53, 8, 108, -56, -34, 15, -41, 76, 23, 42, 10, 7, -39, -83, 4, 40, -34, 37, -3, 12, 13, -61, 72, 17, -45, 54, -44, -23, -7, -46, 55, -72, 27, 10, -65, 46, 18, 41, 21, 23, 45, -55, 45, -28, -14, -58, 63, 22, -53, 21, -45, -8, -64, -19, 15, -23, 20, 31, 18, 26, 47, -54, 39, -14, -32, 24, -9, -13, -15, 9, -82, -2, -13, 43, 7, -34, 19, 23, 10, -22, -9, -47, -31, -20, -7, -9, -17, 62, -6, -5, -29, 0, -38, 49, -93, 72, 34, -83, 46, -59, -14, 15, -42, 54, 24, -29, -43, 17, -35, -27, 21, -30, 86, -41, 34, 4, -6, 78, -59, -6, 0, -68, 4, -17, -22, 70, 24, 10, -54, 9, 15, 14, -53, 14, 30, -11, -82, -12, 11, 10, 5, 60, 24, -22, 74, -29, -4, -28, -3, -43, 19, -36, 30, -28, -14, 18, 36, -37, 18, -18, 73, -69, 32, -79, 12, 24, -27, -14, 47, -86, 94, -3, 36, -7, -6, -27, -36, -15, -64, 93, -17, 48, 13, 15, 51, -60, 43, 26, -7, -52, 21, -27, 6, -35, -48, 6, 12, 2, -2, 31, 75, -56, 7, -62, -14, 8, -57, 36, 23, 4, 61, 2, -29, -25, -6, 8, -65, -17, 79, -43, 63, -44, -17, 28, -66, 127, 1, 37, -42, 12, -23, -53, 19, -41, 25, 18, -55, -6, 48, -12, -3, 1, 42, -14, 0, 47, 53, 35, 38, -7, 14, -15, -17, 20, -37, -61, 42, 30, -51, 58, -37, 70, -1, -20, 75, -14, 23, -60, -21, 8, 1, -13, -19, 12, -13, -11, 11, 21, -1, 52, 85, -4, -19, -21, 15, 7, -36, -25, -41, 64, 7, 9, 0, -8, 54, -43, 1, 9, 23, -8, -35, -5, 15, -43, -11, 54, -56, 85, -56, 37, -15, -18, 90, -3, -55, -10, 35, 8, -22, -41, 20, 6, -21, -11, 39, -17, 91, 5, 4, 35, -77, -17, -19, 59, -46, 1, 9, 38, 27, 8, 39, 24, -37, -26, -51, -49, 19, 25, -48, 64, -92, 32, 8, -72, 114, -30, -20, 52, -71, 44, -17, 2, -6, 52, 25, 7, 81, 0, -60, -18, -17, 18, -5, 12, 0, 8, 20, -4, -31, 42, -3, -82, 12, -31, 37, -72, 18, -44, 6, 8, -35, 32, -39, 66, -2, 57, 51, -13, -45, -3, 10, 13, 53, -19, 3, -36, -39, 30, -68, 37, 0, -9, 83, -20, 53, 31, -19, 97, -23, 23, -70, -38, 1, 30, -12, 34, -35, 38, -11, -9, -60, 6, -60, -51, -22, -13, 13, 5, 7, 62, -7, 51, -34, -14, 21, -28, 6, 32, -9, 19, -52, 45, 31, 17, 5, 7, -15, -25, -1, 46, -42, -10, 5, -38, -30, 46, 24, 7, -25, 68, -58, -7, 0, 21, 9, -59, 42, -9, -60, -34, 0, 18, -38, -37, 19, -65, 40, -63, 34, -8, -56, 64, 19, -23, -7, 20, 41, -47, 34, 53, -30, 18, 24, 48, -82, 5, 0, -48, 52, -3, -37, 39, -41, 35, -44, 8, 55, -2, 29, 1, 0, 3, -48, 22, -77, 74, -22, -18, 9, 22, -5, -65, -3, -22, -23, -1, 0, 0, 13, 34, 45, 9, -8, 5, -21, 13, 11, -30, 77, 0, 9, 14, -22, -46, -46, -46, 14, -2, -60, 7, 11, 18, -58, 27, -15, -48, 45, 20, -29, 38, 7, 3, 43, -31, -4, -10, -22, 6, -6, -1, -6, 34, -25, 27, 38, 54, -42, 9, -45, -17, -22, -57, 39, -64, 45, -30, 65, -37, -12, 22, 40, -35, 74, -20, 5, 19, 8, 2, -42, 55, -48, 28, -43, -4, -56, -24, -57, -2, 36, 2, 27, 11, -1, 46, -42, 61, -9, 26, -24, -6, 4, 17, -17, 35, -65, 0, -51, -42, -18, -37, -41, 103, -7, 44, 54, -58, 78, -31, 5, 57, -85, 7, -63, -35, -1, -1, -28, -44, 70, -46, 11, 23, 5, 65, -61, 5, 39, 3, -10, -11, 42, 0, 64, 2, -32, -6, -55, 32, 36, 25, 52, 0, -28, -29, -76, 3, 17, -40, 44, -95, 41, 18, -30, 49, -24, 72, 17, 2, 18, -46, 19, -31, -45, 39, -19, 2, -54, 99, -52, 4, 53, -5, 42, 34, -13, -10, 21, -86, 51, -42, 1, 47, -7, 58, -5, -5, 45, -47, 47, -7, -45, 10, -37, -1, 39, -62, 74, 12, -53, 28, -58, -14, -89, -6, -4, -15, 29, -39, 37, -5, 52, 21, 3, -12, -1, 51, -19, -21, 69, -62, -22, -18, -46, -34, 96, 4, 13, 17, 6, -18, -25, -48, 10, -12, 48, -22, 19, -47, 0, -48, -51, 55, 23, 41, -37, 46, -62, 20, 24, -62, 79, -120, 30, -13, 23, -6, 0, -38, 0, 17, -53, 23, 60, 2, -4, 58, -22, 36, 27, -39, 6, -2, -70, 9, -13, -5, 53, -55, 32, 11, 14, -47, -2, 54, -70, 0, 11, -82, 59, -17, -38, 43, 10, 7, 46, 30, -44, 95, -68, 20, -10, -22, 21, -63, 15, -87, 36, -1, -27, 44, -37, -40, 18, -32, 10, 37, 10, 75, -34, 8, 4, -74, 83, -1, 0, 14, 28, -42, 22, 17, 56, -22, -2, 3, -51, -5, 41, -59, 31, -20, -45, 18, -15, 85, 18, 8, -57, 35, 3, 39, -7, 36, -32, 29, -42, -85, 59, -68, 102, -4, -8, 59, -72, 26, 8, -51, 31, -15, -55, -40, -20, 61, -24, 61, 0, -28, 81, -72, 85, -13, -17, 49, -53, -77, 46, 9, 7, 46, 17, 18, -13, 30, -17, -64, 66, 23, 11, 9, -62, -12, -46, -2, 11, 9, 36, 0, 76, -83, 40, -22, -77, 27, 35, -7, 1, 1, -2, -2, 7, -69, 20, 30, -30, 6, 48, -75, 6, -30, 74, 0, 37, -12, 77, -49, 52, -35, -57, 36, 14, -12, -13, 48, -37, -47, -43, -52, 10, -36, 66, 52, 38, 10, -21, 37, 11, -35, -11, 4, -13, -80, -21, 12, 37, -59, -18, -15, -12, 27, 25, 58, 49, -37, 14, -23, -7, 11, -92, 17, 36, -26, -17, 45, 86, -8, -42, 22, -13, 12, -58, 12, 21, -66, 44, -35, -60, 13, -32, 66, 1, 73, -13, -20, 7, -30, -15, 12, -87, 44, 0, -13, -69, 35, 19, -72, 55, -34, 13, 8, 27, -15, 110, -58, -34, 9, 0, 35, -63, 7, 10, 47, 20, -29, 8, -23, -38, -53, 2, -62, -5, 0, -98, 43, -47, 42, 17, 44, 78, -55, -29, 11, 19, -13, -30, 12, 29, 56, 9, -19, 0, -44, -12, -9, -44, -2, 57, 0, -46, 28, -54, 25, -21, -92, 65, 13, -9, 13, -31, 121, -5, -13, 53, -100, 5, 15, -83, 71, -30, 11, 127, -24, -29, 18, -26, -19, -26, -14, 85, -79, -29, 24, -5, 1, -27, 51, 22, -11, -70, 19, 7, -44, -10, 63, -46, 57, 42, -1, 32, -11, 29, -114, 38, 0, -4, 14, -61, 26, -18, -35, 115, -23, 34, -51, 14, -7, -60, -2, 54, 27, 23, 12, -18, 27, 15, -102, 71, 17, -63, 41, -71, -8, -18, -59, 46, 22, -8, 25, 5, -8, -43, -65, -21, -21, -11, 12, -25, 24, 87, 2, 30, 25, -63, -19, -53, -22, 64, 10, -10, -2, 42, -15, 41, -68, 17, -30, -51, -61, 53, -12, 11, 59, -51, 49, -18, 45, -71, 4, 35, -18, 13, -61, 75, 0, -29, -20, 25, -1, -18, -70, -11, 15, 25, -40, -44, -17, -17, 5, 20, 44, 28, 27, 23, 48, -99, 18, -11, 22, -45, -32, 68, -23, -1, -52, 56, -5, -53, 49, -48, 3, -32, -30, 78, -60, 58, -37, -7, -12, -60, 29, 17, -35, -28, -2, 38, -53, 38, 14, 19, 17, 13, 72, 24, 51, 5, -8, 26, -26, -76, -2, 52, -11, 22, 22, 30, 77, -29, -8, 3, -40, 35, -6, -14, -21, -13, 15, 21, -34, 30, -28, 32, -2, -94, 53, -51, 14, 5, -42, 34, 39, 4, 27, 40, 41, -106, 61, -7, -18, 22, -77, 14, -27, 25, -91, 39, -31, 45, 43, 23, 9, -15, 1, -40, 12, -11, -24, 73, -70, 1, -42, -21, 28, -40, -3, 41, -42, 6, 27, 15, -14, -3, 9, 4, 2, 5, -68, -4, 38, -4, 9, 0, 55, -40, 28, 44, -85, 25, -39, 56, -4, -29, 48, -52, 41, -24, -86, 41, 38, -41, -30, 41, 8, 0, -6, 1, 56, -86, -12, 91, -5, 48, -26, -20, 29, 0, 6, -2, -9, -7, -2, 41, -21, -27, -40, -26, -45, 63, -31, 17, -23, 98, -11, 39, -35, 8, 23, -43, -55, -2, -24, 21, 13, 31, 1, -11, 43, -14, 72, -65, 26, 32, -69, -6, -62, 23, 32, 23, -25, -12, -25, -53, 28, 28, 71, 8, -36, -13, -46, -13, -17, 0, 62, 0, 41, 38, -7, 71, -82, 26, -36, 5, -8, -26, 52, 34, 2, 38, -76, -7, -45, 26, -15, 34, 31, 52, 22, -18, 40, -81, 57, -27, -24, -32, 21, 88, -36, 31, 15, -5, 10, -70, 11, -39, -41, -2, 12, 47, -29, -24, 27, 29, -24, -30, -21, -2, 27, -28, -2, 70, -62, -22, -58, -17, 29, -28, 27, -77, 3, -6, -29, 52, 24, 55, 36, -19, 75, -31, 36, -38, 7, -64, -61, -35, -32, 45, 7, 4, 28, 31, -80, 2, -36, -64, 44, -49, 20, 0, -37, 32, -29, 2, 37, -30, 46, 22, -13, 47, 0, -9, 35, 24, -27, 70, -18, 17, -23, -24, 9, 40, -25, 40, 4, -81, 21, -1, -8, 28, -10, 57, 27, -24, -73, 6, 11, 19, -38, -58, 45, 1, -83, 81, -25, 82, -18, -59, 14, -25, -28, 60, 27, 12, 41, -8, -20, 17, -40, -5, -71, 22, 15, -66, 68, 29, -70, 8, -7, 32, 6, 0, -28, 55, -14, -23, 76, -51, 76, -57, -9, -10, 2, -21, -80, 58, 14, -48, 13, -10, 60, -86, -12, 82, -7, 47, -24, -19, 1, 48, -37, 54, 18, -25, 25, 3, -58, 86, -69, -23, -55, -40, 55, -58, 94, 28, 5, 90, -87, 81, 0, -71, 13, -81, -13, -38, 17, 37, 2, 22, 32, -30, 12, -56, 60, -69, 73, 7, 86, 47, -30, 17, -56, -31, -21, -22, -36, -40, 52, 18, -11, -39, 58, 3, -14, 69, -5, -15, 20, -56, 7, 0, -73, 0, -9, 35, 44, 2, -32, 2, -62, -15, 26, 4, 45, -34, 53, -23, -63, -35, -41, -21, 59, -10, 12, 44, 37, -36, -22, 2, -15, -24, -80, 34, 23, -28, 29, -5, 18, -45, 21, -3, -82, -1, -38, 14, -30, -27, 17, 24, -26, 49, -20, 18, 40, -47, -19, 25, -42, 27, -93, 2, 44, -19, 22, -3, -40, 19, 60, -28, 5, 27, 11, 10, -2, -11, -35, 65, 13, -44, 5, -40, -1, -64, 70, -77, -18, 80, -59, 34, -2, 58, 1, 9, -35, 55, -2, 57, 23, -2, -13, -34, -13, 42, -24, 24, -32, -3, -45, -45, 3, -52, 70, -37, -28, 22, -25, -3, -18, 25, 47, 32, 71, 11, 53, -36, -8, -7, -87, -5, -1, -29, 39, 0, -59, 99, -38, -23, 77, -75, 68, 6, -53, 97, -36, 10, 56, -70, 13, 40, -85, 12, -51, 3, 41, -42, 34, 29, 18, -30, 15, -22, -71, 58, 4, 6, -9, 59, 43, -80, -44, -8, -25, 28, -57, -25, 59, -70, 57, -21, 51, 68, 41, 10, 7, -41, -3, -14, -1, -35, 40, 28, -6, -85, 19, 0, -42, 25, 37, 2, 23, -83, 25, 31, -4, 21, 23, 7, -31, -15, -30, 7, -32, -11, 73, 9, -27, -13, -25, -17, -5, -48, 68, -15, 20, 86, -11, 54, 10, -53, 19, -32, 45, -43, 40, 30, -79, 17, -40, -39, 37, 7, 34, 58, -24, 32, 6, -37, 76, -68, 60, -14, -28, 5, -25, 0, 5, -102, 60, -46, 64, -12, -6, 48, -49, 51, -22, -52, -14, 8, -17, 26, -2, 32, -38, 9, -9, -14, 88, -41, -5, 51, -82, 59, 2, -57, 45, 0, -28, 11, -13, -21, 5, -55, -32, 26, -40, 11, 38, 65, 0, 40, -53, 53, 20, -75, 6, 41, -7, 64, -19, -43, -23, 20, 28, 21, 31, 6, 35, -21, -14, -62, -10, 60, -17, 17, 14, -47, 11, -23, 15, 23, -41, 41, -22, 19, -42, -25, 38, 31, -2, -34, 45, -53, 86, -52, -44, 52, 12, 13, 24, 10, 90, -57, -17, 32, -35, -39, -44, 1, 35, 0, 36, 24, -58, 34, 31, 14, 23, 40, 44, -57, -8, -45, 35, -41, 71, -4, 34, 14, -66, 0, 1, -6, -31, 8, 13, -6, -14, -61, 58, -72, 74, -7, -29, 22, -48, -7, 54, 11, 64, 23, -30, 64, -32, 5, 5, -44, 1, 27, -29, 127, -18, -19, 18, 4, 21, -46, -22, -72, -6, -1, -6, -5, -28, 53, -26, -21, 28, 5, -52, -26, -2, -23, 3, -40, 66, 25, -10, 12, -6, -9, 77, -10, 20, 30, -91, 22, -32, 8, -7, 39, -7, -21, 83, -24, 61, -28, 41, -8, -11, -71, 0, 48, -66, 18, -5, -25, 52, -15, 34, 14, -2, 3, -39, 51, -12, 5, 48, -35, -36, 15, -2, -73, 25, 9, 38, 38, 11, 87, -77, 4, -43, -68, -5, 2, 10, 26, -28, 54, 39, 7, 34, -26, -2, -13, -70, 37, -28, -7, 74, -17, 2, -10, -1, -54, -55, 64, 21, 10, 5, -27, -10, -52, -6, -77, 20, 38, 14, 36, 21, -58, 65, 4, -46, 62, -7, 68, 6, -38, 30, -20, -29, -40, 31, -5, 22, 28, 45, -65, 52, -64, -18, -7, -17, 14, -24, -9, 52, -9, -12, -37, -15, 42, -24, 38, 26, -14, 49, -12, -2, -1, -1, 8, 20, -30, 71, 2, -7, -42, 0, -24, -44, 63, -5, 56, 11, 70, -41, 2, -42, -20, -26, -9, -69, -6, 29, 11, -46, -3, 38, -13, 4, -6, 78, -48, 18, -25, 30, -94, 86, 15, -5, -1, -12, 12, 45, -34, -5, 43, 57, -39, -48, -3, -46, 47, -9, -6, 6, 63, -56, 0, -11, 62, -13, -35, 29, -44, 37, -32, -3, 74, -4, -2, 76, -20, 54, -30, -45, 5, -47, 77, -25, 23, 31, -60, -5, -43, 47, -42, 47, 77, -45, 34, -41, 56, -7, -6, 80, -124, 23, 4, 25, -12, -37, -5, -32, -22, -40, 46, 15, -14, -2, 6, -49, 10, -70, 28, -44, 60, -51, -12, 48, -81, 78, -22, 88, -10, -12, 17, -68, 32, 62, -31, 21, -56, 39, 17, -44, -30, -10, 35, -7, 7, 35, -1, -11, -38, 9, 36, -63, 10, 0, 10, 1, -38, 19, -30, 21, -46, 51, 71, -54, -34, -1, 4, -15, 38, 11, -3, 82, -66, -23, -15, -34, 36, -1, -6, 37, -27, -47, 23, -15, -9, 11, -1, -20, 2, -2, 2, 51, -5, -21, 39, -39, -29, 11, -38, -28, 72, -57, -18, 47, -15, 6, -1, -42, 10, 39, -41, 10, 34, -38, 111, -24, 29, -58, 5, -46, 0, -47, 20, 9, -8, 31, 10, -100, 79, -37, 48, -31, -28, 55, -86, 99, -3, 76, 7, 14, 39, -75, -19, 12, -26, -49, -51, 62, 17, -28, -45, 23, 31, -46, 100, -56, 13, 32, -51, 22, -93, 19, 31, -83, 57, -45, 19, 56, -7, -2, -4, 42, -34, 56, -40, 3, 5, -10, -56, -61, -26, -43, 32, -29, 83, 9, 9, -11, -30, 3, 39, -61, 35, 0, -35, 21, -8, -11, 24, -53, 74, -28, 28, -18, -6, -58, -41, -39, 12, -14, 21, -22, -14, 96, 19, 38, -8, -28, 40, -40, -15, -13, -51, 70, -36, 20, 65, 77, 61, 12, -19, -27, -53, -5, -60, 53, -28, 23, 68, 12, 19, -19, -4, 40, -35, -8, 20, 32, -37, -17, 18, -4, -3, -3, -6, -14, -26, 21, 57, -3, 9, -23, 65, 2, -44, 44, -14, 24, -59, 11, 72, -53, 10, 45, 2, -34, 9, 27, -72, 76, -29, 49, -7, -59, 35, 42, 4, 37, -40, 17, -4, 37, -29, -70, 45, -22, -29, 61, -23, 74, -32, -7, 14, -9, 8, 20, -76, 38, -38, -44, 31, -69, -14, 45, 39, 22, 57, -24, 22, 6, -39, -31, -7, -17, 0, 15, -39, -18, 15, -5, 68, 1, 45, -30, 38, -54, 7, -6, -40, 58, -72, -17, -42, -15, -7, -51, 21, 61, -9, -10, 30, -57, 64, -5, 22, -13, 24, -41, 73, 2, -28, -23, 29, -38, -28, -52, 106, 4, 45, 37, -41, 66, 9, -46, 48, -43, 12, -46, 1, 26, -49, 98, -92, 56, -28, -62, 24, -34, 77, -64, -14, 4, -14, -57, 0, 77, -10, 42, -14, 40, -14, -59, 0, 11, -40, -45, -24, 1, 17, 9, 35, 36, 18, 11, -25, -1, -57, 11, -68, -21, -2, -83, 116, 8, 35, 0, -5, -31, -11, -29, 25, -17, 1, 18, 39, 25, -53, 55, 13, -85, 77, -56, 15, 14, -58, 58, 11, -71, 26, -9, -91, 38, 54, -46, 9, -53, -4, 14, -26, 7, 34, 8, 39, -54, 59, 30, -40, 56, 2, -43, 43, -15, -57, -39, -31, 1, -28, -28, 49, -89, 23, -9, 1, -18, -9, 54, -10, 78, -21, 0, 23, 25, 15, -27, 49, -61, 54, 12, -22, -46, 58, -11, 30, -41, 4, -12, -45, 55, 11, -27, 38, -105, 85, 30, 12, 32, -34, 25, -22, -26, -31, 0, -82, 90, 18, 11, 40, 14, 63, 20, -34, 38, -105, -37, -62, 18, -10, -11, 45, -38, 81, -17, 11, 46, -79, 22, 15, 11, -2, -31, 26, -28, -1, 21, -80, 32, 27, -48, 27, -27, 57, 73, -35, -49, 42, -17, 4, -113, 28, 44, -34, 61, -5, 83, -14, -38, 15, -3, -49, -40, -11, -2, 34, -123, 47, -34, 13, -14, -64, 54, -2, -17, -53, 20, -76, 53, 15, 42, 45, -40, 83, -85, 17, 43, -74, 65, -100, 34, -13, -12, 0, 98, -70, -11, 10, -28, 41, -52, -32, 26, -82, 24, 14, -29, 53, -5, 29, 37, 36, 69, -37, -5, -41, -64, -56, 5, -29, 43, 41, 30, -26, -32, -23, 29, -44, 59, 59, 19, 2, -5, 48, -40, 9, -55, 52, -36, -53, 35, -5, 26, -60, 36, -30, 71, -24, 32, -26, -21, -27, -24, -18, -6, 23, -39, -7, -4, 82, -46, 34, -11, 12, -19, -60, 44, -92, 69, -19, 9, 19, -24, 60, -53, 41, -24, 17, 64, -6, 23, 44, -62, 31, 29, -54, 57, -17, -10, 11, 4, -26, 17, -43, -22, -9, -8, -55, 34, 0, -37, 81, -48, 59, 4, -35, 0, 25, -53, 61, -40, 27, 24, -94, 15, -32, 43, -10, 7, -29, -7, 30, -7, -42, 61, 20, -15, 43, -79, 26, -2, -14, 44, -25, -30, -9, -41, 20, -57, 58, 4, 36, 40, 47, -8, 12, 7, -8, -1, -48, -20, -44, 65, -78, 57, 30, 7, 68, -56, 12, -29, -56, -22, 28, 11, 36, 21, 48, -28, 80, -20, -55, 12, -51, -11, -22, 22, 40, -42, 21, 23, -57, -2, -51, -21, -48, 7, -31, 44, 46, -4, -9, 42, 24, -19, 32, -19, 54, 9, -21, 7, -31, 15, -5, -58, -10, -44, 1, -8, 59, 2, -22, 21, -83, -14, 43, -31, 20, -12, 38, 14, -5, 0, -51, 45, -1, -14, 56, 43, 23, 39, -20, -30, -3, -54, 69, 9, 13, -23, -2, -41, 3, -2, 12, 7, -11, 32, 17, -89, 43, -54, 52, -2, -34, 0, 4, -63, -26, 29, -17, 51, 1, -13, 18, -34, -8, 57, -61, 37, 32, 25, -71, -20, 42, 5, 22, 12, 6, -11, 37, -26, -40, 34, -55, -30, 1, 39, 26, 27, 20, 0, -40, 0, -31, 4, 55, 39, 27, -12, 7, -32, -35, -71, 74, 2, -30, -26, 37, 19, -44, -17, 39, -13, -34, 22, -8, -96, 36, -41, 8, -14, 86, 48, 59, 52, -56, 11, -13, -17, 1, -49, 25, 23, 6, 22, -44, 17, -27, 49, -44, 72, -13, 20, 72, -79, 1, 12, 5, -22, 4, 15, -56, 22, -32, -9, -24, -4, 29, -45, -19, 18, -10, -41, 58, 18, 22, 12, -35, -12, -12, 4, -57, 46, -22, 44, -8, 41, 43, -49, 56, -28, -5, 20, -24, 47, -56, 26, 40, -29, -41, 66, -10, -6, 82, 4, 6, -82, 2, -27, 15, -51, -23, 85, 3, -8, 10, 9, 32, -28, 29, -94, 8, 24, -76, 75, -9, 35, 6, 23, 72, 27, 25, -45, 10, -49, -51, 18, -40, 48, 73, 0, -5, -19, 13, -52, -4, -45, 38, 26, -59, 40, -29, 90, -71, -14, 0, -7, 35, 58, 14, -9, -12, -34, -8, 5, 14, 71, 4, 0, 42, -11, -13, 4, 13, -88, -4, -20, -6, -34, 63, -2, 36, -70, 8, -14, -23, -92, 45, -100, 82, -17, 56, 82, 13, -10, -14, -27, 14, -49, 44, 38, -74, 3, -4, 56, 22, -4, -13, 11, 17, 35, -31, -39, 28, -37, -38, 32, -52, 21, -81, 27, -15, -14, -7, 36, 35, -90, -37, 17, -2, -35, 42, 27, 72, 5, -1, 37, -1, -12, 35, -26, 17, 9, 21, 23, -76, 40, -25, -17, 39, -46, -59, 31, 46, -21, -18, -2, 29, 19, 19, -18, -9, 34, 11, -95, 30, -14, 20, -14, -3, 52, 24, 19 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
