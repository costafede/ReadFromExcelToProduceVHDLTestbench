-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
            -65, -124, 119, 99, -61, 1, 4, -16, -37, 71, -58, -12, 100, 51     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -6, 25, 99, -48, 127, 9, -99, -97, -87, 118, 89, -77, -40, -34, -3, 100, 75, -107, -43, 96, -114, 112, -98, 36, -41, -86, 105, -65, -68, -115, -23, -70, 24, 121, 29, -50, -83, -78, 56, -78, 11, -56, 6, -43, 97, -93, -50, -40, -116, -89, -49, 112, -71, 8, -104, 103, 34, 37, 61, -109, -77, 61, -59, 101, -61, 42, 102, 68, 42, 56, 80, -76, -38, 123, -103, 52, 42, 71, 123, -99, 88, 15, -42, -47, -64, -72, -46, -104, -42, 95, -112, 43, 39, 112, 50, -51, 84, 126, 109, -68, -108, -123, -19, -67, 23, 67, 6, -69, -33, -11, 94, -112, -113, 89, 108, 58, -109, -50, 56, -117, 54, -1, 121, 61, -92, -124, -49, 90, 63, -80, -66, 33, 14, 97, -120, -102, -23, -74, 70, 88, 50, 122, 15, -76, -44, -38, 53, -50, 10, 20, 65, -127, 9, -56, 117, 78, -25, 100, 48, -71, 106, 67, -1, 126, 76, 17, -15, 40, -49, -8, 18, 62, 9, -66, 84, 66, 63, 44, -51, -79, 63, 106, 47, -4, 9, -1, 9, -99, -15, 0, -111, 118, -45, -83, -110, 39, -23, -93, 27, -44, 118, 24, 9, -11, 90, -29, -72, -59, 55, -116, -5, -80, 122, 118, -98, -60, -89, -35, 29, -14, -60, -6, -111, -44, 97, 19, 2, -13, -106, -14, -31, -36, -60, 26, -59, -83, 105, -58, 93, 69, 57, -98, -103, 35, 67, -65, -11, 17, -41, 4, -2, 92, 37, -93, -60, -69, -94, 1, -23, 47, 22, -8, -58, -54, 58, 95, -28, 58, 96, 104, 19, -85, 89, 93, -39, 81, 115, -81, 30, -75, -15, -42, -113, 59, -105, -27, -106, -40, 117, 60, 99, -79, -60, 97, -41, -2, -15, 27, -43, 58, 117, -25, 106, -82, 20, 117, -32, -67, 77, -123, -86, -57, -38, 119, -96, 92, 3, 104, 63, -3, -27, 75, -29, -99, 27, -29, 122, 87, -24, -49, 127, 47, 59, -105, 50, 68, -93, 84, -105, 90, -65, 87, -83, -45, 97, 127, -84, -70, -111, -82, -23, 11, -102, -43, -51, -77, -99, -71, -31, -57, -20, -27, -44, 17, 31, -12, 25, 98, 116, 54, 108, 18, -92, 2, 48, 63, 7, -37, -60, 8, -57, -73, -118, -105, -102, 14, 46, 16, 85, 34, -113, 72, -118, -108, 113, 68, 61, -43, -20, 108, 37, -27, -9, 71, 72, -2, 62, 66, 56, 75, 35, -127, -23, 31, 107, 35, -10, 82, -106, 27, -77, 24, -57, 126, 16, 54, -60, 32, -69, 120, -92, -13, 37, -27, 97, 62, 85, -66, -76, -95, -64, 96, -28, -73, -122, 26, 125, 109, -12, 58, 111, 98, 75, 0, 112, -35, -102, -119, 95, 88, 89, 78, -2, -106, 20, 22, -13, 49, -42, 46, 92, 68, -12, -13, -37, 120, -20, 122, 85, -37, 44, -19, -110, 71, 103, 74, 56, -123, -79, -60, 106, -55, -78, -94, -67, -2, -62, 123, 77, -109, 64, 10, 98, -120, 71, -1, -97, -99, 126, -33, 1, 4, -53, -27, 58, -108, 10, 107, -117, 33, -119, -89, -83, -118, -53, 98, -58, 113, -27, -37, -24, -32, 70, -9, 99, -42, -120, -10, -63, 75, 93, 34, 31, -105, -8, 43, 83, -30, -6, 6, 126, -122, 39, -77, -40, 109, -125, 15, -33, -120, -109, -43, 23, -123, -38, 9, 65, -35, 11, -53, 100, -31, 102, 4, -5, 76, 120, 68, -57, -106, 111, 45, 55, -113, -8, -66, -61, -55, 98, 85, 63, 71, -76, -72, 93, 7, 20, -79, 54, 122, 39, 21, -78, -24, -15, -56, -124, -29, -9, -75, 3, 88, 82, 123, -67, -48, 103, -80, -44, 0, -54, 18, 80, -7, -62, 2, 42, 1, 90, 55, -50, -21, -29, 14, 123, -33, 21, -127, -75, -7, -106, 103, 54, -46, 53, 12, -73, -45, -39, 99, -16, 68, 72, 17, 15, -4, 121, -57, 19, 30, -78, 91, -126, -9, -14, 89, 3, 67, 88, -1, -110, 80, -61, -76, -86, -117, 89, -104, 113, -87, -94, 123, -41, -32, 21, -110, 49, 121, -8, 108, -17, -41, -92, 73, -86, 91, 82, -79, -58, -57, -75, 32, 16, 75, -30, -92, 20, 87, 30, -7, -128, 62, -71, -12, -62, 94, -24, 49, -38, 38, -109, 73, -90, -54, 39, 46, 9, 68, 65, -107, 93, -100, -48, -121, 37, -55, -60, 109, 51, 50, 115, -22, -26, -84, 36, 1, -99, -52, 115, 114, 47, 80, -48, -47, 70, -41, 48, -6, 118, 63, 52, 87, 12, -125, 19, 16, -123, -89, -17, -125, 96, 106, 108, -47, 22, -25, -91, 117, -113, -75, 34, 55, 29, 117, -47, 12, -119, -30, -13, -65, -25, 30, -120, 75, 36, 49, -123, 105, -48, -22, -37, 99, 74, -59, 82, 39, 90, 86, -49, 66, -58, -13, -30, 17, -50, -51, -55, -85, 11, 82, 50, 100, -5, -90, -88, -19, 45, -77, 81, 30, 59, 51, 115, 66, -19, -63, 70, -62, -56, -68, 113, -15, 5, 124, -79, 48, -49, 113, -76, 120, 19, 8, 106, -37, -23, 119, 83, -18, 31, 127, -9, -16, 124, -54, 23, -66, 80, -117, -110, 112, 50, 40, -4, 32, 67, 116, -55, -26, -106, 111, -38, 41, 11, -80, -7, -123, 24, 98, 43, 7, 11, 113, 101, -86, -103, -117, -7, -12, -123, -53, 53, -127, -66, 34, -35, -121, 87, -21, 75, -54, -47, -49, -52, -85, 102, 78, -37, -15, -63, 105, -108, -35, 7, 102, 21, 52, -85, -34, -77, 9, -118, -36, 81, 92, -31, 100, -38, -48, 22, -72, 107, 81, 35, -100, 125, 48, -93, 88, -71, 51, 106, 7, -37, 97, 48, 91, 61, 66, -86, -25, -100, -117, -68, -35, -3, 55, 45, 127, 100, -30, 32, -62, 46, -83, 38, -35, 35, -121, 115, 112, 77, -19, 115, 92, -72, 82, 110, -111, -100, 100, -10, 2, 26, -51, 40, 126, -11, -93, -8, 47, 23, -3, -102, -116, 28, -40, -90, 64, -33, -65, -111, -82, -110, 18, -70, 72, -40, 100, 1, -104, 107, 90, -19, -105, -28, 4, -125, 6, 92, 5, -103, 17, 52, 115, -32, -26, -63, -68, 120, -83, 102, 60, 10, 118, -66, 0, -116, -68, 70, -28, -80, -62, -11, 44, -116, -77, -87, 68, -48, 117, -80, 49, -67, 105, -84, -20, 114, -26, 97, 100, -111, 85, -86, -30, 5, 102, -100, -36, 41, -69, 96, 48, 95, -105, 126, 112, 127, -17, 113, -11, 96, 125, -41, 108, -109, 113, 16, 95, 75, -19, -101, -48, -36, 42, -100, -14, 81, 16, 97, 78, 113, 44, 88, -60, 7, 121, 98, -114, -78, 83, 56, 96, 93, 27, -35, 13, 8, -42, -2, -12, -93, -116, -4, 119, 29, 42, -113, -46, 47, 104, 19, 127, -5, 14, 119, -18, -86, -6, 104, -15, 67, 25, -46, 124, -125, -111, 121, 91, 107, 93, -56, 51, -2, -67, -101, -83, 109, 82, -88, 54, -6, -44, -29, 108, -42, -24, 26, -121, 42, 58, 17, -102, -58, -17, 38, 93, 116, 1, -73, 113, 29, -114, -27, -93, 45, -118, -11, 71, 124, 48, -118, -107, -120, 80, -54, -124, 62, 94, -104, 110, 126, 34, 118, 59, 12, 98, -5, -101, 121, -111, 84, 7, -6, 35, 43, -89, -85, -110, -67, -24, 27, -90, -123, 14, -120, 78, -104, 86, 36, 3, -84, 115, 61, 123, 69, 59, -25, 67, -120, 49, -21, -50, -42, -60, -89, -59, 120, -100, -125, 49, -45, -93, 118, -18, 106, 27, -100, -21, 25, 93, 68, -127, 111, -46, -73, -67, 62, 10, -113, -87, 71, -1, 100, -46, -37, -67, 77, 85, -30, -62, -80, 77, -18, 110, -70, 83, 68, -50, -121, -48, 38, 82, 76, -47, -19, 49, 74, 58, 117, 122, -107, 53, -37, 82, 107, -17, -78, 114, -90, 85, 22, -9, -90, -109, 42, 30, 97, 17, 113, -122, 108, -103, 90, -11, -65, 3, -1, 13, -118, 91, 124, 74, 30, -67, -126, -62, 124, 42, 40, -6, 127, -105, -111, -14, -104, 90, -65, 42, -55, -23, 74, -72, 85, 22, 18, -7, 15, 51, -109, 124, 45, 40, -50, 60, -87, -53, -37, 44, -8, 49, 83, 37, 9, -16, 77, 78, -39, -109, 117, -124, -81, 122, -101, 122, 85, -17, -118, 1, 23, -33, -8, -28, -120, -84, 56, -40, -105, 84, 60, 103, -110, 56, 13, -93, 85, 4, -73, -4, -97, 111, -45, -98, 79, 70, 57, 64, -12, -42, -97, -55, -60, -26, -113, 45, 38, 94, 84, -69, -93, -101, -76, -36, -125, -115, 4, -47, -93, -18, -128, 24, -120, -53, -75, 113, -39, -34, 65, 4, -109, -128, 50, -101, -54, 98, 20, 51, 113, 101, -23, -15, 7, -3, 89, -22, 127, -41, 53, -54, -8, -116, 84, 21, -34, 80, 76, 50, -60, 89, 31, 68, -96, 118, 110, 16, -117, -124, -109, 103, -23, 26, 48, -1, -24, -85, 115, 31, 69, 111, -112, 107, 55, 19, -39, 74, 92, -41, 9, 110, -31, -14, 40, 92, -111, 50, 89, 1, 8, -71, -46, 41, -30, -52, 104, -127, -72, -34, -28, -35, -50, 77, -30, 119, -97, 42, 40, -7, -92, 113, 104, -14, -50, 39, -113, -102, 108, 100, 9, -12, -112, -23, 10, -58, 90, 109, 116, -5, -49, -37, -124, -65, -66, 62, 96, -11, 38, 89, -114, 19, 112, -77, -108, -13, 101, -29, -27, 52, -29, 66, 87, 67, 113, 121, -126, -126, -33, 119, 103, -71, -96, 58, 97, 95, -59, 119, -1, -106, 106, 73, 111, 51, 121, -58, 74, 74, 90, -61, -9, -41, 22, 53, 72, -23, 4, 92, 10, 26, -35, 124, 4, -116, -53, -31, -53, -96, 111, 48, 122, 0, -78, 59, -19, 0, -84, 101, -70, 79, -103, 70, -47, -28, -12, -115, 91, -36, 83, 97, 75, -78, -27, 86, -63, -99, -49, 40, 126, 66, -89, 120, -33, -11, 12, 59, 113, 127, 56, 70, 59, 95, 49, -123, 32, -88, 3, -50, 54, 31, 61, -41, -4, -76, -72, -123, 98, 46, -45, -113, -41, -20, -50, -11, 19, -110, 63, 104, 85, 39, 85, -96, 21, 46, 117, -2, -107, 56, -15, -23, 6, 44, -108, -119, -19, 99, -98, 17, -69, -103, -61, 44, -96, -83, -27, -47, -78, -107, -19, -39, 93, 26, 103, 2, 13, -46, 1, 45, -33, -104, -113, -95, 87, -13, -66, 33, 85, -33, 51, 126, 76, 84, -96, -113, 60, -18, 42, -40, 30, -115, 86, 2, 37, 5, 56, 16, 31, -89, 6, -84, -4, -68, -3, 106, -110, -45, -119, 23, 0, -85, -48, -123, 32, -56, -92, -91, 105, -118, -79, -91, -37, -87, 5, -2, -38, -101, -116, 112, 91, 124, -8, 19, -128, -47, 109, -127, 102, 103, -84, 15, 7, 82, 7, -75, -50, 0, 33, -21, -128, 38, -41, -25, -45, -71, -65, -66, 9, -90, 0, 3, 34, -20, -90, 86, 103, 8, -6, 13, 75, -34, 81, 91, 22, 35, -91, 15, -41, -24, -32, -117, -122, -108, -36, 7, 110, -43, 96, 85, -5, 127, 84, -121, 102, -44, 1, -52, -52, 14, 31, -29, 47, -103, 17, -67, 70, -16, 120, 52, -52, 122, 120, -97, 102, -112, -102, 57, -5, -26, 35, 89, -69, -9, -21, -128, 94, -6, -93, 126, -5, 80, 23, 11, -85, -66, 35, 33, 42, 0, 43, -102, -21, 94, -103, 51, -77, 36, -35, -122, 99, -10, -125, -25, -69, 97, 58, -26, -4, 45, -15, -98, 58, -2, -65, 36, -127, 94, 102, 113, -42, -124, 38, -9, -54, 89, -41, 77, -14, -20, -8, -14, -117, 66, -122, -19, 71, 23, 69, -7, 105, -69, -40, 59, 60, 41, -40, -105, -56, 115, 36, 40, 91, 4, 125, 75, 81, 58, -9, 100, -70, 28, 75, 17, 61, -17, -85, 41, -120, 14, 21, 69, -51, -10, 46, 14, 20, -105, 112, 37, 56, -2, 19, 65, -10, 102, -101, -113, -5, 105, -88, -97, 24, -11, -102, 57, -18, -61, 47, -75, -1, -21, -1, -89, 60, -122, 105, -43, 35, -11, -68, -91, -76, -7, 114, -1, 80, -120, 23, -75, 3, 127, -87, 79, -61, 49, -48, 81, -51, 124, -72, 65, 0, -101, -96, 15, -51, 116, 34, -1, 70, -111, 18, 23, 50, 76, 21, -37, -10, 124, 1, 119, 14, -23, -43, 25, 7, -13, -65, 114, -90, -89, 54, -105, 81, 124, -55, -59, 102, -116, 115, -42, -60, -40, -110, 14, -36, 57, -70, 70, 76, -95, -49, -86, -87, 92, -31, -97, 82, 31, 52, -127, 72, -6, -4, 33, 69, 111, -108, -114, -19, -19, -105, -26, 15, -82, 118, -35, 17, -60, 58, 76, -125, 104, 21, -99, 32, -71, 114, -4, 13, -104, 116, -48, -9, -76, -31, -71, 21, -47, 121, -114, 72, -69, -3, 47, 86, 106, -11, 40, 9, -99, 41, -66, 103, 45, -111, -36, -76, 39, 108, 7, -31, -109, 98, -57, -67, -125, 6, 97, 53, -103, 9, 1, 86, -121, -93, 41, -76, -8, -107, 100, -47, -37, 5, -8, 50, -110, -122, 56, 34, 78, 53, 124, 55, 56, 82, 36, -1, 100, 93, -105, 84, -78, 121, 76, 3, -18, -15, -57, -125, 80, -62, -125, -43, 106, -107, 110, 70, 6, 82, 113, -15, 87, -116, -33, 105, -50, -87, -127, 46, -111, -127, -106, 32, 39, -102, -95, 100, 95, -91, -46, -104, -84, 81, 43, 104, 79, -57, -70, 20, 54, 96, 120, -114, -59, 110, 32, -16, -118, -35, 8, 41, 49, 52, -99, 79, 16, 57, -69, -31, 84, -104, 65, 76, -36, 55, -34, -28, -108, 96, 57, -89, -10, 78, -13, 103, -86, 58, -118, 1, 55, 79, -20, 103, -4, 5, 100, 9, 110, 19, 19, 29, -128, 78, -18, 72, 82, 45, -40, 44, 123, 117, -98, 44, 54, -38, 38, -33, 81, -45, -110, 122, -56, -37, -115, 112, -72, 38, 67, 43, 55, -56, -70, 2, -38, -124, 63, -24, 92, -124, -46, 39, 98, -20, 6, 26, -87, 51, 47, -50, 109, -72, -78, -31, -24, 23, -116, 38, -96, -65, 119, -83, 94, 2, -26, 87, 91, 25, -11, -59, -101, -78, -87, 102, 16, 30, 57, -42, -116, -45, 7, 52, -26, -32, -21, -96, -21, 0, -37, 10, 86, -3, 125, -116, -106, 116, 73, -4, 77, 42, -11, -13, -15, 87, 64, 7, -37, -51, -96, 63, -104, 100, -110, -5, 38, 94, -20, -79, 24, -8, 49, 100, 20, 91, -127, -77, -65, -88, 122, -91, 59, -24, -20, 87, 3, -54, 126, 42, 97, 20, -30, 107, -101, 38, 41, -52, -123, 64, 56, 116, -107, 112, 3, -128, -104, 6, -15, -31, -125, -75, -49, 37, -128, 30, 73, -57, -82, -111, -109, -32, -64, 34, -60, -19, -21, -21, 12, -121, 34, 125, -75, -69, 74, -45, 107, -109, 113, 30, -25, 33, 102, -75, -128, -46, 99, 116, -45, 30, -21, 118, -17, -76, 34, 7, 21, 29, -94, 109, 72, 67, 98, 66, -14, 37, 113, -114, 117, 1, 50, 25, 86, 46, -59, -119, 126, 1, -3, -5, -50, -96, 124, 48, -41, 101, -83, -86, -94, 39, -102, 112, 89, -36, -40, 2, -67, -87, -106, -56, 62, 41, -43, -9, -21, -21, -112, -27, -71, -49, 46, -58, 93, -14, -27, -16, -6, -90, 46, -77, -73, -98, 49, 60, 14, -107, -102, -57, 54, -98, -3, 8, 88, 49, -127, -102, -71, 48, 89, -62, -17, -10, -107, 84, 101, -51, -74, -94, 45, 121, 45, 83, -82, -73, -92, 89, -1, 1, 114, -58, 78, -126, -97, 32, -79, -122, -52, 82, 90, -65, -69, 89, -110, 29, -75, 16, 97, -53, 33, -88, 28, 23, -23, 33, -82, 103, 71, 65, 84, -23, 50, -103, 60, -19, -58, -64, -68, -103, -91, -81, 7, 29, 89, 72, -50, 36, 37, -65, -98, -26, -14, -37, -52, -93, -118, 85, -68, -17, 36, 70, -36, -54, 116, 36, -122, -128, 114, 83, 56, -19, 89, -23, -75, 124, -67, 81, -7, 28, 54, -38, -73, -11, -122, 91, -84, 124, -20, 70, -75, -124, -54, 112, 87, 65, 65, -116, -90, -28, -108, 55, -123, 82, 116, -57, 94, -54, -110, 117, -126, 32, -118, -16, -44, -100, -117, -25, -40, 34, -77, -80, -40, -22, -94, -54, 120, -98, -58, -45, 30, 117, -68, 2, 52, 117, -20, 16, 45, 112, 23, -87, 103, 105, 48, 112, 92, 44, 111, 119, 36, 58, -61, 92, 73, -30, -123, -76, 87, -89, 47, 23, -24, 31, -35, -33, 122, 89, 119, -64, 62, -1, 13, -124, -107, -90, 94, 28, 97, 29, -88, 43, 118, 95, 8, -71, 115, -82, -52, 51, 75, 67, 111, -57, -90, 14, 123, 38, 89, 30, -104, -61, 101, -45, 8, 69, -35, -112, -103, 4, -90, 30, -63, -119, 55, 59, 101, -5, -81, -109, 101, 33, 106, -100, -101, -100, 14, 72, 68, 20, 42, 27, -50, 44, 16, -2, -87, -111, -5, 85, -89, 120, 20, 126, 104, -39, 56, -90, 115, 24, 7, -32, -47, -63, -33, -97, 89, -102, 98, -117, 12, -51, 4, -6, -89, 55, -46, -53, -34, 5, 7, -70, 82, -62, 60, -3, 0, -93, 118, -92, -105, -104, -95, 49, 104, 42, -97, -44, -122, 51, -13, -93, 126, 41, -120, -55, 54, 52, 119, 61, 87, 110, -3, -91, -40, 17, 2, 55, -32, 84, 88, -92, 12, -5, 105, -69, 25, -50, -74, -5, -31, -47, 71, -44, 113, -124, 55, -113, 61, -95, 43, -42, -48, -14, 70, -97, 125, -111, 63, -60, 59, -78, 77, 98, -22, -68, 54, -21, 110, 105, -112, 97, 24, 6, -31, -41, -89, -46, -51, -12, 50, -60, 76, 103, 42, -105, -76, 126, -78, 105, 104, 86, -3, -34, 104, -9, -93, 112, -76, 68, -114, -22, -98, -58, -121, -123, -67, 49, 109, 51, 94, 68, 79, -11, -54, 78, 73, -27, 121, 97, 19, -92, -48, -67, -10, 100, 52, -15, 114, -111, -26, -18, -22, 89, 9, 17, -91, -114, -85, -38, -12, 39, -83, 10, 45, -76, 26, -20, -18, 73, -123, 78, -1, 29, 117, 124, -77, 12, -63, -82, -107, -88, -55, -27, -78, 100, -9, 105, 48, -16, 53, -11, 108, 44, -75, -93, -87, 26, -86, 78, -114, -13, -8, 11, -61, -85, -38, 116, 17, -122, 111, -116, -99, -93, 46, 28, 60, -10, -23, -19, 112, -64, -21, -49, -113, 7, 55, -70, -40, -24, 123, 24, 75, -58, 79, 89, 14, -22, 36, -127, 117, -13, -3, -118, 92, 125, 34, -19, -116, -21, -58, -68, 27, -128, -83, -33, 46, 94, -107, 109, -118, 110, 18, -113, 65, -101, -14, -38, -45, 99, 67, -122, 79, -69, 50, 11, -27, -12, 18, -84, 37, 101, -58, 10, 58, 39, -42, 103, 48, -100, -27, 45, -103, 64, 39, 100, -89, 14, 104, -6, -39, -80, 69, 124, 29, -68, 108, 123, 111, -125, 32, 48, 17, 119, -44, 14, 40, -40, 94, 108, -28, -74, -91, -77, -20, -39, -20, 115, -116, 123, 108, 92, -118, 65, 19, -86, 55, 16, 33, 53, -82, -12, 95, 57, -48, 61, 92, 95, 1, 2, -48, 62, 54, -13, 88, -59, 81, -100, -68, -4, -27, -52, 113, -106, -49, 89, 114, -44, 34, -29, -79, 113, -89, -60, -6, 121, -104, -64, -1, 86, -106, 111, -105, 78, 8, -38, -71, -119, 69, 35, -105, -40, 39, 15, 84, 16, 49, -102, 100, -81, -56, -93, -35, 10, 85, 70, 10, 47, 0, -32, 45, 54, -15, -126, 74, 18, 97, -72, 53, -31, 120, 18, 6, 52, -26, 62, -63, 118, -51, 10, -69, -85, -9, -102, 79, -17, -4, -62, 4, -112, 3, -82, 99, -65, -110, 93, -98, 100, 9, -109, 17, -111, 121, -47, 97, -83, -81, 84, 47, -82, 60, 13, 91, -117, 72, 99, -15, 26, -87, 19, -66, 56, -33, -108, 41, 92, -117, 29, -69, -81, 57, 27, -83, 76, 44, -43, 40, -77, -94, -81, -106, -47, 107, 6, 74, -48, -114, 34, -84, 52, -126, -63, 8, 48, 105, 7, -4, 48, -124, 118, 15, 126, -14, 44, 39, -99, 120, 68, 77, 27, -80, -125, 90, -17, -74, 26, -122, 87, -24, 32, -59, 16, 14, -93, 62, 29, -113, -32, 79, 88, 79, -24, -1, 72, 87, -43, -28, -86, -2, 69, -79, 62, -3, -85, 111, -124, -74, 34, -98, -23, -47, 98, 62, -128, 62, 125, -32, 73, -90, 20, 122, 120, 110, -58, -88, -24, 81, -112, 80, -81, 51, 59, 29, 86, -93, 53, -63, -57, -66, -122, 73, -9, 125, -49, -25, -7, -64, -117, -15, 96, 17, -104, -117, -81, -107, 14, -68, -10, 107, 33, -63, 44, -24, 58, -120, -45, 0, -117, -116, 110, 82, -59, 37, -33, -59, 69, -115, -16, -55, -103, -96, -4, 47, -79, -59, 39, -53, -66, 102, 99, 47, -72, 1, 59, 83, -103, -53, 60, -20, 9, -31, -26, -41, 14, 52, -90, 106, 102, 43, -50, 85, -88, -81, 27, 17, -22, -128, -77, 23, 53, -93, 12, 72, -55, 21, -88, -11, -109, 118, -66, 106, -120, 99, -15, -17, -28, 90, -127, -75, 9, -83, -35, -90, 72, 124, -77, 10, 127, 11, 47, 120, 56, -98, -85, -87, 93, -38, 108, 52, 95, -120, -76, -59, 54, 64, 77, -100, 116, -58, -91, 33, 4, -28, 58, 57, -19, 31, -64, 16, 100, 24, -8, 58, -50, -56, -90, -119, -53, -3, -106, 12, 91, 78, -36, -89, 98, 66, 0, 24, -116, -105, -126, 124, 20, -39, 16, 58, -10, 35, -6, -97, -40, -83, -34, -6, -36, -94, 9, -112, 21, -76, 85, 71, -41, 107, -45, -40, 79, -98, 36, -96, -7, -103, 39, 88, -26, 68, -61, -58, 105, -53, -50, -54, -26, -121, -30, 99, -35, -82, -93, 78, -2, -114, 38, -57, -85, -89, -39, 79, 113, -45, 33, -66, -11, -92, -47, -20, -99, 27, 19, 14, 14, 24, 62, 95, 28, -46, -74, 65, 45, -108, -124, -127, 42, 41, -16, 81, -79, 22, 20, 125, -17, -116, -102, 25, 56, -38, -11, 26, 48, -114, 96, 32, -68, 5, -75, -103, 125, 79, 77, 43, 46, -125, -83, 42, -104, -90, -85, -42, 68, -85, -25, -2, -60, -72, 118, -3, 118, -30, 111, 28, -90, -78, 82, -55, -23, 98, 71, 51, -58, -94, -44, -24, 62, 112, 64, 116, -10, -101, -72, -35, -106, 97, 8, 34, -85, 33, -3, -89, -24, -82, -81, 37, 77, -92, 56, 34, 89, -115, 120, -29, -113, 58, -110, -69, -83, -2, 55, 14, 0, 69, 123, -92, -83, 83, -125, 63, 20, 28, 93, 53, 12, 88, -124, -126, 59, -51, 30, 116, 96, 46, 89, -54, 75, -64, -120, 118, 24, -31, -94, -38, -12, -74, -108, -44, 37, 92, -119, 83, 3, 17, 104, -79, -11, -87, 30, -106, -46, -60, 78, -68, -29, -91, 29, 0, -6, -80, -53, -117, 32, 106, 25, 52, -58, 58, -13, 114, -44, -128, -27, -110, -87, -42, 104, -59, 97, 123, -113, -9, -125, -117, 63, -63, 55, 24, 30, -75, 11, -120, 28, 68, -25, -28, 0, 77, 127, 52, -61, -88, -42, -57, -31, 75, 43, 39, -77, -63, 124, 58, -69, 13, -127, -73, 25, 122, -43, 32, -78, 100, -93, 109, -119, -27, 120, 111, -30, -76, -89, 33, 117, -14, -40, -113, -67, 124, -77, -30, 83, 1, 75, 114, -95, -70, 24, 57, -81, -51, -118, -111, 29, 47, -128, 58, 127, -37, 13, -121, -103, -45, 50, 94, -59, -2, -87, -57, 24, -7, 14, 22, 12, 64, -116, -76, 107, -120, 114, -4, 73, -61, -25, -39, -5, -93, -119, -103, 2, -18, -4, 33, 24, 74, 0, 81, 8, 122, 123, -55, -26, 15, 70, 87, 123, -42, -75, -92, -26, -63, -35, -48, -120, 97, -53, -87, 112, 84, 109, 26, -106, -119, 104, 14, -27, 24, -16, 96, -14, 68, 4, 66, -81, 48, -23, 12, -96, -53, -52, 62, -90, 88, -124, 119, 71, -30, 17, 29, 121, 71, 116, 121, 95, 118, -115, -34, 12, -104, 73, 113, 26, -115, -128, -27, 39, 28, -7, 106, -62, -16, 127, -11, -12, 122, 4, -112, 43, -5, -78, 2, -60, -23, -101, -57, -120, -43, -88, -31, -65, -8, -90, -74, 22, -44, -125, 34, -108, -63, -52, 124, -33, -76, 66, 61, 91, 31, 18, -19, 10, -8, 81, 68, 87, -61, 5, 84, 67, 109, 95, -128, 82, -32, 46, -99, 52, 73, 78, -54, 98, 43, -111, 50, 65, 36, -21, -100, 67, -15, -27, 53, 45, 104, -51, 69, -30, -82, -79, -26, -78, -48, -19, -12, -15, 28, -127, -82, 60, -118, 18, 62, 36, 90, 95, -108, -4, -68, 112, 117, -128, 112, -87, -100, 101, -42, 109, -84, 33, -53, -76, -3, 24, -98, 43, -10, -93, 4, 32, 117, 69, 104, 24, -122, -51, -21, 95, -30, -75, 1, -13, 39, 91, 123, 103, -10, 52, 24, 80, 23, -115, -88, 13, 16, -16, -128, -30, -65, 72, -76, 32, 71, 73, 83, 52, -35, -120, -78, 100, 76, -85, -93, 16, 31, 32, 116, 5, -128, 104, 51, -113, 44, 119, -85, 95, 119, -43, 84, -39, 63, 56, -44, 88, 119, -108, -27, -24, 17, 108, -40, -21, -63, 97, 6, 95, 0, -33, 111, -93, -120, 36, -41, 88, -7, -67, 86, -126, -12, 108, 83, 94, -5, 52, -90, 66, 34, -84, -123, 53, -104, 88, 78, 62, -81, 126, 116, 31, 91, 77, -73, -22, -103, 4, 87, -29, 94, 20, 100, 95, 65, 6, 83, 80, -76, 117, -124, 17, 24, 95, 99, -88, 55, 59, -112, 120, 95, 62, -3, 44, 9, -11, -67, 83, -116, -64, -16, -72, 98, 45, -14, -66, 13, 82, 8, 55, 31, -40, 0, 49, 4, 12, -108, -125, 65, 126, -6, -32, 21, 17, -1, -74, 5, -41, -97, -36, -20, -24, -123, 98, 117, 69, 65, 2, 110, 77, -49, 112, -48, 92, -95, 116, -58, -113, -81, -59, 74, 69, 62, -16, 68, 53, 79, -9, -48, 42, -117, -110, -126, -81, -83, -16, 34, -95, -97, -30, -65, -113, 68, 59, 54, 41, 5, 74, -14, -122, 16, 21, -11, -107, -95, -104, 16, 24, -19, 63, 15, -112, 5, 117, 102, 1, 66, 31, -66, -9, 106, -6, 119, -46, -49, -67, -20, -100, -27, -29, 66, -8, 113, -12, -13, -95, -26, 69, -4, 50, 62, 42, 80, -44, 58, -55, 3, -123, -12, -7, 110, -97, 100, 74, -128, -105, -64, -3, -39, 97, -6, 41, 35, 112, 36, -94, -41, 22, -104, -9, 15, 20, -113, -49, -71, -7, -65, 84, -89, -33, -94, -118, 17, -122, 58, 61, 4, -109, -47, -34, 47, -100, -110, 56, -70, -59, -48, 68, -41, 108, 76, 106, 47, -106, 66, -109, 20, 124, -9, -128, 43, -25, -46, 115, 99, 117, 103, -36, -9, 28, -34, 38, 50, -54, 62, 22, 85, 83, -50, -107, -121, -76, 9, 100, 96, -26, -74, -61, -36, -123, -51, -125, -33, -47, 23, -18, 123, 1, 118, -96, 48, 69, 87, -65, 57, 57, -25, -97, -55, -72, -39, -72, 106, -65, -39, 66, -112, 41, 47, -95, -21, 76, -26, -4, 25, 116, -94, -24, -7, -28, -127, 123, -44, 36, -97, -88, 113, 1, 111, -107, -104, 19, -58, -82, -47, -9, 58, 60, 69, -54, -69, 1, 64, 66, -77, -66, 6, 50, 111, -36, 22, 48, 68, 108, -28, -116, 81, -67, -7, -29, 89, 106, 87, 100, -81, 110, 14, -44, 35, -103, 80, -12, 90, -86, -118, -54, -37, -12, 96, -2, 48, -113, 77, -58, -124, -51, 124, 52, 118, 72, -126, -113, -72, 30, 125, -25, -48, -117, -80, -113, 20, -62, 1, 10, 46, 20, 26, -25, -81, -112, 48, -76, 88, -125, -45, 105, 16, 60, -7, -33, -52, -49, 81, 120, -42, 21, -62, 118, 116, -95, 31, 13, 53, -95, 123, -115, 52, -16, 100, -39, -1, 121, 113, 25, -3, 75, 69, 59, -126, -97, 8, -89, 32, -100, -121, -41, 121, -103, 63, 10, 86, -62, -89, -43, 47, -108, -45, 98, 14, -20, 112, 47, -96, 77, -30, -110, -71, 27, 84, 55, -109, -109, -118, -107, -122, -35, 115, 0, -120, 26, -71, 85, 71, -85, 61, 44, 85, -58, -90, 95, -11, 36, -44, 102, -28, 63, -103, 59, 21, -117, 15, 46, 127, -29, 126, 104, -6, -74, 99, -92, 114, -11, -97, 16, 72, -17, 103, -34, 105, 52, 104, 19, -18, -90, -78, 72, -46, 33, -56, 38, 90, -43, -10, 80, 107, -26, -66, -118, -49, 101, -90, -57, 85, 39, -86, -31, 114, 50, 11, -26, -64, -96, -47, 24, -12, 98, -27, -79, -24, -63, 28, -91, 32, -24, -101, 29, 19, 4, 75, -105, 3, -84, 58, 115, 3, -119, 16, 122, 75, -122, 91, 12, 47, -106, -73, 44, -114, -63, -96, -69, -109, -109, -61, 80, -16, -7, -65, 54, -101, 74, -88, -99, -49, 90, 92, -62, -127, 127, -84, -73, -124, -4, 4, -57, 64, -13, -28, 121, 86, -72, -20, 127, -13, -42, 109, 90, -97, 85, 89, -66, -26, 9, -70, 4, 23, 74, -75, 98, 37, 94, -100, 72, 85, 105, 112, -26, -50, 2, -43, 36, -77, 49, 26, 11, -17, 43, -95, -97, -104, 7, 122, -8, -49, -47, -68, -107, 31, 116, 57, 86, 34, -90, -41, -103, -29, -108, -117, 109, 119, 44, 85, -103, -7, -92, 116, -73, -88, 83, -62, 43, -51, 1, 52, 36, -46, 116, -74, -72, 29, -13, 30, -6, -101, -55, 120, -58, 127, -119, 70, 45, -114, -19, 86, 117, -37, -3, -80, -63, 109, 15, -43, -74, 20, 115, 40, -79, 113, 37, -112, 78, -74, -101, 3, 9, 98, 59, 106, 17, 110, 75, 3, 6, -123, 53, -45, 98, 61, -67, -114, 38, -89, -9, -91, -24, 78, -70, -71, -84, 46, 93, 25, 112, -11, -70, -89, -51, 125, -89, -59, 29, 5, -85, -4, 111, 123, -118, 0, -106, -77, -104, -28, 13, -51, 64, -93, -96, -75, 14, -79, -9, 118, -33, -68, 56, 53, -6, -77, -39, -45, -40, -116, -58, -112, -70, -109, -125, 21, 55, 4, -103, 92, -91, 120, -78, 39, -68, 107, 55, -44, -26, 71, 63, 93, -101, 58, -58, -84, -7, 70, -84, 36, -55, 31, 30, 15, 52, 79, 64, -88, -40, -17, 45, 13, 116, -22, -112, -11, 111, -59, 102, 51, -6, 101, 19, -55, -112, -83, 55, -109, 8, -7, 38, -40, -15, -38, -44, -85, -100, -81, 32, 123, -90, 7, -122, -84, -64, 123, -41, -26, -52, -29, 46, -119, 51, -26, 14, -49, 69, -72, 11, -116, 48, -118, 73, -38, -111, -100, 43, -108, 68, -2, -3, 20, -81, -58, 92, -9, -118, 69, -104, -26, -96, 46, 0, -44, -66, -15, 46, 105, -20, -33, 20, 126, -73, -44, -30, 3, 109, 42, -49, -113, -87, -49, -70, -123, -48, 93, 105, 94, 86, -34, -45, -110, -23, -118, 83, 48, -72, 57, -125, -91, -66, -63, -47, -1, 20, 100, -67, -28, -113, -31, -69, -85, -116, 127, -20, 104, 48, 42, 37, -109, 26, 113, 6, -107, -4, 54, -38, -12, -52, 113, -62, 34, 8, 97, -86, 32, 107, -68, -96, 3, -14, 80, 97, 31, 71, 124, 13, 106, -114, -21, 44, 99, 28, 116, -39, -76, 45, -3, -8, -59, -25, -11, 125, -18, -14, 121, 27, -115, -127, -101, 28, 124, 56, 112, 125, 76, 83, 71, 103, -119, 124, 60, -20, 49, 117, 15, -29, -47, 121, -92, 20, 122, 111, 121, -54, 6, 16, -1, 87, 96, -106, 46, 107, -38, -52, 84, 36, -97, -19, 95, 7, -87, 13, -82, 91, -46, -7, 101, -89, -109, -43, 126, -102, -64, 75, 14, 8, -16, -73, -51, -14, -97, 100, -11, 45, -74, 19, 114, 109, -14, 23, -74, 127, -117, -62, -33, -10, 14, -125, -48, -124, 76, 31, 97, 76, -21, -23, 69, -67, -110, 81, 80, 93, 28, -84, -12, 126, 123, 39, -2, 107, 5, 14, -8, 70, 41, -108, 10, -74, -59, 61, 52, 11, -108, 113, 74, 114, 14, 34, -64, -24, 29, 42, -46, 81, -71, -77, -66, -62, -54, -74, 46, 4, -28, 15, -122, 93, 0, -54, -8, 82, 76, 6, -61, 29, 72, -106, 108, -127, 37, 71, -66, 16, 72, 60, -78, 51, -108, 30, 45, -67, 1, -83, 13, -55, 22, 15, -113, 24, -24, 46, -66, 4, 2, 57, -60, -36, -108, 78, -22, 50, -124, -84, 4, -54, -78, -2, -75, -64, 121, -49, -5, 32, -123, 32, 81, -44, -110, -73, -117, -5, 77, 34, -88, 25, -94, -68, -78, 1, 26, -46, -2, 14, 40, -115, -92, -38, -55, -125, 11, 60, -36, 94, 77, -110, 14, 117, 75, 1, 48, -61, 20, 75, -15, 17, 73, -126, 0, -83, 68, 42, 62, 33, 77, -114, 80, -121, -69, -5, 75, -47, 13, -59, 93, 35, 37, 93, -126, 19, -115, 118, -97, -93, -119, 78, -37, -125, -111, 63, 54, 73, 50, -44, -111, 40, 15, 112, 16, -46, -92, -8, -18, -83, -1, -34, -100, 29, -28, -67, -48, 32, -102, -93, -73, -51, 76, 2, -4, -110, 120, -114, -43, -6, -126, -105, 4, 90, 61, 38, 19, 68, -50, -101, 55, -19, 30, -116, 120, 49, 27, 80, 91, 76, -27, -49, -124, -59, 53, -84, 18, 79, 69, 114, 126, -49, 105, -12, -57, -114, 127, -64, 25, -59, 120, -97, 45, 8, 56, -67, -36, 102, -106, -34, -12, -63, -48, -96, 121, 11, 119, -89, 27, 79, 78, 93, -34, 73, 113, -120, -97, -24, -38, 104, 2, -58, 26, -77, -32, -59, -116, -6, -22, -106, 34, -16, 65, -97, -90, -44, 91, 99, -11, 73, -99, -79, -37, -112, -73, 99, -105, -44, 75, -32, -108, 18, 119, 83, 90, -118, 122, 79, -4, -97, -1, -16, 110, -57, -101, 113, 103, 108, 96, -20, 37, -29, -85, 126, 112, -65, -94, 126, 12, -11, -87, 88, -12, 51, -25, 8, 127, 110, 33, 57, 84, -66, 41, 118, 79, 94, 93, 120, -118, -94, 103, 103, -28, 65, -84, 111, -114, -50, -59, -8, -116, 122, -21, -90, -112, 83, 24, -46, 13, -78, 108, 27, -7, -125, 43, -74, -83, 7, -118, -93, -1, 92, 98, -120, -79, 86, 41, -105, 69, 3, -58, -89, 52, -117, -99, -53, -118, -100, -56, 81, -38, -99, 33, -52, 80, 127, 18, -48, 115, -23, 115, -122, -35, 106, -46, -7, -40, -100, 69, 67, -7, 67, 22, 21, 50, -20, 35, -113, 105, -11, 97, 8, 81, 0, -78, -11, 8, -20, -93, 53, -6, 52, -56, -122, 16, 56, 51, 124, 118, 101, -11, -29, -88, 95, -28, -112, 0, 83, 4, 15, 17, 70, 99, 43, -76, -76, -56, 43, -112, -65, -85, 29, 98, 28, -43, 119, 89, -44, -122, -77, 119, -84, -50, 93, 11, -34, -82, 94, -60, -45, -109, 60, -62, 3, 79, 94, -23, -61, 72, -21, 67, -34, -88, 75, -63, 57, -24, -30, 72, -23, -6, 58, -124, -113, 52, 81, 8, -83, 87, 97, 20, 12, 111, -35, -50, 25, 123, 23, 68, -6, 64, -10, 74, 48, -58, -74, 43, 58, 25, 97, 20, -88, -82, 28, 6, -62, 54, -58, -80, 116, -58, 78, 118, 127, 36, -86, -37, -39, 2, 18, -50, -4, 101, -47, 66, -22, 125, 118, -28, -10, 21, -46, 7, 104, -4, -23, 11, 62, -39, -95, -75, -68, 38, 72, -41, 23, -34, -51, -7, -100, 48, -26, -31, 120, -31, 62, 60, -90, -116, 100, 105, -22, 33, 3, 19, 48, -22, 46, -34, -77, -69, 100, -15, 19, -94, 32, -87, -121, 73, 78, 52, -22, 45, -17, -109, 63, 118, -67, -39, -65, 87, -14, 114, -107, -46, -67, 95, 110, -95, 108, -91, 23, 45, -75, -19, -36, 88, -79, 39, -35, -18, -73, 35, -12, 42, -81, -98, -99, 10, -78, 83, -32, 42, -9, -120, 49, -114, -72, -16, 126, 33, -7, 12, -84, -95, 83, -67, -74, 82, -35, 54, 35, -105, 38, -50, 14, 61, -122, -120, 50, 112, -79, 59, 1, -66, -40, -121, -96, -89, 35, 22, -20, 84, -39, -37, -4, 123, 12, -30, 111, 99, -63, -108, 3, 89, -109, 120, 13, 55, -99, 51, 47, 98, -18, 86, -126, 108, 3, 95, -105, -45, -118, 122, -23, 105, -102, 21, 67, 64, 45, -118, 30, -81, 95, 41, -80, -15, -60, 117, -5, -122, 15, -107, -103, -105, -25, 102, -91, -85, 40, 106, 104, 98, 77, -100, 3, 100, 25, -79, 7, 93, 74, -24, 97, -19, -91, -39, -21, -120, 127, -54, 36, 46, 88, -4, 50, 48, 65, -65, -53, 14, 90, 37, 31, -17, -128, 104, 32, 30, -72, 11, -11, 97, -90, -56, -120, -100, 118, 14, -100, -33, 44, -36, -69, 76, -40, -103, -114, -114, 92, -98, -42, 52, 118, -77, 113, -69, -77, -71, 50, -43, 42, -122, -124, 71, -91, -1, 47, -116, 97, 126, 29, 9, 82, 113, -111, -40, -20, 86, 27, -10, -44, -112, -29, -71, 39, 125, -33, 112, -123, 74, -92, -21, 87, 120, -53, -112, -56, -4, -48, 84, -33, 34, -10, 37, 17, -108, 37, -128, -51, 86, -77, -94, 57, 93, -52, -21, -124, -26, 71, -21, -106, 72, 81, -54, -38, -89, 90, 84, -127, -88, -28, 120, -28, -116, -2, 57, 47, -37, -53, 17, 58, 7, -28, -93, -50, -2, -43, 82, -51, -84, -36, 80, 16, -93, -71, 57, 30, 112, 107, -28, -27, 22, 32, 127, -51, -90, -48, -106, 126, 123, 9, -97, 76, -96, 31, -25, 93, -77, 70, 64, -9, 44, 57, 35, 70, -65, -27, -82, -47, 14, -15, -88, 37, 59, -98, -2, -78, -25, 10, 15, 85, -71, 115, -59, 30, -20, 19, 64, -24, 125, -5, -63, -120, 10, 79, -106, -12, -115, -39, -23, 51, 66, 80, -80, -47, -90, 58, -2, -115, -22, -20, -105, -121, 106, 41, -74, -53, 45, 103, -77, -98, 57, 126, 7, 28, -67, 3, 122, -53, 19, -37, 80, -93, 108, -30, -108, -50, 77, -74, 71, 116, -96, -17, -23, 64, -83, -60, 45, -93, -66, 55, -38, 119, -123, 54, 93, -85, 93, 121, -17, 120, -30, -18, -6, -30, -16, 120, 4, -47, 88, 120, 64, 86, -80, -8, -47, -49, 112, -102, 76, -43, -46, -71, -7, -90, 81, 126, 119, -3, 77, 59, 44, 119, -95, 44, -118, 26, 46, 46, 17, 2, -21, -50, 36, 122, -13, -6, 26, 19, -46, 11, 105, 118, -38, 27, -114, 19, -4, 115, 65, 15, -8, 77, 121, 107, -29, -65, -59, 35, -104, 95, 110, -72, -120, -65, 22, -88, -37, 75, 14, -128, -108, -15, 47, 3, 118, -96, 21, 127, -26, -59, 58, -27, -120, -21, 19, 74, 75, -84, 46, 2, 19, -77, -44, -42, -23, 90, -53, 84, 4, 4, 16, -21, 54, 60, -116, -81, -116, 60, 41, 44, 121, -65, -48, -100, -39, 64, -117, -69, -30, -38, -82, 85, -106, -16, -67, 14, -36, -46, 112, -25, 46, -120, -35, -11, -73, 48, 93, 29, 74, 35, -80, 102, 47, -123, 6, 49, -76, 19, 87, 10, -26, -65, 0, 102, 11, -102, -63, 18, 44, -52, 120, -102, 71, 71, 32, -37, 7, -32, -22, 119, 82, 99, 25, 13, 117, -128, -74, -23, -6, 63, 17, 105, -112, -45, -18, 16, -46, 59, -119, 125, -48, -14, -53, -10, -69, 42, 3, 69, 38, -53, -89, 71, 48, -1, 118, 38, -48, -84, -102, 11, -15, -5, -56, -48, 1, 70, 122, -80, 80, 111, -121, -72, 93, -119, 39, -19, 47, -123, 34, -117, 112, 10, -4, 50, 1, -49, 111, -105, 65, -115, 127, 114, -111, 66, 65, 26, -21, -92, 55, -70, 103, 85, 67, -103, -16, 108, -46, 80, -97, -33, 107, -90, 111, 47, -10, 95, -55, 18, -60, 12, -52, 104, -81, -106, -67, -125, -55, 3, -6, 68, -105, 120, -106, -123, 6, -90, -108, -117, 47, -89, 116, -47, 11, -31, -94, 63, 7, -118, 3, 8, -9, 57, -22, -19, 79, 88, -64, 13, -37, 75, 12, -27, -103, -77, 16, 27, -105, 106, -126, 83, 20, 84, 24, -21, -58, 67, 53, 26, -122, 84, -21, 65, 16, -21, -60, -119, -107, -87, -57, 116, 13, 59, -31, 97, 108, -18, 40, -92, 108, -124, -106, -115, -89, 87, -66, 121, 13, -86, -23, 4, 102, 29, -10, 74, 45, -123, 77, -39, 124, -96, -19, 121, -43, -108, 58, 30, 117, 109, 63, -51, 80, -86, 9, -20, 101, -77, -50, -72, -79, 111, 67, -76, 55, 125, -60, 46, -40, -83, -39, 56, 37, -88, 110, -112, -13, -80, 111, 42, -44, 14, 108, -65, 46, 84, 48, -109, -98, -15, -57, -105, -41, 25, -96, 96, -4, 11, -56, 14, -122, 101, -116, 27, -100, 109, -22, 125, 104, -6, -8, -89, 56, 5, 52, -104, -46, 117, -87, -2, 81, 37, 62, 36, -75, 103, 114, 115, -106, 123, 60, 59, -16, 35, -123, -104, 115, 72, -72, -81, 81, 22, -31, -55, -92, -126, 92, 124, 126, -71, 38, 60, -35, -72, 124, -19, -100, -92, -7, -20, -60, -123, 38, -96, -26, 16, -123, -125, -75, 99, 78, 4, -22, 47, 86, -37, -107, -31, -51, 54, -118, 51, 30, 87, -113, 123, -108, 53, -4, -28, 70, -100, -48, -123, 53, -91, -67, -119, -97, -60, -10, -104, 84, 42, -19, -50, -68, 30, 97, -10, 94, -62, -121, 8, -33, 58, 124, -119, -69, -16, -127, -49, -27, 95, 9, -64, 80, 0, -128, -90, 49, -100, -40, -2, -12, 95, -121, -12, -23, 16, 93, -50, 1, -63, 42, 49, -127, -23, -30, -11, -27, -98, 88, -76, -26, 9, 47, 76, -27, -63, -25, -1, 90, 24, 118, -43, -27, 74, 101, -110, 41, 57, 120, 12, 10, 60, -64, 117, 57, 56, 69, -106, 100, -71, -102, 41, 26, -72, -51, -89, 33, -76, 111, 22, -8, 1, 102, 106, -63, -83, -5, 125, -77, 28, 90, -103, 16, 99, 56, -23, -83, 83, -2, -39, 127, -66, 68, 115, -63, -71, -37, 77, 55, -80, 87, 116, 49, 19, 107, -91, 55, 45, -27, -99, 53, 115, 124, 76, -57, 98, -75, -47, -94, -74, 103, -93, 11, -1, 20, 90, 87, -33, 22, 52, 14, 81, 62, -5, -120, -103, 63, 54, 37, -128, 69, -100, -91, -119, 68, 9, -98, -112, -101, 66, 78, 43, 77, -65, -85, -44, 75, 77, -117, -12, -19, 57, 12, 8, 45, -87, 14, 60, -46, 29, -75, -94, 36, 98, 80, -40, 108, 116, 76, -1, 66, -9, -3, -57, -125, 71, 62, 93, -10, 59, -120, 114, 73, -55, 118, -7, 123, 87, 25, 73, -107, 122, 110, 119, -63, 117, 99, 127, 85, 54, -5, -40, -34, -120, 9, 118, 3, 87, -83, 50, 78, 67, -5, 83, 97, -110, 11, 81, -101, -94, -83, 91, -9, 5, -35, -85, 26, 116, -28, -1, 76, 26, -112, -83, 22, 121, -29, 83, 3, 10, 70, 96, 67, 89, -52, 63, 66, -127, 41, -112, 63, 100, 46, 39, 15, -12, -108, -100, -81, -86, 72, 23, 99, 64, 79, -62, 104, 4, 88, 27, -82, -37, 21, 21, -105, 113, 90, -85, -75, 81, -19, -20, 101, -26, -90, 72, -96, -71, 121, -7, -67, -46, -82, 97, 16, 112, -32, 108, -100, 91, -35, 107, -34, -90, -60, 7, -38, 112, -111, 127, 98, 76, 53, -25, 25, 121, -5, 48, 115, 1, 122, -91, -6, -81, 123, -67, 78, 33, -14, -108, -44, 48, 108, 36, 25, 62, 91, 61, 106, -128, -88, 118, -10, 32, 52, 14, 103, 44, -58, -52, -95, -112, 32, -22, 102, 88, -77, 77, 90, 78, -14, 122, 1, -107, -70, -99, 125, 92, 96, -97, 75, 26, 55, -5, -47, -126, 4, 42, -106, -81, -8, -121, 120, -35, 109, 107, 48, -87, 55, -12, 10, 23, -60, -64, -13, 112, 34, 55, 92, -88, -115, -79, -64, -74, -121, 75, 49, 46, -56, 62, -42, -105, 5, -69, -60, -48, 81, 1, 66, 96, 110, -78, 60, -102, 71, -1, 21, 21, -121, -43, 17, -79, -59, -99, 90, 75, 8, -18, 110, 78, -23, 11, -97, 33, -29, -49, 41, -41, -80, 20, -45, -55, 17, -20, 28, 89, -97, 17, 15, 100, -47, -39, -59, 75, 34, -91, 76, 103, -75, 51, 16, 48, 58, -25, -53, -15, -112, -27, 65, 73, -125, 110, 96, -88, 24, -43, -67, 69, 44, -30, -22, 74, 46, -42, 62, -14, -114, 0, 114, 85, 77, -116, -104, 109, 98, -76, -9, 118, -39, 69, 74, 7, 4, -121, 114, -37, 77, -110, 54, 76, 76, 30, 125, 37, -69, -39, -81, -61, -116, 106, -7, 123, 47, -10, -71, 79, -45, -109, 23, -49, -111, 72, -126, -60, -73, -22, -21, -51, -44, -53, -87, 45, 111, 65, -110, 81, -85, 116, -62, 82, 106, 55, -9, -17, 3, 121, -20, 26, 65, 23, -74, 104, -33, -123, -115, 36, -126, -59, 4, -101, 99, -12, -119, 111, -26, -76, 59, 41, 119, 71, 59, 15, -9, -96, -23, 93, 56, -26, 21, -7, 102, -113, 16, 52, -38, 60, 97, -11, 51, -91, -75, -61, 43, -21, 113, -89, 16, -11, -91, 73, -68, 74, -5, -73, 64, 56, -97, 111, 31, 45, 110, -80, -118, -14, 64, 103, 118, 73, -14, -78, -58, 78, 7, -126, 35, -114, 105, -40, -6, 18, -125, 35, -80, -76, 56, 21, 92, 65, -98, -91, 92, 76, 109, -118, -26, 67, -84, -102, -18, 29, -16, 75, 66, 37, 83, -125, -93, 80, 119, -81, -33, -46, -2, -40, 16, -53, -28, -128, 50, -31, 26, 105, 114, 60, -34, -66, -120, 16, -62, -21, -51, -27, -16, -36, 121, -1, 100, -18, -24, 59, -74, 111, -91, -84, -91, -35, -66, 83, -124, -33, 127, 98, -2, 109, 93, -33, -80, 19, -127, 6, -103, 87, 50, 95, -97, -60, -28, -128, -73, 82, 20, -50, -91, 39, 57, 20, 20, 70, 47, -70, 60, -28, -23, -61, -13, -100, -65, 36, 17, -105, 98, -108, -69, -35, -19, 19, -127, 55, 54, 97, -83, -82, -118, -17, -96, 63, -13, 1, 50, -27, 78, 36, -7, -62, 39, 65, -2, 85, 36, 108, -120, -36, 96, 126, -73, -33, -44, -45, -106, 31, -32, -52, 98, -32, -113, 59, 55, -85, -13, -123, -60, 7, 15, 67, -42, -4, 4, -120, -51, -63, 28, 75, 48, 0, -44, 53, 90, -86, -12, -98, -86, -93, 107, -112, 52, 126, 92, -70, 0, -23, 60, -67, -115, -54, -46, 114, 29, 93, -78, 88, -82, 79, 8, -22, -30, 32, -53, -78, 40, 5, -53, -52, 64, -79, 28, 126, 10, 121, 49, -33, -98, -4, 110, -41, -32, 57, 125, -26, -9, -12, -113, -90, -108, -65, 16, 118, -42, 65, -47, -108, -10, -85, 32, -128, -89, -112, 84, 105, 18, 87, 86, -11, -3, 78, -58, -46, -32, 44, -113, 105, 104, 54, 27, -118, -111, -79, 87, -54, 3, 74, 74, 69, -3, 26, -98, 106, -42, 101, -76, -128, 65, 1, 66, 46, -125, 4, -79, 6, -25, -93, 53, -18, -125, -27, -46, 107, -62, 86, 24, -79, 125, 34, -63, -49, -42, 6, 82, -25, 83, -100, -115, 127, -98, 37, -18, -89, -82, -91, -41, -106, 57, 23, 72, 126, -105, 14, 6, 90, 83, 95, 33, -26, 80, 32, -100, 127, 100, -90, 100, -53, 65, -65, -36, 97, -128, 94, -80, -35, -52, -14, 29, -21, -22, 111, 19, 26, 106, -21, 45, 37, 68, -21, 88, 106, -63, 42, 58, 108, 41, -11, 24, -1, 43, -87, 12, -97, -36, -73, 84, -26, -125, -120, -96, 127, -25, 96, -58, -75, -97, 117, -96, 45, -93, 67, 117, 15, -66, 94, 42, 85, -95, -27, -97, 47, 119, 36, -21, 24, -9, -25, -92, 74, -108, -13, -93, 3, -92, 93, -26, 17, -20, -106, 36, -81, -127, -61, -94, 120, 95, -52, -11, -77, 32, 11, -71, 10, 122, 103, -82, -34, 95, -103, -81, -66, 14, -87, -76, -67, -84, 23, 23, 50, -2, -32, 122, -60, -117, -115, 44, 114, -84, 107, -76, 0, 51, 3, -71, 101, -23, -32, -115, -60, 17, -88, 59, -39, 40, 40, 41, 68, 15, 68, -26, 39, 58, 115, 55, -26, -81, 24, 7, -108, 110, -91, 36, 69, -70, -103, -68, -67, 50, -47, -115, -53, 32, 33, 70, -67, -120, -82, 50, -57, -93, -121, 64, -8, -115, -99, 54, 107, -127, -117, 22, 111, 57, -122, 86, 126, -3, -109, 124, 25, 120, -91, -91, -13, 82, -74, -38, -63, 112, 23, -23, -86, -112, -18, 111, -31, -17, 78, -6, 63, 80, 27, 9, -90, -85, -118, 92, 123, -29, -92, 100, -18, -79, -32, 67, -7, 89, -30, -111, 67, -79, -36, 59, 2, 31, 34, -119, -124, -90, -106, 40, 25, 113, -73, -77, 123, 114, -125, 114, 15, 88, 90, -123, 34, 52, -8, -63, 92, -48, -11, 79, 127, -27, 59, 64, 94, -88, -120, 100, 1, 30, 13, 111, -23, 105, -12, 80, -116, 24, 23, 78, 49, -100, 94, 6, -89, 41, -17, -35, 92, 24, 76, 22, 28, 0, 19, -90, -107, 87, -78, 11, -128, 103, 15, -35, -42, -66, -34, -114, 87, 3, -53, 13, 124, 24, -2, 18, 14, -78, 87, 62, 0, -127, 38, 25, -59, -79, -128, -54, -10, 43, -119, -105, -1, -113, -95, 124, 25, -27, -14, -94, 50, -124, 4, 29, 66, 24, -16, -6, -20, -38, 50, -123, -99, 87, 17, 119, 114, 16, 40, -28, 113, 94, -8, -7, 83, 55, 122, -95, -61, -46, 30, 99, -46, 47, 101, -107, 57, 85, 46, 93, 87, 93, 120, 103, 25, -98, 32, -102, -114, 56, -72, -37, 123, -60, -49, 47, 38, -64, -122, -123, 64, 97, 110, -3, 6, 115, -29, -100, -101, -126, -19, 28, 91, 104, -21, -42, -60, 110, -69, 78, -45, -26, 98, -121, -41, 104, -62, 21, 75, 107, 103, -33, -80, -28, 8, -28, -22, -36, -112, 16, -127, -36, -120, 20, -1, -2, 85, 36, 55, -15, 5, 120, -117, -21, 19, -93, 42, -115, -28, 90, -46, -5, 122, -7, -12, -32, 72, -44, -123, 81, 30, -55, -24, -57, -122, -28, 70, 82, 35, 110, 44, -23, 86, 41, -104, -122, 16, 30, -17, 125, 107, -2, 76, -53, 62, -34, 32, 69, -66, -31, 112, -79, -75, 52, 46, -97, -75, -56, 111, -2, -39, -64, -109, -69, 28, 35, 36, 30, 47, 76, -78, 38, -46, -51, -112, 83, 96, 109, 109, 48, -6, -99, 19, -17, 15, -11, 88, -94, -41, -11, 52, 118, 9, -60, 28, 50, -92, 105, 90, 52, 51, 67, 6, -49, 82, -94, 85, -100, -62, 70, -102, 41, -115, -43, 98, -79, -29, 73, -77, -68, 104, -86, 83, 7, -48, -70, -67, 102, 22, -114, 103, -126, -108, 8, -67, -66, -64, 70, 61, 101, 112, 91, -105, 102, -89, 110, -95, 101, 3, 4, 41, 23, -41, -87, 63, -94, 18, -9, -35, 28, -60, 67, -97, -119, -32, 85, -104, -24, 51, 30, -91, -2, -1, 47, -110, 58, 32, -39, 42, 28, 82, -58, -98, -85, 124, -62, -19, 115, 11, -88, 17, 116, -20, -7, -88, 127, 58, 97, 107, 103, -106, 101, -46, 15, 29, -13, 98, 79, 54, 2, -78, -11, -55, -58, -6, -6, 13, 90, 92, 118, 92, 17, -87, -2, -43, 82, -40, -124, 77, 70, -17, 122, 97, -75, 107, 113, -97, -9, -42, 38, -58, -45, 109, 73, -52, -32, -22, 115, -106, 102, 78, -20, -40, 33, -46, 70, 78, -4, 38, -94, 22, -125, -7, -19, 15, -17, 19, -28, -86, -12, 14, 6, -28, 45, -92, -70, 124, 80, -110, -71, 54, -3, -101, 51, -79, 65, 4, 17, 79, 60, -62, -63, -31, 127, -113, 84, 1, -66, -29, -71, -84, 91, -76, 83, -71, -2, 110, 68, 68, 124, -10, -5, -117, -66, -34, 113, 107, 29, 29, 12, 0, -38, 8, 98, 127, 104, 37, -72, 16, 110, 126, 82, -66, 94, -76, -115, 109, 39, -127, 70, -84, 20, -124, 80, 121, -101, -71, -61, 125, 55, -89, -54, -22, 5, -106, 32, -93, 74, 54, 21, -30, 19, 51, 120, -76, -85, 60, -29, -120, 115, 28, 37, 19, 114, -4, 102, -106, 12, -15, -54, 64, -69, 34, -50, -42, 3, -55, -126, 9, 68, -99, -110, -36, 69, -124, 15, -68, 55, -57, 98, -126, -24, -66, 50, -34, 120, -50, 62, 99, 97, 49, 26, 99, 115, 74, -4, 93, -62, 35, -71, -49, -83, 122, -16, -80, -27, -90, 78, 71, -74, 73, 53, 68, 41, -13, 28, -110, -53, -24, 118, -91, 126, -39, -61, 53, 44, -116, 77, -84, 72, 28, 98, 62, 104, 84, -69, -88, -58, 34, -47, 100, -96, 104, 125, 100, -28, 16, -93, 89, 90, -98, -63, -97, -20, -114, -124, -98, 85, -66, -92, -55, -51, -73, -121, 25, 108, 107, -7, 37, -118, -42, -125, 7, 50, 57, 11, -62, -110, 108, 125, -82, -35, 89, 117, -113, -24, 20, -35, -45, 117, -4, -128, -13, 117, -34, 125, 110, -126, 116, -12, -37, -60, -45, 114, 53, 72, 30, 67, 61, -40, -53, 41, 95, 7, 100, 4, -6, 4, -88, -19, -24, 86, 76, 72, 26, -63, -55, 38, 3, -105, 74, -91, 49, -58, 20, -50, -35, -20, 122, -68, 123, -123, 86, -25, -30, 72, 50, -54, 93, -69, -32, 16, 67, -7, 123, 33, 59, -10, -57, 58, -52, 99, 117, -49, 7, -1, -87, 108, -44, -64, -95, -84, 110, 30, -123, -75, -70, -63, -21, 125, -88, 61, -19, -115, -55, -37, -33, 42, 87, -89, 124, -80, -96, 33, 11, 120, 93, 99, -89, 89, 5, -27, -3, -67, -45, 85, 22, 20, 98, -36, -108, 42, 103, 63, 34, 123, 84, -7, 60, -9, 123, 33, -92, -18, -58, -13, 74, 11, -93, 46, 109, 10, -17, -42, 76, -36, -79, 110, -24, -100, -13, -61, 65, 63, -74, 10, -27, -95, -8, 85, -11, -104, 29, -1, 51, -53, 111, 36, -101, 14, -15, -66, -104, 93, 50, -89, 87, -46, 56, 70, 34, 10, -27, -36, -55, 13, -4, -31, -94, 119, 67, -43, 26, -61, 84, -98, -104, 30, -79, 40, -44, -19, -57, 70, 25, 119, 99, 58, -39, 7, -67, 1, 12, 73, -28, 101, -32, 73, -55, -33, 52, -52, -66, 69, 19, -103, -28, -68, -2, 92, -119, -24, 53, -116, 53, 123, -46, -9, 33, 0, 13, 106, -102, 10, -79, -95, -63, -105, -126, -21, 104, -38, 117, 25, -87, 8, 40, -117, -48, -122, 91, -127, -108, -72, -96, -1, -17, 101, -48, 25, 120, -128, -115, -52, -79, 62, -97, 37, 70, -42, -80, -86, 68, 17, -128, 84, 44, -48, -86, 51, -97, -18, -45, 47, 76, -126, -96, -5, -38, 46, 13, 13, -66, -4, 24, 54, 112, -79, 9, -74, -71, 109, 57, -47, -79, -4, 54, -8, 85, -33, 86, -15, -97, -22, -70, -36, 121, 115, 86, 39, -22, 113, -44, 66, -87, 75, 15, 125, 97, 23, 71, -110, -125, -36, 16, -38, 97, -74, -115, -66, 57, 28, 6, 91, -36, -61, 66, 6, -16, 117, 87, -30, -76, 106, -58, 53, 54, 70, 25, -83, 57, -29, 7, 108, 27, 6, 62, 21, -112, 48, -41, -2, -121, 8, -19, 87, 26, -97, 58, 114, 56, 35, 39, -20, -94, 9, -46, 17, -86, 4, -23, 12, -22, -66, 108, -108, 18, -44, -88, -49, 7, -41, -6, -121, 44, 10, 123, 55, 56, -79, 3, 44, -128, -26, -41, 108, 126, 55, 72, -95, 79, -123, -65, -102, 46, 27, 63, -119, -115, -18, -19, -126, 41, 40, 78, 118, -73, 97, 108, -8, 113, 29, 37, -38, 35, 6, 92, 123, -81, -49, -124, -32, 124, -127, 111, -109, -13, -35, 127, -92, -85, 0, -26, -87, -126, -55, -114, -35, 22, 57, 72, 8, -12, -75, 120, -5, 57, 48, -37, 3, -26, 33, 63, 62, -96, 78, 2, 90, 66, -105, -84, 72, 28, 126, 11, -55, -19, -91, 108, 3, 63, -70, -28, 125, 33, -125, -72, 110, -77, -39, 22, -91, 1, -25, 63, -96, 64, 92, 2, -17, 71, 122, -125, 1, 31, 74, 14, 8, 117, 80, -113, 94, 11, -101, 58, -23, 52, -122, 100, -93, -80, 31, 34, 26, 2, 99, 20, 23, -17, 6, -113, -78, -69, 79, 60, -56, -33, 120, -68, -125, 106, -38, -32, 85, 67, 14, -109, -10, 115, -71, 107, 71, -27, -18, -89, 89, 94, -69, -78, -121, 124, 103, 105, 34, 67, 83, -63, 33, 12, 117, -63, -41, -111, 19, -78, -86, 48, -122, -100, 8, 34, -94, 1, 77, -42, 32, 14, -69, -91, -54, 40, -96, 70, -38, -62, 14, -111, 39, 56, 79, -10, -30, 31, -111, 8, 108, 111, 4, -53, 73, -78, 114, 74, 41, 95, 89, 72, 122, -32, -114, -2, 79, 28, -118, 42, 62, 100, 2, 27, -12, -68, 93, -118, -27, 31, 46, 36, 33, 19, 54, -117, -124, 14, 121, 57, 117, 53, 60, -59, -89, 47, 0, -25, -6, -14, -83, -115, 127, 97, -21, -116, -58, -89, 90, -81, -66, -127, -35, -31, 126, 88, 112, -51, -4, 99, 58, 101, -103, 64, -3, 25, -24, -92, 9, -44, 104, -126, 56, 107, -108, -13, 64, 103, -31, 28, -101, 115, 127, -4, 46, 127, 118, 70, 87, 43, 87, 122, -71, 62, -71, 56, 75, -126, 7, 115, 84, 103, 74, -51, 19, -26, 121, -71, 75, 65, -19, -10, 95, -4, 93, 91, -111, 43, 16, -126, -84, 76, -62, 72, 9, -78, 28, 127, -112, 127, 72, 38, 61, -82, 125, 82, 114, 44, -36, 54, -63, -97, 78, 127, -26, -68, -124, -76, 24, 94, -122, -53, -102, 110, -3, -113, 34, -124, -108, 59, 23, -26, 16, 90, -24, -62, 125, -31, -40, -23, -35, 66, -44, 64, -95, 53, 19, -7, 83, -11, 73, -26, -128, 19, 113, -9, 58, -85, 99, 111, -53, 24, 42, -52, -109, -111, -91, 52, -53, 109, -37, 0, 116, 120, 21, 76, 54, -18, 8, -125, 24, -22, -74, 127, 115, 53, -43, 58, -10, -97, -67, 54, 57, -91, 82, -45, -45, 44, -121, 44, 121, -118, 111, 40, 8, -27, 78, -14, -64, -67, 52, 45, -88, 89, 45, 59, 37, -17, 14, 110, -5, -95, 122, -72, -117, 58, 17, -92, -103, -74, -108, -39, -16, 18, 8, -3, 77, 103, 28, 125, -32, 121, -110, 75, -51, 103, 96, -126, -68, -46, 57, -91, -39, -68, 54, 57, -6, 84, 87, -128, -98, 115, -10, 124, -23, 100, 17, 85, 49, -33, 35, 25, 40, -110, -70, 9, -1, -110, -55, -65, 61, -107, -55, 123, 10, -91, 97, -93, 92, 19, -25, 31, -48, 102, 8, -89, 95, -63, 109, -34, -11, -112, 96, 67, 86, 54, -120, 33, -103, 50, 34, -33, 24, -71, -11, -20, -22, -126, 58, 103, 42, 48, 33, -34, -81, 79, -26, 3, -2, -111, 121, 74, -76, -18, -48, -21, -45, 85, 9, -105, 71, 85, 11, 92, -98, 26, -45, -102, -84, 39, -37, -32, 82, -58, 26, -117, -28, 74, 116, 89, 94, 85, 47, 94, 0, 53, -71, 36, 51, 89, -91, -5, -47, 96, 35, -20, -24, -10, 116, -23, 60, -51, 127, 70, 9, -54, 88, -73, -22, -11, -9, -3, 55, -57, 93, 94, 11, -19, 13, 48, -12, 8, -52, 23, 66, -97, -92, -54, 68, -112, -54, 43, 18, -36, 127, 17, -57, -26, 72, -108, -105, 53, -119, -41, 111, -69, -26, 15, 39, -59, 35, -64, 45, 64, 65, -17, -124, 60, -66, -121, 76, 17, -113, 0, 92, -35, 45, -90, -67, 125, 41, -25, 8, -1, 95, -75, 14, -72, -58, 35, -58, 126, -127, -80, -12, -71, -19, 83, -98, 43, 95, -112, 37, -70, 58, 63, 7, -93, -124, -1, 26, -82, 51, -74, -111, 60, 49, -104, -76, 44, 92, -111, -97, -22, 19, -91, 120, -55, -93, 122, -66, -46, 38, 7, -5, 26, -120, -11, -37, -12, -94, 72, 64, -11, -126, 54, -6, 120, -24, -30, -41, -128, -91, -11, 113, 109, -50, -69, -57, -9, 92, 52, 80, 15, -75, 88, 5, 52, 0, 116, -79, 71, 6, -18, -21, 106, 122, -9, -66, -48, -96, -41, 103, -18, 70, -10, -67, -51, -93, -122, 11, 89, -61, 89, 100, 115, -117, 89, 3, -47, 8, 74, -65, 31, -81, -75, 100, 101, 127, 70, -40, -50, -116, 105, 37, -33, 16, -120, 120, 26, 100, -22, -11, 80, 57, 64, 69, -118, 48, 42, -79, 63, 1, 89, -3, 113, 56, -29, -25, 6, -89, -34, 0, 95, -11, 42, 106, -43, -27, -43, -73, 76, 82, 85, -28, -68, -128, 39, 9, 34, -112, -116, -46, -60, 46, 29, -11, 49, -10, -9, -116, -103, 46, 64, 91, -88, -57, -97, 114, -2, -72, 39, -103, 59, 32, -70, -6, -84, 58, 111, -116, 47, 125, -89, -70, -63, -35, -119, 67, 92, -56, -57, -1, 101, 92, 44, -67, 61, -7, 95, -87, -45, -92, -5, -73, 9, -61, 48, -16, 18, 95, -84, 70, -79, -128, -69, -37, 86, 28, -6, 18, 12, -87, 37, 57, -26, -107, 66, 17, 5, -60, -44, -50, 81, -104, 70, 8, 84, -62, 14, 74, -79, 71, -62, -21, -15, -48, 5, -108, -64, -47, 90, -114, 28, 34, -65, 100, -3, 34, -76, -98, 100, 27, -54, -13, -3, -29, -28, -57, 11, -3, -98, 100, 33, 85, 46, -47, -69, -34, 68, -22, -40, -123, -114, -108, 94, 124, -56, -8, 104, 79, 57, 42, 59, 0, -93, -29, -32, -16, 7, -19, 69, 36, 120, 111, -118, -103, 25, -21, 97, -50, -41, -26, -19, -27, 48, 93, 99, 61, -4, 9, 36, 81, -103, 90, -12, 105, -67, 104, -48, -57, -27, 48, 19, -104, -24, -13, 5, 40, 123, -8, -124, -113, -62, -101, 61, -26, 94, -31, -95, 1, 67, -128, 34, -114, -49, -116, -79, 26, 88, -75, 104, 61, -77, 105, 79, -69, 75, 81, 120, 42, -32, 81, -40, -110, -97, 27, 28, 42, 60, 127, -90, 66, -16, -6, -72, 64, -124, 33, 73, -95, -65, 43, 60, 26, -119, 6, -81, -88, -109, -72, 28, 84, 73, 88, -18, 38, -125, 115, -43, -83, -62, -42, 52, -115, -71, 69, -93, 60, -31, 96, -67, -122, -86, -79, -108, -37, -43, 20, -99, -80, 64, 104, -25, 53, 83, 29, -41, 24, 29, -107, 100, 13, 106, 49, 51, 4, -3, 95, -64, -55, -6, -65, -68, 80, 13, 37, 117, 53, 126, -31, 75, -108, 106, 114, -121, 55, 92, -31, -27, -29, 77, -109, 70, 80, -4, 48, -124, -101, 54, -9, 116, -22, 48, -124, -56, -109, -95, 120, -56, -82, -113, -94, -24, 72, 22, -87, 67, -10, -92, -59, 52, 81, -12, -111, 103, -67, 57, -125, -2, -120, 35, 2, 98, -85, -121, 0, -96, 108, -34, 28, 65, -110, 21, 56, 6, 75, 76, -62, -40, -117, -107, 16, -35, -113, -97, -62, -3, 82, -61, 111, 41, 9, -54, 79, 117, 77, -96, -53, -92, -27, -42, -110, 45, 120, 83, -35, -102, -81, 29, -115, 114, -98, -23, -16, -45, 53, -115, 7, 12, 12, -89, 13, 107, 32, 126, -83, 45, 66, 98, -119, 54, -65, -46, 40, 123, -112, -114, 73, 110, -128, -114, -112, -51, -108, -43, -37, -123, -110, 4, 26, 14, -109, 122, -35, -58, -73, 78, -116, 92, -84, -91, -6, -47, 80, -38, 90, 74, -76, -69, -114, 124, -87, -86, 62, -42, 73, 0, 97, -61, -43, -88, 63, -47, 52, -111, -38, 97, 49, 103, -109, -40, 65, 45, -2, -58, -98, -84, 104, 126, -94, -9, 28, 83, -87, 36, 82, 90, -40, 51, -112, 92, 84, 110, 16, -40, -81, -75, -70, -93, -92, -114, -72, -128, 106, -83, 92, -15, 56, 95, 37, -16, 0, 111, -82, 110, -2, -38, 11, -127, 103, -14, -21, -107, -100, -28, 63, -104, 117, 36, 20, -3, -72, 109, -70, -110, -63, -39, 35, -30, 16, -1, -128, 45, -89, 27, -73, -17, -16, 106, -43, -118, 3, -107, 2, 101, 62, 124, -15, 37, -22, 56, -24, 23, 27, -9, -123, 89, -64, 61, 46, 106, 124, -86, 3, 37, 2, 21, 62, -56, -37, 120, -65, 64, 22, -71, -51, -31, 12, -25, 109, -38, -100, 43, -116, -92, 24, -24, -102, 2, -94, -44, -7, -76, 97, -35, 63, 1, 97, 2, 96, 1, -98, 76, -63, -76, -48, 106, -11, 97, 95, 51, 101, -116, 120, 116, 99, -79, 43, -101, 61, 66, -101, -83, 69, 109, 18, -104, 17, -13, -6, 124, -110, -1, -87, 45, 83, -110, 97, -4, 98, 58, -35, 124, 49, 85, -35, -15, 3, 113, -106, 3, -32, 34, 64, -19, -45, 103, -15, 69, 51, -87, -43, 105, -126, -106, 61, 13, -17, 127, 109, -117, 61, 126, -59, 75, 14, -59, 67, -69, 28, -31, -71, -45, 63, -104, -59, 98, -73, -120, 106, -14, -27, -27, -87, 92, -51, 0, -12, 30, 99, 3, 111, -102, -34, -115, 106, 49, 89, 91, 109, 52, 97, 21, 41, 49, -103, -85, -105, -117, 27, -98, -109, -42, 33, -88, 113, 78, -12, -52, 76, -114, -18, -13, -76, -26, -127, 102, -28, -18, -71, 31, -26, 34, 82, -111, -121, -102, 19, 93, 32, -125, 23, 79, -70, -52, 68, 120, 99, -12, -99, -110, 80, 51, 118, -19, -120, 10, 59, -69, 75, -70, -110, -102, 122, -118, -127, -95, -95, 105, 72, -37, 67, -80, 86, -61, -120, 54, 106, 61, 50, 46, 16, 43, -81, 109, -65, 15, -62, -88, -32, 106, 2, -16, -2, 87, 97, -6, 69, -83, 50, 114, 105, 77, 55, -63, 111, 80, -66, 8, -73, 10, -95, -75, 94, -40, -6, -79, 14, 127, -105, -63, -68, -3, -65, 24, 121, -51, -11, -72, 20, 27, 51, 20, -80, 84, 15, -53, -35, 5, -122, -7, -72, -86, -121, -77, 13, 121, 55, -78, -85, -53, -48, 101, 5, -54, 55, -78, 109, -26, -56, 72, 85, 55, -125, 20, 48, -50, -10, -120, -27, 32, -41, -61, -14, -49, 39, -77, 93, 112, -87, 101, 88, -126, -52, -119, -27, 121, -92, 9, -120, -3, -111, 60, 113, 94, -48, 105, 12, 87, 76, -96, -105, 101, -2, -78, 94, 4, -97, -13, 16, 36, 11, 8, -112, -34, 37, 83, -49, -72, 72, -89, 20, -79, 34, -47, -14, -49, 79, -44, -32, -82, 112, 14, 57, -78, -43, -48, 118, -94, 18, -58, 7, 124, -65, -124, -107, -1, 0, -125, 127, -24, 123, -97, 45, -80, -118, 2, -36, 112, 47, 20, -47, 83, 0, -96, -120, -32, 99, -99, 82, -70, -47, -126, -108, -32, -19, -6, 74, 107, 38, 115, -84, -44, -33, 114, 30, 57, -34, -22, 84, -39, -90, -9, -78, -111, -39, -117, -21, -82, 111, -100, -111, -47, -107, -38, 68, 25, 13, -47, -9, 119, -63, 124, 21, 39, -98, -39, -85, 4, 100, 101, 38, -17, -17, -5, -83, 12, 29, 113, -91, -34, -65, -120, 0, -86, -17, 65, -86, 41, 17, -40, 79, -2, 68, 31, -85, -28, 106, -123, 100, 79, 110, 101, -29, 95, -122, 103, -126, 2, 109, 56, 75, -63, -7, 44, -112, 70, -66, 44, 47, 83, 26, -2, -36, -23, -52, 20, 7, 28, 56, -18, -59, -33, 69, 59, -111, -39, -22, -72, -31, -85, 108, 52, 25, -103, 74, 91, -83, 88, 126, -105, -69, 78, 7, 52, -32, 0, 106, 8, -20, 57, 82, -115, 65, -85, 126, 5, 68, -52, -38, -58, -17, 93, -11, 27, 110, 25, -19, -19, -109, 15, 95, 54, -121, 69, -6, -36, -117, -30, -71, 21, 36, 73, -52, -2, -122, -61, -99, 35, -90, 54, -92, 95, 51, 95, 108, -62, 108, 40, -118, -12, 116, -34, -98, -123, 110, 94, 93, -37, 30, 25, -93, 51, -29, -86, 114, -126, -19, 113, 72, -116, 85, 3, 97, -64, 49, -109, 72, -28, -38, -25, -44, -38, 92, 103, -56, 22, 24, -71, 109, 29, -35, 96, 97, -45, 70, 52, -75, -43, 51, 21, -59, -121, -10, -3, 6, 75, -128, -117, -27, -91, 3, -45, -122, 79, -104, 10, 84, -69, -36, -51, 65, -58, -119, 27, 60, -5, 88, 89, -102, -33, 103, 11, -63, -118, -37, -90, 18, 84, -9, 101, 77, -95, 9, -77, -128, 23, 58, 49, 48, -3, -79, -50, 81, -57, 100, 58, -73, 80, 127, 94, 47, -46, -106, 71, 11, -76, -2, 94, -44, -2, -32, 63, -128, -36, 125, -104, 107, 97, 18, -60, 59, 94, -20, -119, 16, 116, 106, 117, 49, 90, 102, 54, 18, -32, 123, -92, 54, 111, -126, -28, -93, -88, -27, 10, -111, 41, 74, -19, 67, -108, 111, 96, -89, 108, 103, -86, -58, 59, 61, 102, 24, 55, 75, -16, -55, -108, -4, -58, -65, -109, 122, -64, -29, -73, 119, -110, -55, 92, 84, -111, 24, 96, 10, 45, 10, 69, 4, -80, 5, 95, 114, -79, 21, 21, 63, 47, 39, -83, 110, 84, 92, 32, 51, -68, 75, -36, -4, 71, -77, -9, -109, 85, 103, -58, -57, 123, -85, 41, -98, -106, -58, 2, -81, 50, -86, 107, -67, -60, 71, -18, -113, -66, -68, -37, 36, -81, -28, 16, -1, -53, 70, -41, 98, 114, -36, -88, -56, 16, -76, 104, -36, -125, 25, 61, -113, -62, -75, -112, 99, -24, -29, -53, 100, 124, 27, -24, 16, -121, 87, 28, -21, -5, -15, 23, -81, -101, -25, 106, -23, 59, 47, 2, -100, -6, 11, 118, -105, -45, 65, 65, -123, -110, 6, -7, -78, 86, -119, 89, 106, 2, 55, 79, -117, -52, -50, 109, 102, -5, -70, 37, 56, 49, -78, 110, 71, -104, -22, 113, 110, 18, 113, -13, -119, 29, 4, -4, 47, 108, -113, -90, 35, 116, -75, -105, -117, 62, -24, 76, 5, 98, -44, 33, 121, 80, 77, -82, -85, 91, -65, 63, 80, -4, -35, 94, -94, -35, 88, 27, -28, 120, -81, -57, 67, -12, 45, 52, -90, 117, -127, -103, 96, 62, 114, -124, 124, 69, -22, -11, 44, 40, 22, -128, -63, 20, 24, -112, -10, -65, -92, -50, -36, 93, 22, -94, -53, -62, 90, 78, -112, -64, 103, 16, -29, 26, 58, 14, -76, -56, -49, 16, -102, 6, -97, 39, 2, -60, -120, 76, 20, 62, 127, 97, 5, 106, -106, -116, 112, -45, 76, 83, 107, 81, 7, -42, 2, 98, 48, 103, 2, 104, 0, -89, 38, -100, -10, 43, -107, 40, 118, -10, 71, -7, -116, -28, -103, -62, -114, 8, 121, 108, -17, -70, 48, 45, 51, -115, 30, -71, -102, -28, -115, -76, 20, 92, -90, 4, -105, -68, -19, -91, -51, -31, -98, -2, -85, 75, 93, 90, 114, 113, -104, 115, -58, -14, -63, -7, -88, 93, 15, -80, -116, 3, 124, -17, 100, 126, -83, -16, 31, -41, 103, 36, 71, -25, -43, -54, -26, 2, -124, 65, -45, 77, -67, 66, -10, 18, 11, 116, 106, -76, -94, -4, 95, 61, -118, -92, -22, -3, 79, 9, 29, 116, -26, -29, -41, -40, 46, 43, -73, -98, 109, -89, 112, -98, 7, 48, -18, 97, -117, 62, 81, -75, -72, -116, -77, -22, -66, -59, 113, 1, 44, -8, -98, -72, 126, 27, -26, 72, 41, 124, -11, -127, -35, -119, -32, -95, 35, 44, -50, 52, -2, -32, -26, 42, 79, -100, -106, 29, 81, -108, 76, -84, -105, -6, 32, -83, -108, 99, -37, 65, 102, 91, -70, 70, -48, -65, 33, 41, 80, -7, -94, -125, -116, -21, -107, -99, -117, -67, 117, -92, -100, 16, -58, 127, -67, -120, 89, 74, -108, -74, -80, -23, -90, 50, -81, -115, 86, 32, -22, -43, -80, -103, -82, 3, -87, -87, -63, 5, 21, -112, 98, 64, -95, 125, -60, -2, -11, -32, -108, -14, 96, -44, 40, 60, -61, -48, -39, 39, 5, -20, 5, 111, -14, 85, 28, -116, 106, -77, 63, -29, -94, -47, -77, -106, 107, 103, 60, -118, 16, 55, -2, -20, 34, -82, -108, 77, 37, -73, 71, -95, -51, 42, -112, 116, 56, -60, -113, -111, 94, -18, -125, 4, 74, -33, -90, 113, 95, -43, -96, 55, -11, -7, -27, 123, -5, -104, 14, -6, -100, -34, 2, 102, -36, 108, 32, -2, -76, -51, -22, 16, 51, 73, -118, 65, 124, -51, 91, 48, 127, -1, 79, -2, -56, 2, -22, 45, 104, 19, -26, 46, -1, -109, 45, 5, -17, 32, -81, 106, -91, -25, -122, -76, 38, -22, -27, 25, -27, -40, -44, 46, -102, -1, 84, -43, -126, 48, 62, -53, 64, -50, 121, 2, 111, -47, -126, 93, -20, -98, -63, -96, -9, -126, 88, -3, 81, -120, 116, 117, -52, 24, 9, 98, 84, 54, 122, 8, 94, 92, 25, -46, 49, -80, -42, -89, 80, -69, -10, -114, -119, 14, 80, 63, 55, -19, -107, -114, 36, 43, -9, -127, -82, -83, 104, -62, 52, 119, 4, -113, -118, -59, 52, 13, 0, -93, 62, 33, -101, -79, 50, 122, 61, 126, -85, 92, 114, 98, 42, -124, -93, -121, -125, -110, 17, -108, 108, -42, -63, 38, 35, 31, 64, 71, 122, 82, 88, -12, 72, 122, -47, 69, -53, 95, -91, -96, -55, 126, 79, 85, 8, 12, -39, 54, 49, -67, 94, -114, 37, -104, -81, -60, -70, 122, -74, 53, -19, -118, 90, 40, 74, -69, -1, 84, 80, 86, -88, 100, -108, 100, 45, -43, 16, -11, 26, -106, -48, 7, -19, -77, -49, 100, -21, -113, -115, 94, 90, 7, -24, -60, 85, -80, -71, -27, 57, 51, -76, -121, -12, 36, -111, 1, -77, 53, -28, 121, -93, 0, 92, 54, -61, -34, 98, 56, 49, -21, 36, -41, -37, 42, 125, -84, 62, 127, -18, -32, -106, -102, 7, -70, -83, 127, -19, -102, 118, -39, -86, -55, -12, 43, 68, -108, 58, 104, -76, 85, -100, -5, 45, 47, -24, 98, 85, -90, 96, 95, 123, -85, 106, 110, 54, -101, 99, 28, 61, -44, 71, -60, 62, -27, -92, -32, -31, 90, -53, -26, 30, 2, -67, -90, -63, 20, 12, 59, 45, 84, -18, 46, -103, -73, 95, -29, -47, 55, 93, -31, -56, -116, 7, 102, -19, -75, 15, -7, -65, -37, 36, -103, 88, 26, -113, -33, -116, 116, -83, 9, -4, 31, 75, -32, 37, 5, -63, 52, -100, -50, -77, 107, 87, -20, -127, 36, 105, 69, -128, 127, 88, -126, 33, -28, 78, -64, -15, -8, 58, -15, 120, -3, -123, 19, 5, 43, -6, -122, -28, 37, -66, 73, 70, -4, -105, -91, -119, -43, 127, -67, -44, 82, -19, -6, -75, -123, 16, -75, 58, 29, 97, 29, 117, 27, 56, 87, 37, -31, -57, -109, -33, 119, -21, -96, 109, -89, 3, 74, -110, -79, 20, 23, 71, 9, 125, -98, 0, -18, -16, 123, -57, 60, 127, 11, -26, 76, -36, -74, -8, 21, 14, -45, -77, 55, 0, -57, -44, -44, 106, -57, -66, -17, 28, -89, 98, 6, 103, -4, 106, 88, -14, 35, -42, -35, -109, 89, 88, 30, -102, 65, 127, -109, -108, -119, -93, -99, -85, 96, -30, -121, 20, -10, -101, -25, -58, -105, -41, -42, 118, -73, 75, 74, 69, 116, 127, -28, -52, -48, -33, 53, -3, 109, -45, -23, -7, 27, 74, 120, -107, 22, 30, -112, 33, -84, 75, 72, -33, -52, 60, -87, 98, 49, 21, 120, 48, -13, -83, -125, -32, -12, -126, 3, 108, 19, -41, 87, 22, 52, 122, -91, -105, 48, -55, 104, 7, -90, -59, -11, 79, -8, 16, 95, -58, 67, 91, 56, -122, -43, -62, -7, 50, -112, -117, 8, -118, -98, -98, 51, -109, -20, 30, 13, -104, 116, -26, -57, -95, -76, 67, 32, -39, -56, 90, 33, -39, -9, 70, 81, 93, 112, -52, -19, -6, 37, 109, -54, -116, 43, 73, -70, 90, 101, 125, 3, 34, -25, -82, 30, -108, 20, -15, -60, -118, -119, 121, -87, -78, -38, -41, -70, 63, -80, 34, -16, 114, -89, -120, 68, -112, -39, 14, -56, 118, -13, -9, 96, 12, -38, -63, -54, -58, -32, 60, 36, 54, 32, 106, -122, -89, 83, -103, -26, -87, -114, 77, -51, 3, 33, -64, 110, -11, -29, -115, 71, 71, -39, -64, -7, 123, -30, 12, 59, 28, -21, 54, 44, -102, -122, 12, 4, -114, -23, 17, -114, -86, 34, -61, 38, 47, 116, -34, -127, -64, -23, 20, 110, 78, 10, 35, 74, 70, -24, 44, 46, -100, -15, -119, -33, -85, 7, 5, 55, 100, -12, -47, -47, 122, 1, -15, 110, 18, 8, -86, 75, -4, 78, 27, -106, 104, -71, 111, 73, 59, 69, -120, -24, -16, 13, 80, 72, 93, 124, 6, -100, 94, 80, -12, -95, -86, 65, 49, -126, -76, 94, 110, -34, 34, 8, 92, -88, 102, -95, 124, 86, 104, 80, -82, -91, 90, 87, -80, 58, 40, 19, -123, 84, 94, -50, 14, 7, 111, 61, -100, 63, -36, -28, 109, -116, -63, 39, -57, 44, 79, -11, 40, 113, 109, 40, 75, 84, -42, 72, 66, -61, 47, -61, -48, 48, 104, -77, -101, -10, -62, 89, 29, -37, -117, 31, -102, 111, 0, 44, -32, -26, -32, -114, -55, -109, 116, -72, 6, 11, -76, 11, 69, -99, 110, 58, 59, 88, -32, -71, -115, 41, 55, -31, 81, 35, 79, 36, 78, 4, -29, -8, -98, 111, -118, 60, -10, -81, -11, 27, 99, 55, 50, 71, 120, -10, 28, -77, -72, -68, 59, 119, -54, 127, -63, -56, -120, -70, 62, -58, 14, -115, -37, 22, -119, 90, -105, -73, 4, 80, -59, 38, -92, 13, 16, -24, -66, 39, 122, -80, 122, -66, -64, -14, -67, 98, -84, -55, 21, 40, 5, 22, -30, 69, -57, 52, -66, -68, 4, 22, -93, 127, 103, -22, 46, 11, 81, -43, -57, 114, 77, 60, -102, 65, -71, 118, -85, -97, -4, 57, -109, -109, 21, -97, -43, -7, 121, -82, -112, -41, 79, -56, 127, -105, -25, 92, -34, -107, 96, -77, 68, -44, 34, -102, -111, -96, 103, -2, -94, 70, -54, 55, 36, 40, -78, 121, -30, -104, -6, 35, 72, 87, -37, 103, 30, 48, 41, -80, -84, -69, 42, -108, 14, 10, -113, 104, 91, 7, 65, 15, 3, 27, 3, -97, -9, 113, -86, -19, 11, 74, -43, 119, 110, -54, -94, 82, 15, -110, -81, -78, -127, -51, -49, 121, -109, 9, -73, -100, -85, -121, -91, -125, -15, 125, 67, 127, 27, -61, -44, -75, 63, 58, -54, 76, 23, 102, 95, 36, 53, 83, 62, -13, 71, -76, 8, -89, 102, -34, 105, 42, -80, 24, 123, 76, 44, -3, -103, -70, -44, 12, -94, -55, -14, 9, -77, -52, -4, -48, -83, 7, -22, -124, -60, -67, -63, 18, 36, -92, -96, -56, -128, -35, -88, 71, -68, 117, 2, 126, -42, -63, -111, 96, 42, -11, 64, 84, -2, 36, 12, -41, 41, 117, 101, 29, -38, 8, 105, 88, -115, -78, -86, -128, 74, 18, -16, -12, 9, 78, 113, 88, -84, 60, 50, 46, -122, 79, -107, 122, 13, -54, -56, 28, 21, 57, -32, 111, 83, -122, 91, -80, 60, 40, -109, 111, 64, 119, 8, -85, -10, 36, 99, 6, -56, 12, -92, -111, 61, -76, 33, 93, 70, 114, -4, -53, 68, -41, -38, 15, 81, 5, -61, 120, 28, -119, -35, 54, -98, 109, -117, 19, -55, -123, -43, 29, -3, -69, -1, 39, -110, -7, 13, -15, -38, 56, 103, 62, 39, -51, -87, 122, 33, -92, -113, 77, 114, 90, -67, 115, -22, 66, 37, 88, 124, 73, 79, -51, 96, 93, 76, 120, -16, -112, -77, -107, -81, 83, -57, -62, 78, -124, 8, 25, 117, 44, 31, -1, -7, 25, -53, -57, 27, 95, 66, 38, 9, -121, 35, 104, -44, -11, -23, 11, 56, -111, -123, -52, 127, -49, 14, 44, 12, -108, 58, -54, -42, 70, 51, 0, 101, -85, 10, -16, -52, 90, 59, 64, -29, 66, -117, 72, -22, 79, 19, 3, -52, -41, 51, 82, 38, -60, 33, 54, -104, 87, 126, 11, 75, -46, -64, -9, 57, -122, -92, 86, -77, 42, -46, 4, 10, -13, 90, -59, -117, -34, 96, -63, 122, -19, -26, 56, 95, 42, 105, 91, -69, 88, -62, 108, 13, 118, -49, 21, -21, -106, -96, -64, 126, -3, 55, -87, -67, 94, 33, -128, 2, -56, -48, -11, -114, 15, 21, -20, -38, 55, -80, 9, 7, 88, -76, 45, 40, -128, -102, 89, -95, 72, 122, -91, -125, 28, -59, -114, -69, 14, -15, 116, 13, 10, -63, -109, -11, 33, 3, -43, 20, -90, -65, -69, -91, -87, 24, 42, -69, -3, -121, 55, -12, 102, 93, -68, -40, -75, 58, -4, 27, -55, -10, -69, 73, -97, -110, 13, -25, 92, -34, 123, -52, -41, 83, 14, -35, -121, 34, 43, -72, 73, -54, 86, -100, -83, 115, 125, 123, -74, -9, -109, 16, 117, -62, -82, 94, 103, -20, 83, 50, 124, -22, -83, 33, -37, 28, 36, -69, 62, 99, 12, 89, -26, 113, 4, -111, 127, -95, -71, 44, 40, -113, -108, -65, 46, 36, -70, 77, -59, 113, 106, 32, 102, -80, -77, -92, 32, 121, 37, 78, -100, 117, 19, 87, 67, -29, -26, 53, -82, 0, -41, 120, 96, 47, -38, -83, -62, 68, -33, 50, 87, 106, -102, 34, 21, -103, 117, -17, -73, 71, 17, -34, -92, -30, -102, -100, 70, -127, 70, 110, 57, -22, 72, 56, 42, -47, -14, -69, 110, -71, 74, 22, -99, -121, -127, 17, -80, 3, -94, 112, 90, 53, -9, -16, 118, 56, 34, -86, -105, 29, 113, 29, -6, 44, -5, -53, -98, 1, -59, 25, -110, -48, 127, -101, -96, 99, 19, -24, 81, 82, -97, 32, -110, -16, 56, 2, 24, -55, 40, -116, -125, -99, 60, 121, 94, 106, -91, 70, 50, 53, 36, -101, 52, -16, -57, 127, -44, 56, -36, -42, -119, 48, -113, 34, 108, 78, 2, 94, 68, -118, -108, 30, -66, -38, 15, 100, 125, -16, -119, 15, 4, -109, 15, 24, -12, 86, 90, -98, 15, 84, 62, 23, 60, -16, -93, -29, -98, 67, -98, -110, 103, -121, -67, 113, 69, 123, -123, -77, 42, -94, 63, -112, -119, 80, -93, 45, 0, 68, -44, -28, 61, -109, -83, -107, 38, 54, 104, -92, 97, 21, -66, 37, 39, -89, 87, -42, -75, 59, 18, -102, 40, -8, -25, -42, 110, 103, 40, -97, 64, -71, 124, 125, -107, -83, 54, -105, -1, -69, -35, 22, -37, 102, 76, 49, 50, -107, 29, -57, 123, 122, 4, 9, 65, 80, 39, -84, 118, -40, 81, 47, -66, 66, -80, 65, 121, -1, -18, 127, -99, -12, -99, -24, -110, 126, 43, 26, 114, 74, -5, -100, 14, -80, -90, -5, -80, -86, -53, -82, 93, -35, -67, -64, 77, -95, 127, -12, 31, -107, 49, -44, -82, 48, 86, 102, 92, 36, 85, -62, -104, -91, -28, 89, -100, 78, 102, 100, -122, 53, 34, 24, 28, -53, 104, 44, 121, -13, -99, -101, 90, 118, 63, -75, 93, -40, 81, 17, 114, -5, 62, 36, -28, 46, 18, 20, 41, -76, -3, 40, -88, 44, -70, -80, -5, 0, -116, -112, -28, -121, 84, -116, 36, -10, 69, 111, 27, 1, 8, 89, -121, 30, 43, 59, 54, 84, -74, -105, -94, -48, -30, 91, 49, 65, 49, 86, -102, 103, 47, -92, 41, -100, 106, 49, 126, -27, -114, -101, -91, -98, -81, -121, -64, 66, 34, -65, -71, 63, 70, -73, -82, 126, -32, 28, -37, -122, 25, -56, 29, 40, 29, 99, 30, -53, 18, 97, 49, 27, 77, -109, -120, 70, 49, -37, 104, 40, -26, 125, -110, 56, -100, -76, 53, -2, 127, -63, 79, 14, -47, 111, -95, -41, 43, 59, -20, 33, -104, -38, 115, 69, -23, 12, 41, 39, -30, 76, 44, 44, 101, 120, 53, 57, 53, 24, -23, 64, 72, -17, -102, 25, -112, -23, 34, 53, -35, -17, -101, 48, 21, -51, 103, 89, 1, -34, 87, 50, 99, 23, 7, -29, -114, 12, 61, 126, -11, 81, -99, 44, 48, 62, -126, -12, -53, -59, 49, 35, -112, -114, 111, 30, -12, 77, -90, 0, 18, 78, -84, -44, -44, -63, 59, -56, -17, -84, 53, 50, 125, 56, -47, -107, -115, -73, 9, 65, 0, -91, 38, -58, -50, 25, -31, 73, -60, -4, 11, 49, -30, 93, -27, 61, 31, -13, -75, -94, -77, 25, -95, -113, -122, 14, 38, -92, 9, 79, -1, 21, 98, -4, 91, -2, 45, 57, -14, 23, -54, -125, 111, 124, -51, -61, -10, -47, -64, -74, -24, 127, -5, 113, -37, 33, 0, 24, -62, -71, -109, 95, -32, -92, -53, -15, -32, -37, -28, 74, 84, -23, 51, 70, -128, -74, -37, 83, 29, 82, 74, 53, -99, 62, 52, -112, 56, 110, -117, 124, 108, 10, -114, -28, -118, -91, -61, 7, 114, 75, -44, -1, 5, -115, 37, 84, -6, 62, 63, -26, 7, 115, 54, 60, -103, -113, -42, 109, -93, 82, 69, 72, -121, 85, 95, -88, 94, -31, -42, 74, 65, -66, -70, -80, 43, -126, 46, 110, 16, 14, 97, -114, 9, -49, -34, 113, 101, -107, -52, -101, 109, 53, -111, -29, -1, 27, -78, 55, -82, -50, 116, -109, -62, -92, -126, 113, 79, 6, 26, -35, 100, 4, -13, -1, 7, -43, -89, -64, 42, -64, -116, 100, 41, -33, 57, 47, 91, -18, -113, -85, 114, 27, -64, -91, -63, 54, 122, -84, -96, 62, 115, 113, -119, -61, 76, -116, -88, -98, 117, -56, -121, 75, 84, -78, -127, 35, -65, 108, -89, -27, 23, -9, -3, -34, 69, -114, 104, -7, -103, 120, 24, 114, -96, -49, 90, 50, -100, -97, 97, -11, 123, 8, -60, -54, -78, 13, 69, 67, 29, -89, -87, -94, 37, 23, -18, -14, -73, -6, 34, -91, 107, -58, 105, -22, 67, -117, 67, 105, -44, -125, -29, -102, -48, -4, -91, -117, -26, -62, 13, 43, -58, 65, 39, -30, 122, 62, -123, 23, -4, -75, 67, -64, 117, 103, -31, 82, 80, 116, -19, 13, 21, 104, 126, -3, 125, 47, -116, -41, -83, 68, -98, -35, -31, -127, -51, -21, 49, 80, 75, 101, 22, 102, -16, 57, 46, -92, -48, 86, -108, 98, 5, -28, 79, 115, -94, -97, 103, -56, 117, -92, 10, 82, -104, 2, -21, -43, -37, -124, 126, 124, 23, -97, 53, -31, -106, 95, 123, 90, 3, 122, -90, 45, 22, 48, -128, -113, 70, -85, -74, 37, 79, -119, -39, 5, -120, 24, 55, 90, -70, -46, 35, 83, 83, 20, 61, 101, -85, 4, 51, 57, 88, 126, -84, 125, 117, 11, 62, -17, 13, 73, -105, 114, 78, -117, -11, 107, 79, 88, -9, 40, -99, -78, 106, 80, -53, 66, -116, 41, -58, 5, 67, -77, -60, -55, -22, -32, 99, -61, -116, 113, -71, -98, 76, -98, 94, 116, 31, -32, 58, -120, -1, -83, -44, 80, 110, -126, 39, -126, -45, -4, 33, 77, 62, -35, 17, 90, -9, -126, 124, -50, -12, -29, 57, 63, 101, -70, 83, -68, -86, -113, 66, 99, 7, 35, 111, 123, 107, 56, 124, -83, 97, -64, -38, -61, -111, -53, 104, -83, 67, 108, 53, -45, -113, -26, 121, 36, -122, 25, -68, 22, 121, 54, 20, -57, -69, -23, -103, 127, -7, -6, 103, -61, -9, 82, -74, -45, -126, 5, 74, -118, 14, 11, 65, 96, 90, -103, -7, -14, 114, 71, -45, -101, -7, 56, 2, -86, -86, -109, 90, 19, -63, 90, 61, -106, -60, 47, 43, -105, -8, -1, -127, -116, 3, -92, 82, -47, 0, 27, -63, -81, -19, -89, -10, 120, 45, -54, 73, 95, 125, -84, 15, -47, -34, -36, -57, 35, 8, -16, 119, 122, 61, 59, -111, -113, 45, 97, 40, -119, 90, 14, -84, -43, -19, 21, -98, -67, -120, -38, -41, 44, 6, -10, 113, -49, -53, 49, -16, 10, 38, 120, 8, -115, -51, 34, 124, -73, 115, 18, -31, 12, 73, -84, 13, -102, 9, 68, -99, -60, 74, -47, -97, 56, 75, 64, -87, 64, -1, 91, -121, 40, 14, -8, -49, 116, 17, -10, -73, -34, 16, -23, 45, -113, -128, 37, -108, -112, -53, 68, 126, 22, -63, -16, -103, 127, 45, -66, 35, -120, -83, 3, 23, 69, -38, -77, 94, 121, 109, -94, -12, -99, -73, 80, -49, 37, -77, 12, 103, -28, -121, -18, 41, 126, -116, -103, -119, 46, -93, 24, 123, -42, 113, 122, 68, 11, -101, 25, -111, 79, -2, 72, -27, -117, -49, 60, -5, -28, -107, 96, -16, 65, -48, 8, -31, 71, 56, -54, -20, -47, -112, -119, 2, -35, 110, -45, -110, 25, -121, 95, 76, -3, 72, -14, 38, -36, -116, 60, 46, -50, 106, -115, -45, -28, -70, 44, 61, 126, 33, 92, 98, 85, 55, 103, -11, -86, -27, -104, -20, 109, 42, 98, -17, -24, -38, -117, -119, -84, 14, 102, 42, 16, 63, -88, -119, 19, -10, 102, 20, 117, 28, -51, -94, -34, -122, 88, -80, 124, 118, -70, 108, 111, -112, -18, 80, 3, 117, -115, 43, -109, -17, -56, -43, -25, -80, -101, -27, -38, -66, -19, 125, 46, -121, 15, -109, -120, -97, 106, -4, 54, -21, -25, -65, -110, 119, -3, 23, -97, 24, -75, -123, -56, 8, 123, -104, 105, -50, -62, 25, -128, -106, 85, 42, 101, -75, -99, -14, -94, -100, -3, -10, -67, 43, 90, -93, -45, -55, -32, -97, -57, 33, 122, -60, -60, -99, 12, 106, 13, -116, 24, -55, 6, 80, -84, -93, -73, -61, -36, -75, 12, -72, -39, -44, -32, 3, -93, 107, 64, -59, -95, 21, 41, 125, -11, 17, -4, 63, -124, 118, 60, -70, 97, 18, 123, -15, -124, -23, 54, -114, -83, 95, -121, -30, 41, -83, 82, -86, -24, -124, -18, -95, 120, -28, 12, 66, 106, 78, -48, -98, 53, -50, 41, -105, -112, -101, 118, -95, 89, 24, 117, -125, 49, -99, -11, 40, 28, -116, 114, 96, -118, 2, 15, -6, -61, 77, 101, 26, -72, 26, -109, -91, 86, 64, 58, 22, 13, 77, 125, 72, 42, -6, -107, -71, -112, -128, -76, -84, 33, 0, 29, -59, -80, -78, 109, 3, -79, 121, 14, 46, 53, 13, 100, 33, -112, 94, -95, 64, 61, -38, 31, 58, -10, -69, 18, -121, -128, 102, 36, -75, 36, 55, -95, 103, -87, 58, 75, -97, 124, -128, -74, -52, -14, -100, -12, -64, -17, -82, -91, -24, -10, 114, -83, -70, 19, -66, -63, -35, -11, 114, 75, 70, 16, 15, 77, -33, -47, 104, 82, -11, 107, -80, 73, -69, -31, -25, 102, 85, 64, 126, 0, -20, -46, 52, 33, -58, -4, -95, -97, -25, -34, 43, -72, 99, 82, 68, 67, -8, 33, -117, 71, -63, -29, 2, -45, 11, -104, 65, 101, 76, -41, 94, -109, 67, -32, 79, -118, -128, 81, 86, 11, -124, 3, 109, -59, -52, -31, 81, -9, 107, -4, 123, -42, 58, 127, -117, -52, -20, 3, -78, 84, -123, 31, 47, -29, 89, -128, -65, -114, 93, 122, -54, -86, -18, -34, -6, -10, -47, -11, 97, 106, 126, 88, -124, 10, 53, -100, -4, 64, -54, 119, 46, 23, 27, -127, 1, -43, 51, 26, 113, -92, -22, -125, 100, -17, 93, -107, 75, -25, 125, 112, -119, 122, 21, -15, -55, 24, 113, -32, 86, -45, -99, 73, -78, 80, -100, 112, -84, -51, 2, 0, 69, -98, 86, -112, -95, 1, 124, -117, -70, -55, 116, -51, -74, -49, -1, -86, 95, -51, -13, -106, -112, 109, 51, -75, 104, 40, 86, 88, 72, 30, -40, 123, -40, 7, 110, -44, -83, -94, 64, 43, 39, -22, -59, -61, -73, 115, -10, 81, 29, -47, -54, 59, -119, -99, -4, 20, 59, 11, -95, -52, 126, -81, -12, -123, 33, -57, 123, -64, 3, 108, -22, -88, -99, -51, 59, -125, -117, -87, -92, 58, -32, 55, -47, 95, -59, -35, 33, 6, 98, -30, -72, 24, 76, 70, 108, 34, -61, 5, 68, -5, 42, 114, 84, 119, 5, 75, 107, -76, -74, 14, 25, 33, 14, -66, -48, -42, 19, 104, 49, -100, -105, -96, 112, 95, 62, -76, 31, 70, 47, -102, -67, 36, 115, -64, 38, 5, -14, -19, 7, -43, -33, 119, 117, -105, 119, -95, -38, -3, -28, -92, 125, 50, -17, 111, 118, -68, 32, 18, 20, -89, 70, -17, 89, -84, 97, -23, -18, -92, 69, 78, -67, 52, 69, 93, -14, 6, -1, 2, -105, -53, 60, -110, -41, 73, 26, 45, -123, 116, 59, -34, 105, -24, 94, -11, 71, 17, -112, -84, -5, -24, 9, 82, 58, 114, -102, -44, 56, 41, 23, 107, -92, -37, -109, -58, -125, -71, -67, 90, -47, -61, 71, 1, 101, 22, -7, 118, 64, -82, -5, 14, -83, 53, -60, -11, 85, 52, 33, -20, 52, -115, 15, 96, 63, -20, 121, -62, 54, 26, 115, 36, 126, -96, 101, -86, -46, 90, 32, -16, -84, -111, -29, -44, 24, 48, -87, -60, -102, 91, -123, -46, 59, 10, -100, 55, -120, -117, -4, -37, -18, 73, 22, 3, 4, -70, -76, 65, -47, 23, 54, 82, 107, 115, -77, -112, -81, -122, 10, 33, -54, 99, -6, 74, 0, 55, 91, -52, 12, -118, -4, -25, 61, 80, 25, 12, 68, 53, -24, 46, 65, 14, 41, 40, -27, 64, 96, -14, -83, -46, -71, -66, -69, -69, 120, -4, -57, -124, 84, 17, 17, -6, -25, 43, -9, 60, 97, 30, -22, -89, 72, -122, 58, -120, -100, -97, 74, -46, -52, 43, -62, -28, -72, -118, 61, 7, -76, 103, -25, 56, -9, -31, 65, -92, -106, -67, 95, 116, -93, -70, -39, -81, 106, -29, 78, 96, 82, 13, 127, 7, -69, 110, -65, 80, -11, -109, 33, 70, -119, -117, 114, 35, 55, 31, 30, 108, 11, 12, -108, 119, -89, 38, 75, 117, 52, 98, 48, 121, -107, -125, -1, 86, 33, 20, 9, 17, 113, 13, 98, 121, 34, -9, -114, 30, 11, -61, -30, -31, 61, -22, 93, -116, -122, 29, -108, 90, -68, 91, -120, 1, 101, 108, -108, -43, 26, -65, 69, 120, -124, -90, -86, 53, 85, -96, 123, 26, 101, -28, -107, 7, 98, 29, 27, 107, 25, -49, -46, 121, -7, 51, 35, -28, 66, 99, 119, -59, 4, 85, 113, -101, 27, 104, 68, -71, -93, 122, -98, 38, -39, 51, 107, 116, 24, -23, -1, 106, -3, 77, -31, 40, 38, 47, -123, -120, 33, -86, -29, -39, -94, 109, 74, -97, 64, -16, 66, 124, -57, 110, -79, 48, -40, 37, -32, -85, 5, 117, -37, 40, -11, 11, 115, 77, 8, -45, 52, 98, -58, -83, 86, -29, 46, 82, -86, -29, -122, -110, 15, -40, -3, -126, 126, 108, -20, -100, 44, 29, -22, 87, -88, -35, 34, 14, 118, 11, -68, 28, 82, 65, -12, 110, 0, -56, 103, 107, 59, 7, 17, -42, 23, -84, -38, -94, 96, 56, 114, 126, -1, -73, 3, -108, 80, -11, -85, 31, -122, 103, 87, -19, 75, -48, -48, -56, 38, 123, 102, -86, -48, 79, -9, 85, 47, 63, -6, 127, 113, 8, -87, 87, -67, -89, -120, 115, -106, -122, 7, 112, -119, -22, 113, 122, 18, 91, 94, -121, 116, 92, 34, -126, -22, -78, -89, 7, 84, -98, -30, -120, -112, -124, -31, 85, 17, -38, 63, -48, 121, 0, -13, 25, -128, 125, 2, -84, -58, 52, -10, -20, 44, 68, 22, -67, 53, -68, -11, 25, -65, -19, -101, -32, 99, -111, 79, -6, -97, 85, 125, -127, -20, -122, 62, 91, -67, -104, 108, 56, -81, 48, -23, -72, 63, 99, 104, -122, 13, -39, 71, 79, 1, 86, -73, 52, -21, 41, -28, 109, 51, -16, -94, 44, 65, -34, 106, 12, -109, -37, 68, -103, 59, -65, 33, 39, -35, 1, 14, -111, -121, 80, -83, -96, -71, 68, -115, 104, 9, -3, -39, 24, 80, 75, 23, -18, 51, 12, 75, -89, -87, 39, 82, 9, 67, 112, 110, -116, 34, -33, 54, -79, 48, -103, -25, -75, 104, 93, 9, -23, -112, 31, -41, 56, -118, -83, 124, -97, -52, -66, -44, 6, 62, -44, -24, -62, 83, -10, -53, -66, -42, -29, -84, -120, 121, -49, 100, 49, 122, 55, 106, 54, -21, 115, -18, 17, 114, 50, -33, -63, 110, 25, 42, -93, 17, 113, 61, -118, -9, 123, -109, -23, -111, 65, -122, -14, -29, 69, -8, -22, 2, -88, -70, -86, 116, 18, 58, -86, 20, -86, -12, 62, 32, 57, 0, -25, 106, 103, 95, -25, 31, -78, 7, -13, -92, -33, 38, 57, -16, -40, -106, 34, -22, 55, 57, 113, -122, 34, -32, 86, 26, 30, 78, 109, 84, -80, -67, -111, -122, -2, -85, 98, 59, -106, 22, 18, -97, 75, -16, 23, -110, -90, -13, 10, 41, 14, -24, 65, -69, -4, 20, -29, 32, -81, 13, -50, -22, -83, 72, 78, -13, 67, 121, -77, 115, -7, -96, -25, -34, -10, -76, -16, 61, -99, -15, 103, 41, -46, -64, -41, 82, 20, -88, 100, 53, -32, -112, -123, 95, -47, -95, -45, 54, 2, -69, 44, -33, -124, -73, 32, -49, -77, 51, -104, 96, 119, -99, -18, -104, 67, -119, -125, -69, -9, -120, 120, -119, 67, 122, -109, 73, -51, -40, 76, 98, 51, -78, -51, 49, -77, 106, 19, 103, 31, 100, 85, 82, 114, 103, 59, -34, 127, -30, 22, 47, -97, -116, -108, -106, 74, -92, -126, 71, 118, 99, -82, -65, 31, 79, -94, 80, 18, 106, -23, 74, 125, -14, 117, 33, 49, 122, -110, 52, 34, -64, -101, -40, -91, -32, 43, -105, -9, -57, 41, 71, -85, -31, 8, 51, -103, -11, 116, 56, 38, 9, -87, 17, -30, 93, 65, -73, -78, 61, -43, 89, -96, -102, 11, -98, 22, -80, -10, -78, -126, -37, 59, 44, 62, -14, -55, -97, 122, 13, 111, -19, 41, 87, 115, -50, 24, -66, -17, 5, 80, -31, -46, -2, -51, -17, -123, 81, -125, 127, -14, -37, 18, -3, 27, 70, -45, -10, -52, 22, -4, -62, 123, 84, -35, -3, 2, -17, -62, 110, -101, -115, -32, 119, 33, -14, -128, -4, 1, 71, -52, -31, -32, 86, -9, -94, 38, 34, 79, -98, 4, -108, 20, 71, 23, 69, 60, -12, 37, 98, 52, 52, 87, 77, 106, -96, -72, -93, 124, 114, -56, -86, -88, -70, -2, -67, -23, 50, 4, 74, 53, -123, 11, -100, -103, 60, -48, 118, 4, 25, 71, -110, 25, -96, 78, 69, 99, -76, 84, -98, -12, 21, -52, -60, 25, -71, 20, 118, -13, 70, -119, 24, 1, -62, 11, 101, 118, -25, -79, -76, -1, -88, 104, 114, 127, 14, 38, -92, -55, -97, -126, -60, 113, 107, -75, -114, 111, -69, -101, 64, 12, -97, -28, 68, 98, 23, 103, -125, 94, -39, -23, 23, 34, 67, 124, 73, 82, -18, -36, 86, -32, -78, -127, -34, 89, -92, 115, -71, -115, -84, -55, -69, -67, 15, 111, 45, 52, 8, 27, -125, -65, -58, -89, -102, 17, -39, 123, -62, 86, 122, -65, -83, 103, 20, -75, -89, 126, -67, 125, -92, -87, -67, 58, 75, 79, -90, -121, 98, -31, -45, -125, -33, -65, 85, 41, 57, -68, 57, -51, -10, 97, 14, 1, 12, 11, -118, -71, 64, -122, 82, -115, -51, -116, 106, -127, 53, 8, -60, -3, 88, -93, 68, -117, -83, 33, 87, -89, -83, -97, 51, 103, -114, -38, -14, -25, 16, -53, 59, -112, -38, -22, 52, -39, -8, 24, 72, -103, 122, -16, 123, -55, -51, 1, -62, -75, 86, -87, 54, -62, 19, -75, 87, 101, -84, -73, 83, -103, 33, 85, 67, -44, 15, 36, -20, 115, 31, 2, -26, -36, -77, 23, 46, -115, 70, 44, 58, 77, -126, 62, 102, -10, -99, 68, -92, 40, 59, 63, -121, 52, -61, -118, -26, -30, 69, -57, -77, -57, -114, -110, -18, 29, 74, -20, 49, -115, -52, 18, -1, -12, 51, -85, -38, -27, 123, 63, 96, 6, -87, 11, 47, -20, -8, -21, -90, -68, -63, -80, -8, -10, 30, 105, -87, 63, -120, -8, 10, -21, -116, 106, 58, 7, -100, -67, 97, -67, 84, 80, 58, -101, 49, -4, -127, -7, -120, -60, -45, 19, -120, -37, 72, 99, 113, -23, -116, 9, 20, 44, -107, 40, -87, 42, 68, -5, -51, 61, 99, -2, 80, -69, 101, 127, -45, -37, -116, 7, -42, 5, 50, 4, 70, -103, -27, -11, 15, -62, -45, -9, 36, 77, -64, 47, -105, -86, 24, -92, -33, -124, 74, -79, 58, 96, -68, -15, 75, 13, -26, -82, 35, 37, 47, -115, -66, -62, 113, 77, 82, 69, -104, -41, -40, 56, 69, 103, -51, -48, -118, 80, -92, -70, -28, -119, -62, -126, -32, 36, 16, 58, -112, 120, -61, 75, 89, 79, -106, 8, 3, -105, -111, -24, 16, -115, 100, -59, -106, -124, 11, -75, -9, 76, -39, -38, -127, 30, 0, -109, 115, -65, 124, 34, 102, 111, 116, -117, -50, -1, -122, -90, -90, -104, 7, -6, -58, 14, 120, 107, -93, 34, -83, 44, 2, -45, 13, 85, 66, 9, -28, -25, -4, 19, 99, 31, 3, 119, 35, -97, 1, -117, -23, 22, 61, -34, 24, 66, 126, 14, -84, 81, 4, 127, -65, 11, 85, 19, -28, 67, -114, 98, -107, 30, -18, 29, 6, 75, 43, -96, -60, -45, -87, 119, -123, 98, 100, 102, 97, -101, -64, 58, -56, -124, 102, 125, -74, -33, 31, 77, 56, 81, 25, -63, 108, -123, 105, -88, -11, 12, 92, -113, 48, 88, 23, 76, -29, 47, -78, 101, -123, -100, 122, 43, 77, -21, 6, -9, 56, 109, -123, 75, -89, -111, -101, 26, 43, -89, 64, -25, 120, 45, -111, -106, 99, 114, 35, 127, -72, -120, -57, 1, -69, -105, 37, 114, -120, -81, 115, 25, 41, -25, 111, -82, 42, -99, 19, -9, -7, -87, 122, 77, -127, 31, -72, -96, -111, -9, 10, -109, -6, 6, -109, 32, 61, -57, 70, -21, 10, -53, 22, 54, -97, -20, 2, 14, 100, -54, -125, 97, 18, -19, 94, 20, -2, -60, 84, 121, 77, -26, -22, -118, -59, 44, -116, 16, 0, -7, 125, 124, 76, 28, -21, 40, -45, -35, -18, -49, -47, 75, -124, -93, -121, 64, -15, 22, -7, -107, 100, 48, -97, 102, 33, 54, -5, 29, -50, 87, -112, 71, 47, 112, 102, 21, 72, 124, 52, 24, -38, 77, 27, 71, 35, -112, -28, 8, 124, 48, -60, 7, 71, 90, -107, -30, -51, 67, -80, -68, -22, -111, 31, 24, -62, -71, -83, 38, 51, -72, -37, 125, -111, -62, 112, -55, -38, 88, -9, 54, 95, 80, -73, 85, 73, -46, 84, 4, -62, -1, -27, -69, -41, -39, 17, 17, 85, 105, 76, 53, -47, 54, -125, 67, 78, 2, 1, 72, 32, 113, -95, 21, -6, 79, 94, 80, 18, 50, -43, -9, -16, -95, 56, -99, 117, -24, 90, 39, -6, -34, -70, 26, 17, 5, -7, 119, 82, -128, 126, 97, -46, -26, -87, -85, -52, 52, -72, 48, -112, 54, 118, -18, 43, 13, 66, -107, -57, -114, 25, 111, 83, -6, -73, 85, 18, -92, 40, 101, 65, -95, 92, -56, 5, -124, 0, 75, -106, -112, 8, -89, -6, 27, -104, 122, 123, -26, 78, -23, 2, 114, -23, -119, -38, -78, -26, 57, 126, 54, 50, 94, 3, 44, 58, -84, 93, -72, -5, 100, -47, -25, 115, -83, 64, 92, 80, -76, 95, -102, 39, -67, 8, -82, 121, 79, 25, -113, 31, -119, 5, 62, 59, -87, 5, -18, -116, 118, 78, -106, 20, 27, 64, -8, -76, 92, -39, -14, -66, -4, -114, 80, 11, 60, 20, 85, 44, 127, 44, 120, 20, 14, -50, 39, 37, 9, 90, -124, 53, -59, 121, -16, -8, -118, -102, -111, 90, -126, 26, -72, -91, -46, -76, -18, -97, 77, -122, 113, 89, 76, 35, -24, 20, -57, 122, -1, 70, -83, 106, 69, 89, 26, -55, 111, -100, -22, -12, -91, 35, 26, 64, -27, 104, -114, 2, 39, 72, -96, 84, 65, -101, -32, -88, -114, -104, 65, 117, 118, 75, 97, -41, -26, 83, -31, 92, -57, -105, -11, -79, 61, 120, 65, -74, -118, 90, -14, 62, 94, -26, 46, -81, 23, 123, -92, 105, 109, 12, -32, 12, 69, -42, -106, 109, 125, -33, -28, -37, -116, 126, -78, -104, 37, 75, 125, 101, -109, 123, -23, -40, -37, -36, -19, -104, 25, 69, 25, 105, 24, -40, 11, -38, -53, 103, 4, 0, -113, -83, -39, -112, 110, 27, -13, 106, 122, -48, 57, -61, 52, -75, -115, 76, -110, -27, -36, -95, -29, -53, 110, 92, -55, 22, -105, 124, -116, 84, -64, 74, -92, 60, 21, 96, 63, 7, 72, -124, -121, -101, 64, -68, -72, -83, 96, -16, 119, -71, -58, 103, 78, 97, -92, 65, 119, -86, -7, -32, 33, 102, -55, 45, -128, 31, 70, -113, -83, -39, -69, 87, 112, 71, -125, 126, -11, 113, -15, 114, 74, 37, -60, -38, 90, -67, -40, -34, -3, -83, -29, -4, -53, -53, 55, -94, 24, -9, 29, 102, 4, -18, -34, -9, -6, 62, -96, 96, 2, -28, -40, -22, 41, 80, 102, 1, 33, 119, -110, -74, -111, 62, -84, 68, -108, 74, -37, -15, -73, -102, 125, -35, 99, 50, 60, 0, -20, -32, 115, 50, 125, -67, 1, -92, 80, 63, -121, -32, -76, -122, -37, 119, -3, 40, 61, -9, -124, 44, 102, -88, -3, 0, 7, -70, -123, -6, 0, -38, 41, 25, -83, -5, 48, 11, 108, -69, -11, 4, 111, 66, -71, -65, 126, -124, -107, 85, 109, -11, -38, 110, -17, 13, -22, -93, 60, -104, -30, 4, -51, 97, 117, -41, -123, -74, 30, -44, 55, -1, -36, 123, -122, 67, -71, 27, 60, 87, 29, -60, -88, -9, 120, -61, 35, 109, -43, 35, 101, 103, -124, -51, -85, -1, 75, -126, -34, 68, 5, 118, 85, 20, -112, 116, 92, -88, -55, 121, 98, 64, -46, -58, -115, -105, 109, -58, -99, -53, -96, -86, 31, -5, 48, -48, 51, 97, 71, 87, -83, 57, 106, 69, -47, -35, 5, 53, 106, -71, 18, -65, -34, -19, -122, -23, 80, -103, 125, -58, 7, -72, 89, 8, -8, -11, 9, 119, 97, 52, 93, 67, -123, -66, 20, -82, -123, -96, -75, -93, -118, -92, 35, 57, 63, -87, -37, 109, -106, 52, -21, 36, 23, 34, -54, 95, 44, 17, 25, 71, -119, 95, -4, 92, 122, 58, 30, 69, -76, 67, 107, -14, 30, -13, 17, 45, 103, 101, 65, 49, -64, -85, -11, 107, -69, -48, -21, 86, 102, 126, -79, 59, -108, 108, -63, 42, -3, 64, -64, -41, -104, -25, -41, -9, 89, 63, -32, -35, -78, 67, 127, 62, -21, 123, 20, -10, -117, 62, 84, 10, 122, 71, -26, -122, -98, 52, 19, -25, -55, -21, -103, 123, 26, -37, 118, -125, -50, -23, 121, -118, -72, 68, -67, -26, 90, 71, 83, -74, 13, -108, 63, -50, -24, 40, 55, 14, -93, 68, -61, -33, 94, -24, -59, -89, -16, -36, -101, -125, -43, -35, 73, 17, -77, 87, -42, 89, 85, -15, 31, 4, -83, -104, 93, -70, 66, -84, 106, -2, -114, -64, -64, -25, -23, -22, -116, 82, -83, 86, -38, -27, -91, 9, 86, -97, 51, 17, -37, -78, 33, 74, 24, -121, -42, -88, 42, -16, -55, 114, 107, 98, -24, -39, -119, 46, -68, -68, -9, -104, -88, 100, -122, -127, 54, -51, 100, 3, -80, -125, -113, 86, -118, -58, -110, -106, 101, -97, 103, 113, 114, 29, 46, -9, -32, -92, 116, -115, 58, -11, -33, 107, -66, 63, -57, 19, 25, 64, 46, -84, 120, 41, -53, 23, 56, -67, -76, 111, -91, 123, 27, 0, -21, 73, -89, -63, 14, 23, 123, 54, 86, 22, -61, 102, 88, 26, 60, 37, -127, 115, 125, 31, 34, 70, -82, 100, 87, -33, -89, -21, -45, -13, 84, -27, -120, 116, 102, 118, 9, 18, -65, -99, 98, 3, -28, 58, 25, -14, 106, 60, -87, 115, -63, 53, 15, -60, 7, -111, 102, 106, 102, 25, -36, 27, 79, 49, -90, 31, -44, -90, -77, -55, 122, 75, -15, -67, -46, -36, -76, 50, -36, -26, 52, -61, -65, 64, 2, 40, -103, 35, 5, 93, 85, -91, 63, -75, -83, 115, -103, 11, -88, 5, -35, 63, -47, -8, -93, 110, -29, 124, -26, 82, -118, 125, 104, 92, 16, -56, 30, 61, -52, 39, -111, 10, 92, 96, 14, -96, 29, -3, 26, 77, 28, -70, 23, -74, 104, 101, 117, 39, -66, 62, 101, -88, 57, 103, -61, 98, -14, -65, -127, -124, -42, 44, -31, 64, -23, -51, 86, -104, 31, -21, 69, 73, -54, 81, -3, -61, -81, -95, 43, 121, 0, 25, -107, 56, -104, 79, -95, 68, 57, -96, -121, 36, -23, -30, -109, -3, 11, 69, 81, -111, 24, -75, 119, 50, 38, -56, -106, -66, 16, 97, 30, 86, 62, -32, -116, 62, 97, 29, -67, 45, -124, -36, -87, -97, 92, -31, 107, -23, 33, 45, -71, 7, 116, -40, -90, -93, 41, 81, 12, 125, 115, -89, -77, 5, 9, 126, -7, -66, 91, -55, -66, -124, 53, -1, -107, -107, 92, 16, -119, -114, 28, 6, -27, 126, 40, 93, 73, -83, 64, -83, 2, 14, 80, 93, -29, 88, 8, -41, -52, -88, -20, 65, 96, 107, 29, -89, -82, 0, 59, 1, 118, 46, 82, 26, 4, -11, -69, -100, -70, 42, -101, -97, 116, -55, -2, -63, -6, -25, -73, 80, 44, 93, 122, -107, -61, 46, -75, 62, -34, -1, -101, 82, 120, -18, -5, -75, -34, 89, 93, 106, 65, 97, 98, -69, -12, -3, 57, 115, -40, -113, 92, -84, 113, 104, -106, 73, -108, 21, -15, -37, -124, -80, 118, -106, 114, -79, -121, -12, 4, -7, -26, 80, -25, -52, -81, 116, 7, 54, -51, -11, -46, -119, 114, 58, -78, -67, 35, -24, -110, 64, -98, 121, 125, -59, 27, 97, -115, 69, 32, 0, 91, 28, 23, -44, -72, -68, -116, -82, 17, -34, -3, 106, -9, -90, -98, -17, -76, -89, -104, -20, 121, 48, -99, -58, -88, 93, 42, -80, -102, 50, 80, -30, -30, 93, 31, 36, 65, -32, 101, -11, 46, 114, 39, -80, -65, 79, 125, -13, -1, -25, 102, 53, -50, -32, -111, -38, -43, -52, -108, 32, -119, 112, 19, -74, 119, 70, 63, 36, 4, -114, 33, -51, 96, -100, -12, 20, -90, 38, -98, -90, -90, 61, 67, 76, -76, -21, -103, 42, -126, -13, 48, 66, 4, -5, -75, -73, 41, -108, 58, 23, -46, 22, 79, -45, -62, -104, 107, -76, 106, 73, 118, 122, -82, 86, -76, -113, 120, 65, -95, 37, -110, 21, -85, 106, 33, 22, -121, 10, 43, -75, -29, 75, -14, 110, -120, -123, -125, -63, -48, -27, -57, 125, 51, 100, 109, 17, 112, 101, -66, 122, 33, -122, -45, 118, -12, -93, -51, -126, -3, 91, 67, -27, 99, 80, -55, -73, 74, 125, -80, -13, -115, -77, -88, -27, 57, -124, -74, -118, -107, 82, -4, 33, -10, -67, -73, 91, 31, -121, 86, -97, 77, 7, 43, 43, 125, 15, -11, -92, 91, -108, 39, 42, -10, 11, 26, 126, 74, 74, 29, 77, -81, -109, 65, 118, 102, -36, 18, 79, -29, 34, -49, -115, 98, 122, -17, -4, -89, 9, -81, -121, -72, -18, 79, -7, -80, 105, 79, -110, 111, -51, -24, -26, 23, 110, 64, 79, -77, -90, -30, -110, -88, 1, 56, 102, -112, -73, 40, 81, 5, 109, -62, 119, -126, 18, -56, -46, -112, -80, -125, 95, -63, 97, 116, 120, 22, -69, 51, -83, 88, -28, -127, -51, -128, 104, -106, -16, -119, -102, 35, -58, -125, 123, 106, 111, 82, 76, -84, 67, -47, -79, 98, 119, -36, -83, 83, 91, 64, 83, -25, 86, 35, -70, -73, 122, 14, 64, -45, -41, -119, -73, -116, 95, -120, -104, 45, 53, -61, -58, 52, 42, 89, -37, -13, -125, 32, -23, -63, -11, -67, -87, -109, -118, 100, 3, -61, -85, 50, -15, -110, 121, 56, 106, -60, -118, 2, -100, 89, -2, -88, 7, 34, 37, 46, -108, 50, 8, -50, -117, -27, 32, 104, -60, -32, -55, 22, -68, 100, 44, -94, -28, -11, -59, -37, -128, -93, -15, -45, 83, -20, -78, -34, -23, 12, -13, 70, -36, 99, -62, 73, -53, -71, -4, -42, 118, -110, 21, -45, -22, -94, -84, -39, 1, 83, -78, 39, -25, 86, 20, -61, 64, -14, 5, 57, -8, -60, 75, 46, -65, 49, 33, 8, -26, 59, 82, -72, 3, 4, -68, 36, -13, 87, 33, -115, -10, 29, 64, -19, 112, -101, -83, -25, -94, -84, 53, -104, -100, -65, -69, -20, 109, 67, -53, -62, -59, -66, 56, 51, 83, 10, -58, 98, -14, -72, -112, 122, 107, 61, -29, -84, 65, 81, -5, -61, 65, 9, -75, -33, -83, -60, -69, 114, -63, 122, 53, 27, -102, 103, -30, -112, -98, -117, 92, 62, 53, 87, -97, -68, 94, 56, 60, 19, -76, -8, -87, 0, -7, -128, 5, 50, 40, 63, 100, 11, 81, 4, 5, -3, -55, 3, 75, -104, 55, 7, 27, 65, 37, -14, 87, 23, -112, -1, 75, 22, 11, 108, -9, -34, 117, 12, 95, -42, 84, 19, -76, 48, -102, 81, 99, -21, 84, -55, 65, -28, -57, -109, 108, 36, 127, -46, -88, 110, -48, -80, -87, 88, 8, -64, 16, 61, 6, 74, 16, 93, -95, 126, 14, 107, -19, 86, 58, 24, 106, 109, -110, -117, -25, -55, -121, 65, 104, 48, -64, 48, -116, -23, 5, -11, 6, 48, 11, 13, 31, -49, -116, -65, -67, 92, 10, 4, 93, -74, 19, 105, -119, 31, -94, 98, 54, 70, 26, 116, -63, 82, -14, -4, -45, -23, -118, 57, 102, -17, 45, 75, 55, 27, 19, 73, -44, -33, 21, 53, 99, -113, -92, 36, -52, 47, -16, 23, -17, 69, -46, -11, -112, 74, 73, 32, -55, 65, 124, -86, 15, -115, -20, -74, 69, 107, 107, -35, 127, 117, 30, -86, 15, -49, -85, 109, -44, -35, -55, -67, -75, -58, -48, -57, 92, -125, -127, -41, 78, 100, -16, 33, -125, -67, 77, 13, 68, -64, 88, 67, -94, -116, 21, -5, 94, -49, -34, -17, 96, -114, -116, 32, -126, -5, -106, -67, -44, 90, 64, 120, 0, -15, -126, -90, -20, 109, 96, -61, 81, 43, -105, 33, 51, -39, -85, 112, -105, 20, -19, 15, 59, -91, 31, 81, 15, 20, 2, 44, 20, -2, -14, -111, 116, 30, -96, -102, -88, -123, -14, 83, -10, -21, -52, 19, 71, 52, 54, 105, -58, 71, 90, -45, 44, 120, -95, 60, 126, -68, 1, 67, -81, -53, -59, -117, -85, -125, 86, -33, 56, 2, -2, 25, 96, 3, 4, -91, -8, -125, -41, -78, 96, -92, 44, 3, -76, -87, -109, -32, -30, -94, 82, 77, -70, -70, -128, -77, 15, -26, -108, -61, -56, -73, 12, -90, -41, 113, 2, -106, 105, -77, -110, -85, 9, -72, -124, 96, -42, 122, 0, 42, 39, -118, -114, 83, -125, -2, 31, -123, 38, -20, 20, -83, -91, 74, 98, -72, -13, -107, 117, 3, 2, 61, -35, -14, 111, 3, -61, 30, -67, 106, -7, 105, 112, 114, 22, -56, -14, -81, -68, -23, -43, 113, -27, -27, -128, -109, -33, -92, -84, -127, 2, -115, -56, -73, 72, 102, 121, -38, 17, -11, 63, 123, -100, -27, 35, 81, -35, -62, 39, 71, -61, 125, 21, 61, -42, 62, -34, 4, 23, 26, -1, 60, 76, 55, -72, -58, 38, 92, 121, -105, -70, -124, -69, 25, -117, -82, -58, 51, 76, -77, -53, -40, -47, -67, -92, 40, -111, 45, -41, -75, 34, -68, -45, 13, 79, 52, -128, -55, 70, 9, 101, -122, 51, 49, 62, 9, -100, -23, -70, -94, 49, 82, -86, 118, 118, -75, -99, 11, 14, 42, 102, -57, -110, 34, 70, 1, 41, 96, 6, 2, -55, -99, 54, -53, 82, 84, 113, -108, 41, 103, -13, 90, 86, 29, -117, 18, -20, 40, -114, -42, -4, -51, 124, 84, -90, -98, 12, -70, -103, -11, 104, 77, 38, -19, 92, 106, 19, 59, 57, 100, 35, 11, -87, 109, -40, -63, 25, -67, 51, 43, -72, -17, 82, 19, -127, 44, -124, -24, 42, -98, 108, 18, 115, 29, 13, 8, 48, 35, -108, 75, 106, 120, 20, -52, 36, 62, 20, 1, -18, -105, 124, -62, -95, -53, -66, 51, -80, -89, -42, -128, -100, -43, -93, -100, -77, -61, -3, -59, 65, -22, -113, 16, 112, -17, 20, -33, -14, 9, -9, -127, -10, 67, 21, 8, 120, 29, 9, 126, -5, -55, 18, 65, -107, 62, 98, -27, -33, -67, 112, 23, 73, 26, -25, 113, -6, 46, -110, 82, 36, 108, 54, 81, 20, 120, -105, -65, 24, 96, 14, -72, -87, -19, -20, 104, -126, 100, -64, -107, -6, 68, -36, -93, 41, -72, 59, -111, 117, 26, 41, 34, 117, -52, 87, 44, 11, -36, -128, -2, -40, -49, 100, -60, -22, 42, 108, 35, -120, -23, 61, 13, -91, -123, 107, -112, -53, 120, -93, 13, -71, -73, -4, -27, -85, 36, -49, -128, -40, -113, 88, 85, 126, 58, -71, -100, -4, -8, -59, 22, 54, -88, -110, 106, 42, 16, 39, 54, -25, -35, 46, -21, -123, 5, -104, -41, 49, -20, 118, 69, -26, 108, 14, 54, 55, -106, 0, 24, 51, 46, 106, 34, -13, -45, -102, 83, 118, -16, -79, 78, 72, -53, -29, 92, 92, -89, 25, 118, -110, -22, 70, 63, -61, 59, -73, -103, -50, -18, 15, 97, -42, -91, 112, -77, 38, -68, 49, -64, 9, 118, -52, -120, -57, 12, 41, -117, -45, 69, -95, 82, -66, -20, -4, 20, -103, 67, -53, 41, -55, 22, -23, -107, 61, 75, 117, 53, -37, 52, -81, -95, -56, -65, -12, -98, 100, 37, -104, -63, 81, 44, -44, 90, -21, -62, 6, 57, -126, 109, -43, -27, -50, 64, -1, 22, -11, -118, 110, 18, -43, 7, -10, -39, -19, -103, -24, -102, -48, -31, -71, -109, -69, 126, -52, -108, -48, -100, 14, 97, -35, 29, -90, 64, 87, -80, -95, 24, 98, -86, -105, -80, -59, -64, 41, -76, 119, -43, 22, 32, -17, 9, -36, 4, 52, -10, -41, 90, -110, -74, -25, -115, -20, 118, 27, -54, 47, 76, 125, 36, -48, 80, 110, -11, 45, -28, 94, 13, -22, -105, 66, -54, 11, 22, 32, 61, -88, 79, -9, -112, -55, 15, -62, 97, -43, -52, -78, 35, -40, 111, -49, 120, 100, 25, 5, -33, 111, 69, 31, -112, 116, 73, 75, 8, 122, 34, 5, 98, -62, -34, -1, -62, 39, 79, -16, -121, 37, -100, -107, -100, -113, -108, 123, 5, 20, 45, -41, -126, -12, -125, -64, 90, -128, -40, -102, -73, -14, 99, 85, -79, 68, 11, -51, 10, 92, 89, -85, -8, 43, 35, -123, -74, 79, 101, -119, 72, -39, 105, -86, -125, 105, 8, 123, 56, 63, 26, 29, 75, -65, 4, 47, -58, 54, -112, -51, 119, -2, 49, 0, 23, 88, 97, 15, 25, 78, 15, 85, -37, 72, 53, -33, 127, 21, -19, 41, -47, 67, 101, 55, -44, -46, -43, -120, 6, -9, 10, -11, -37, 109, -99, 99, -83, 66, 36, 55, -105, -106, -95, 6, -11, 25, -116, 87, 7, -24, 20, 38, 11, 54, -3, -22, -35, -86, -9, 92, -120, 10, -120, -59, 126, 69, 92, 108, 92, 5, 31, 15, -59, -86, 82, -10, 126, 107, 17, -16, 20, -46, -27, 32, 87, -22, 52, 32, 105, -88, -2, -23, -18, 96, -68, 127, -84, 67, -120, -17, 26, 107, 92, 79, -47, 105, 41, 40, -58, 52, 97, -119, -113, -120, -115, -104, -38, 8, -126, -12, -113, 72, 81, 27, -85, -21, 118, 57, -125, -128, 24, -30, 19, -86, 21, 31, 69, 120, -45, -70, 27, 51, 31, -96, -118, -58, -11, -114, -95, -4, 25, -91, 32, -125, 88, 92, -76, 13, -74, 77, -11, 8, 118, 38, 110, 61, -24, 45, 80, -50, 51, 99, 55, -39, -63, -33, -39, 0, 82, 79, 73, 51, 19, -13, 8, -79, -37, -3, 119, -28, -2, -111, 36, -30, 25, 38, 59, 84, 37, 90, -18, 61, -33, 92, 42, -63, -69, 43, 41, -100, 4, -43, 118, -50, -90, -11, 108, 38, -91, 68, 50, -69, -84, 23, 77, 17, -7, -73, -9, 10, 74, 91, -66, 109, -65, 91, -106, 106, 53, 22, 127, 111, -80, -86, 84, 90, 58, 81, -45, 71, 8, -4, 1, -6, -108, 111, 97, -79, 43, 3, 89, -97, -56, -4, 91, -10, -42, 58, -72, 97, -40, 3, -118, -55, -107, 77, -83, 1, 38, 81, -36, 14, 42, 79, -14, 124, -50, -84, -17, -54, -22, 45, 101, -11, 10, 92, -110, -20, 68, -54, -91, 126, -15, -65, -51, -77, -13, -24, 13, -84, -109, 81, 7, -71, 118, 66, 34, -78, 38, -73, 122, 21, -26, 88, 76, -90, -77, -97, 39, 57, 79, 77, -69, -1, 42, 90, 110, -21, 79, -16, 38, -113, 93, 65, -46, -47, -25, -120, 109, -20, 83, 52, 126, -92, 73, -62, -44, 70, -11, -121, -4, -100, 27, 53, -125, 62, 44, 20, 67, -41, 85, -106, 124, -38, 44, -57, 39, -29, 66, 59, 58, 109, 127, 35, 33, -43, -71, 28, -90, -26, 17, -70, 69, 3, -31, -33, 11, 113, -114, -82, -89, -70, -115, -76, 100, 78, -45, 126, 8, 75, -35, -54, 85, 102, 116, -10, -41, 59, 72, 123, 126, 94, 123, -41, 91, 83, 54, 49, 28, 49, -52, -110, -128, 64, 42, -20, -128, -92, -83, -17, 92, -95, 113, 22, 59, 18, -112, 19, -18, 31, -18, 29, -94, 99, -57, 48, 60, -42, -109, -6, 42, 108, -63, 27, -23, 24, 39, 122, -44, -39, -28, -13, -73, -88, -44, -116, -69, 13, 122, 97, 0, -85, 45, 30, 115, 51, -9, 120, 23, 38, -14, 38, -33, 34, -75, -62, 86, -106, 107, 61, -12, -99, 8, -114, 99, -79, 33, -33, -47, -6, 65, -106, -35, -107, -120, -23, -15, -120, -124, 68, -49, 90, 7, 117, -115, -119, 12, -48, -6, -126, 32, 59, 105, 27, -19, -59, -38, -4, -27, 59, -89, 122, 80, 101, -48, -12, 85, -118, -29, -93, -108, 97, 98, -29, -81, -66, -24, -87, 51, 121, 16, 69, 42, 18, -111, 105, -103, -33, -115, -43, 55, -38, 33, -105, 6, 121, -36, 6, -113, -69, 15, -76, 1, 84, -17, -27, 6, -75, 50, -107, 51, -34, -5, -81, -56, 43, 19, -63, -22, 107, -28, 50, -72, 116, 35, 44, 22, 87, -69, -30, 8, -11, -94, 98, 113, 49, 106, 120, -38, 86, 59, -89, -30, 11, -43, 85, -31, -75, -60, -112, -52, -85, 108, 16, 111, 4, -82, 71, -16, -28, 63, 65, -61, -26, -89, 90, 90, -3, 19, 43, -22, -84, -99, 23, 101, -91, -89, 24, 1, -93, -51, 9, 39, 100, -107, 118, 105, 28, 84, -59, -84, 120, 116, -108, 7, 97, 33, -50, 70, -64, -125, -73, -42, 109, -69, 25, 78, -36, -122, -18, -47, 13, -12, -52, 119, -109, -118, 101, 15, 72, 93, -112, -123, 103, 32, -43, 91, -42, 8, 112, 114, 96, -117, -31, 19, -23, -118, -44, 15, -93, 109, 119, -30, -101, 72, 7, -5, -119, 54, -108, -82, -24, -27, 106, -111, -55, -53, -120, 54, -4, 14, -63, 0, 25, -49, 68, -105, 12, -100, 112, 15, -87, -67, 61, 70, 67, -120, 26, -46, 71, -24, 94, -92, 1, -92, 103, 91, -4, 102, 1, -23, -64, 85, -87, 68, -97, 52, -84, 6, -31, -66, -125, -122, -16, 14, -101, -114, 6, -103, 118, -12, 80, 13, -50, 123, -113, 126, -103, -29, 80, -10, 69, -20, 30, 90, 66, -3, -108, -126, 52, -70, -86, 108, -49, 118, -66, -21, -29, -58, 88, 49, -47, 125, 86, -4, -1, -79, -44, -8, 97, 59, 16, -80, 42, -65, 81, -18, 91, -99, 91, 55, -13, 96, -31, 8, 31, -24, -70, 102, 13, -52, 66, 59, -73, 17, -70, 100, 120, -2, -42, -67, -1, -54, 1, -28, 127, -72, 30, -66, 95, -92, -70, -112, 21, -96, -100, 58, 1, 8, 12, -13, 97, 72, 73, 57, -55, -96, -88, -6, -14, -89, -30, -73, 6, 41, -13, 98, 31, 35, 53, -35, -49, -94, -46, 21, 17, -25, -70, -100, 108, -37, -108, 14, -81, -96, 71, -35, 48, 87, 120, 69, 24, -121, 44, 21, -41, 31, 1, -17, -85, -127, 32, 60, 52, -50, -45, 106, -36, -67, -47, 94, 123, 40, 118, -16, 104, 13, 60, -27, -122, -34, 90, -62, 0, 58, 56, -79, -94, 5, 14, -33, 63, 53, 59, -32, -33, -60, -88, -65, -57, -21, -63, 68, -91, 38, 96, -59, -15, -30, -29, 20, 77, -88, -86, -40, -44, -51, 53, 49, 23, 89, -125, -31, -85, -15, 86, -81, -121, 52, -87, -37, -111, 9, -118, -14, -23, 127, -26, -12, 120, 61, -85, 41, 104, -62, 30, -90, 37, 76, 113, -54, 57, 31, -45, -24, 31, -17, -10, -11, -120, 10, 126, -83, 59, -67, 69, 28, 18, -65, 36, -79, -123, 100, 75, 15, -21, -83, -57, -102, 20, 120, 41, -79, -120, 87, -28, -23, 67, 29, -54, -57, -20, -19, -51, -117, -120, -91, 84, -25, 45, -75, -80, -23, -101, -56, -36, 4, 62, 126, -90, -91, 92, 117, -51, -68, 2, -115, 118, -58, 46, 126, 33, -42, 57, 75, 92, 54, 0, 102, 36, -118, 96, 77, -28, -94, -109, 112, 72, -91, -50, 71, -73, -16, -76, -110, -48, 63, 107, -42, 3, -125, 94, -69, 26, -12, 125, -44, -78, 44, -9, 84, -80, -50, 121, 127, -65, 19, 21, 73, 20, 116, -75, 46, 14, -62, 88, -5, 17, 65, 85, -125, -37, 0, 59, 60, -89, -7, -3, 75, -114, -102, 27, -111, 72, 50, -28, -55, -42, 41, -110, -50, 46, 101, -107, 20, -68, 68, 38, -33, 7, -17, 117, -23, 99, 125, 103, -105, 12, 81, -44, 47, 115, -120, -44, 100, 126, -57, -56, 19, -55, 63, 110, 102, -78, -117, 0, 57, 123, -87, -42, -76, -57, 108, 127, 48, 93, 126, 37, -60, 92, -98, -79, 73, 76, -88, 96, 13, 40, 112, -105, 8, -67, -49, -25, 94, 109, -115, -30, -53, 54, -109, 68, 7, -119, -82, -94, -110, 7, -34, 37, -47, -90, -73, 116, -108, -20, -1, -125, 106, -44, 64, 40, 2, 90, -36, -85, 120, 21, 81, -4, -122, -95, 120, 42, -115, -51, 7, -114, -61, 120, -11, -54, -88, -55, 80, 32, -108, -104, 51, 22, 115, -43, 67, -104, 96, -44, 47, -62, -61, -64, -70, 127, -1, -91, -124, 80, -5, -97, -88, 13, 60, 52, 13, -46, 69, -72, 0, -89, 76, 74, -113, -85, -5, 101, 0, -26, -54, 52, -40, -97, -1, 14, -65, -73, 44, -43, -13, -122, -48, 26, -86, -29, -97, -34, -76, 107, 72, 24, 65, 93, 18, -79, -27, 61, -96, -80, 101, 54, 85, -122, -51, 7, 26, 11, -43, 43, -109, 61, -47, -40, -90, -90, 119, -46, 111, -64, -47, 34, 12, -21, -14, -63, 115, 19, -103, 80, 88, -79, 41, -89, -79, 75, 25, -70, -72, 100, -65, -49, 118, -90, 93, -125, -96, 86, -105, 108, -110, -78, 4, 33, -11, -17, -98, 38, -79, 9, 103, -61, -125, -26, -106, -120, 9, 22, -54, 55, 77, 20, 13, 52, 117, -78, -102, 14, -127, -43, 101, -42, 64, -34, 95, -87, -111, 9, -36, 97, 21, -4, 30, -19, -22, -38, -119, 75, -126, -21, 57, -40, 0, 30, -43, 112, 115, 84, 52, -111, -40, -87, 17, -49, -111, 37, 67, 114, -122, 63, -90, 20, -85, -2, 66, -55, -102, 102, 11, -61, -125, -12, -87, -96, 85, 84, -125, 9, -57, 49, 121, 106, 29, 49, -3, 16, 71, -76, -51, -40, 57, 29, 30, 78, 75, -114, -58, -42, -63, 64, 36, -21, -8, 6, 118, 77, -15, 3, -56, -116, 79, -79, 1, 13, -91, -85, -115, 37, -36, -46, -7, -66, -95, 121, 60, -28, -52, -104, 37, -116, 1, 85, -74, -69, -60, 8, -97, -98, -94, 46, 63, -84, 25, 110, -58, 109, -103, -52, -40, -33, 71, -113, -44, 37, -88, 94, 124, -45, 102, 9, 74, 85, -106, 75, 127, 9, -48, 32, -5, 26, 22, -117, 53, -47, -48, -98, -85, -1, 7, -106, 57, 7, -60, 58, -121, 82, -109, 29, -41, -14, -122, -58, 27, 12, 71, 80, 77, 60, -18, -2, 10, 109, 97, 96, -100, -10, 58, -42, -89, -23, 23, 46, 54, 81, 92, -56, 27, 99, -80, -72, -45, -45, -108, -40, 81, -115, -102, 33, -60, 124, 52, 55, 79, 113, 118, 45, -45, -117, -42, 1, -113, 52, 21, -55, 20, -105, -111, -58, 82, -20, 41, -79, 75, -26, -81, 35, -74, 28, 40, -45, -125, 30, 73, 27, 79, -84, 39, 76, -1, -52, -41, -55, -88, 94, 13, 85, -106, -85, -43, -30, 120, -110, -84, -91, -3, -114, -2, 62, 6, -41, -15, -69, -4, 107, -89, -34, -16, -56, -32, -3, -103, -17, -69, -55, 3, -42, -90, 70, -73, 75, 81, 16, 95, 127, 127, -45, 117, 93, -10, 98, -100, -97, 63, 78, 120, -60, -5, 56, 42, -15, -51, 54, -91, 101, 43, -6, 47, 126, 95, -23, -52, 36, -102, -75, -16, 55, 49, 35, 34, 31, -112, -66, 51, 47, 126, -37, -85, -96, 125, -41, 19, 92, 51, -36, 14, 121, -96, 51, -30, -45, -95, -22, 121, -109, -85, -113, -45, -108, -50, -12, -16, 106, -34, -99, -63, 45, 36, 37, 110, -68, 15, 117, -5, -106, -46, 119, 97, 37, -98, 53, -88, 122, -110, -26, 92, 87, 105, 26, 51, -28, 113, -98, -20, -63, -108, -117, -60, 45, 85, 100, -18, 26, -1, -126, 49, -86, 36, -94, 50, -71, 120, 13, -115, 75, 90, -57, 4, 63, -73, -39, -103, -124, -104, 17, -75, -92, 126, 35, 111, -85, 43, 69, -16, -4, -120, 37, -112, -15, 85, -33, 67, -84, -83, -103, 53, -103, -19, 103, 87, 91, 51, 36, 38, 44, -51, -104, -127, -59, 126, -6, 44, 10, 107, -32, 45, 42, -19, -17, 127, -61, 57, 16, 68, -22, -112, 40, 111, -125, 29, -81, 108, 10, 24, -9, 76, 46, -123, 31, 20, -62, -95, 65, 54, -88, -127, 49, 64, -7, -69, -116, 95, 110, 38, 38, 78, -51, -47, -41, -105, -62, 94, -42, 27, -105, -14, 72, -46, 7, -50, -57, 28, -75, -18, -63, -58, 0, 1, -76, 44, -64, 67, -62, -105, -48, -84, 96, 75, 102, -66, 82, -128, -14, -108, 82, 2, 15, -123, 2, 35, 116, -31, -65, -116, -101, -78, 89, -92, 110, -29, -47, 48, 48, -124, 33, -14, -70, -68, 12, -115, -32, -3, 9, -46, 5, -36, -20, 56, -52, -42, 25, -84, -50, 127, -42, 38, 89, -70, 122, -82, 6, -66, -106, 48, 1, -125, -44, 6, -14, -9, 56, -96, -113, 43, 84, -4, -13, 77, -3, 97, -15, -26, -62, 94, 57, -13, 98, 126, -42, -68, -88, 82, -114, -41, -72, -47, -54, -7, -98, -90, -54, 3, -111, 88, 46, 117, -59, -106, -94, 103, 117, 57, -79, 52, 81, 53, -92, -28, 75, 77, -5, 79, 108, -126, -105, 3, 26, -90, -61, -96, 117, -110, -34, 58, -52, 47, -11, -50, 127, 21, -97, -58, -40, 117, 127, -70, 6, 6, -28, 14, 1, 46, 57, -59, -27, 36, 14, 75, 0, 62, -9, -110, 9, 51, 95, -24, 75, 101, 95, 86, -31, 61, -87, -16, 42, -110, -121, 58, 62, 123, -128, -64, 111, 44, -10, -51, -89, -40, -28, 102, -9, -55, -24, 49, -125, -15, 80, 8, 40, -22, 98, -20, 45, 64, 18, -110, -93, -56, -3, -18, -78, 24, -48, 116, -106, -66, -86, 40, 38, 6, 13, -54, 10, -82, -55, -95, 86, -89, 43, -93, -124, 47, 58, 20, 7, -125, 8, 101, -62, -41, 62, -59, -59, -98, 49, 77, -124, 17, 57, -27, -113, 52, 49, -21, -116, 27, -40, 124, -117, 70, -110, -52, 76, -65, -8, 20, 32, -61, 109, -110, -5, 80, 68, -26, -71, -61, -100, -47, -57, 8, 125, -123, 74, -101, 35, 108, -92, -33, 37, 78, 95, -21, 17, 48, 103, -110, -67, 111, -49, 92, -49, 49, -61, -18, 69, 6, -49, -20, -66, 26, -45, -73, -62, -104, -48, 29, -120, 86, 100, 32, 74, 38, 55, -25, 59, 101, -21, 118, -120, -99, -112, 87, -9, 36, 127, -11, 122, 13, 53, 80, -26, 11, -97, -36, 1, 116, -42, 21, 97, -29, -74, 32, -18, 40, -55, -15, -29, 118, 104, -89, -39, 77, -1, -115, -14, 81, -126, -61, -127, 37, 9, -30, -94, 74, -113, -40, 74, -93, 107, -46, -42, 109, -127, 110, 45, 120, -21, -124, -5, -51, 62, 77, -119, -13, 20, -60, -68, -59, 54, -19, -44, -110, 84, -88, 42, -28, -4, 9, -127, -61, -83, -21, -58, 67, -65, -71, 21, -103, 74, -79, -116, 26, -60, 81, 70, 94, 122, 88, -54, 15, -77, -21, 91, 73, 42, -39, 80, 23, -97, -80, 71, -39, -109, 100, -72, -63, -30, -113, -124 );
    signal scenario_output : scenario_type :=( 124, -22, 127, 54, -128, -70, 14, 127, 86, -128, 52, 78, -51, 127, 21, -128, 87, 127, -128, 27, 122, -128, 122, -128, 127, -128, -128, 53, -126, -47, 100, 127, -78, -128, -74, -63, 12, -128, -94, 120, -128, 109, 32, -128, -128, 73, -128, -128, 127, 122, -108, -128, 127, 73, 127, -100, 127, -128, -116, 127, -125, 28, 119, -14, 127, -29, 64, 127, 22, -128, 1, 127, -128, 4, 127, -22, 127, -128, 104, 127, -128, -6, -126, -128, -121, -128, 42, 127, -128, 61, 127, 0, 73, -81, 127, 127, -103, -128, -128, -104, -128, -83, 65, 127, -117, -128, 25, 93, -7, -128, -128, 127, 127, -128, -128, 31, 87, -128, 49, 127, 41, 120, -128, -128, 105, 127, -39, -128, 42, 127, 5, -20, -128, -128, 127, -128, 127, 127, 55, 127, -30, -128, -13, -6, -35, -57, -4, 127, -94, -128, -38, 127, 66, 127, -122, 127, 58, -128, 127, 127, -128, 127, 127, -128, 62, 23, -128, -74, 127, 36, -60, -60, 127, 127, -51, 90, -128, -97, 127, 127, -79, 25, 76, -18, -128, -128, -19, 12, -128, 127, -25, -128, 116, 51, -120, -128, 127, 88, 92, 127, -128, 127, 85, -128, -128, 100, -11, -128, -123, 127, 127, 127, -128, -74, 13, -128, 86, -87, -99, 0, -128, -31, 127, -54, -86, 40, -128, -49, 1, -128, 10, 39, -128, -102, 127, -27, 54, 127, -128, -128, -128, 127, -20, -128, 74, 127, -128, 5, 127, 124, -7, -128, -65, -104, -128, 43, 71, 46, 119, -114, -91, -18, 127, 104, -97, 127, 127, 6, -92, -83, 127, 117, -128, 127, 127, -128, -12, 30, -128, -35, -128, 91, -120, -128, 46, -49, 127, 117, -1, -68, -87, 127, -128, -128, 127, -78, -15, 127, 127, -93, 86, -2, -70, 127, -128, -106, 127, -128, -128, 127, -42, 127, -49, 72, 127, -39, 127, -128, 54, 116, -128, -128, 127, 71, 127, 127, -128, 100, 127, 35, -128, -2, 94, 127, -128, 110, 51, -128, 127, -128, 17, -128, 127, 28, -128, -128, -56, -128, 28, -49, -128, -52, 5, -128, -128, -56, -38, -92, -17, 9, -62, 108, 75, -51, 127, 127, 127, 91, 127, -51, -128, 107, 127, -48, -23, -93, -47, -29, -128, -128, -128, -128, -75, 104, 127, 51, 127, 1, -128, 87, -128, -128, 127, 92, -128, 64, 46, 127, -69, -128, 127, 127, 28, -37, 127, 127, 18, 127, -77, -128, 15, 127, 31, 39, 26, 127, -128, -128, 81, -128, 127, 127, 127, -128, 77, -88, 58, -3, -60, -128, 127, -121, 127, 127, -71, -128, -128, -96, -78, 127, -112, -128, 38, 127, 127, 28, 11, 127, 127, 32, 44, 82, 115, -128, -128, 48, 127, 127, 36, 127, -116, -128, 88, 48, -128, 115, 12, 80, 127, -35, -65, -24, 64, 121, 55, 127, 127, -128, 106, -66, -128, 127, 127, -47, 30, -128, -128, 116, 18, -128, -128, 38, -128, -38, 17, 127, 127, -128, 127, 127, -128, -45, 47, 109, -128, 93, 127, -115, -128, 127, -128, 0, 73, -128, 72, 127, -128, -62, -18, -128, -22, -128, 57, 127, -32, 113, 127, -128, 108, -38, 80, 87, 49, -73, -128, 97, -30, 82, 127, -43, -3, -128, -22, 127, -39, -65, 4, 127, 11, -128, -78, 93, -128, 127, -128, -92, 127, -128, -95, 70, -77, -128, -4, 127, -34, -45, -14, 108, 55, 82, 22, 127, -126, 127, 127, -66, -128, -39, 127, 59, -128, -37, -86, -42, -128, 112, 127, 127, 43, 124, -128, -97, 127, -70, -128, 77, 127, 127, -100, -48, -59, -99, -23, -128, -128, 40, -3, -128, 127, 127, 127, 97, -128, -55, 127, -128, -128, 127, -128, 77, 127, -128, -122, 127, 66, -22, 127, 94, -128, -7, 24, 36, 127, -82, -128, -102, -128, 47, -128, 127, 127, -128, 127, 20, -128, -27, 91, 93, 37, 81, 127, -107, 11, 123, 96, -110, -65, 127, -128, 56, -120, -128, 127, -21, 99, 121, 127, -128, -128, 127, -128, -128, -5, -120, 92, -20, -14, 53, -128, 127, -128, -128, 127, -128, 127, 127, -126, 127, 64, -128, 32, 21, -57, 88, 127, -128, -66, -6, -128, 94, 127, 26, -58, -128, 127, 127, -102, -121, -72, 51, -65, -128, 127, 71, 55, -82, 127, -128, -42, -38, -48, -128, 127, 5, -1, 127, 39, -128, 90, -89, -128, 93, -60, -52, -117, 127, 107, 18, 127, -120, -128, 8, -7, -55, -128, 127, 127, 127, 10, 127, -103, -128, 127, -113, -30, 127, 125, 127, 7, 127, -128, -128, 111, -13, -128, -56, 42, -128, 127, 127, -87, 10, 19, -40, -128, 127, -128, -128, 127, 0, 53, 127, -54, -128, -74, -128, 55, -128, 43, 49, -128, 127, 127, -128, -5, 127, 14, -128, 127, 127, 63, -128, 127, 127, -5, 127, -117, 46, -37, -128, 107, -91, -97, -128, -62, -128, 123, 127, 87, 127, -39, -128, -73, 29, -30, -96, 127, 127, -55, 127, 127, 51, -128, -15, 87, -128, -128, 127, 127, -23, -21, 127, -128, -79, 127, -82, 72, 55, 127, -128, 127, -128, -65, 127, 9, -128, 127, 127, -128, -15, 127, -128, -128, 127, -110, -128, -128, 127, 30, -128, 127, 91, 127, 58, -128, -128, 62, 43, 23, -115, 127, -128, -68, -107, 41, 127, -83, 23, 127, 127, 17, -128, -128, -49, -92, -105, -128, 82, 127, -128, -89, 127, -128, -128, 127, 82, -128, 61, -128, 13, -128, -39, 127, 127, -128, 39, 74, -8, -128, -128, 127, 43, 48, -28, -74, -128, -9, -128, -128, -23, 127, 20, -35, 127, -25, -128, 127, -85, 127, 127, -128, 19, 127, 35, -128, 127, 3, -68, 127, -128, -2, 127, 102, 23, 127, -55, -128, -128, -128, -128, -17, -13, 43, 127, 127, 127, 127, -128, 17, -12, -128, -24, -78, 127, -128, 6, 127, 127, -128, 127, 127, 77, -128, 127, 127, -128, -47, 127, -128, -128, 127, -104, 127, 127, -128, -128, 127, 87, -102, -90, -128, -128, 103, -128, -128, 127, -69, -128, -66, -128, -116, -10, 35, 31, 127, 40, 55, -128, 127, 127, -128, -90, 63, -97, -128, 127, 127, -128, -128, 127, 127, -11, -65, -122, -26, -95, 127, -59, 86, 127, -128, 127, -111, -128, -69, -128, 127, -128, -128, 85, 49, -58, -128, -128, 114, 2, 57, 45, 85, -128, 127, -83, -36, -108, 127, -109, 127, 127, -128, 93, -12, -128, 127, -10, -128, -55, 127, -128, 127, 127, -128, 11, 127, 127, -128, 121, 127, 104, 29, 127, -128, 63, 23, -30, 127, -74, 127, -128, -128, -45, -10, -88, -128, 38, 127, -27, 127, 127, 88, 127, 5, -93, 2, 127, -100, -128, 23, 127, 5, 98, 127, -59, -85, 44, -41, -128, 15, -46, -128, -128, 127, 127, -11, -54, -89, -91, 127, 56, 76, 127, 65, -51, 127, -128, -128, 127, 127, -104, 85, 127, -120, 127, -128, -128, 127, 112, 34, 127, -108, 42, 3, -128, -128, 20, 127, 41, -128, 127, 77, -128, 127, 127, -128, -119, 127, -128, 86, 127, -128, -128, -31, 86, 54, 127, 127, -102, -45, 127, -94, -128, 48, -15, -128, -93, -40, 127, 99, -64, -128, -128, -34, 11, -128, -128, 127, 93, -128, 127, 127, -128, 127, 127, -88, 127, -128, -128, 127, -108, -90, 127, -128, 127, -18, -128, -128, -105, -128, 44, -14, -128, -128, 96, -128, -44, 115, 1, 127, -128, 66, 127, 127, 28, 127, -30, 13, -52, -128, -60, 106, -128, 22, -128, -128, 65, 127, -128, -128, 127, -128, -128, 127, 75, -5, 127, -128, 83, 127, 63, -7, -128, 127, -21, -128, 127, 106, -113, -128, 61, 127, -2, 22, 40, -128, 105, 127, 122, -128, -104, 43, 79, 46, 4, 105, 55, 127, -128, -128, 72, 127, 108, 63, -80, 31, 127, 56, 119, 127, 94, -128, 42, 127, -48, 127, -128, -26, 127, -128, -41, 127, -128, -128, -121, 127, 121, 57, 127, 25, -64, -39, 97, -128, 127, -128, 127, 29, -128, -73, 127, 127, -110, 35, -128, -128, 47, 127, 22, -43, 127, 74, -128, -128, 127, -128, 27, 89, -128, 116, -108, 127, -112, 97, 127, -128, 100, 44, -18, -125, 127, 127, -128, 115, 3, -128, -128, 127, -1, 29, 122, 127, -21, -34, 70, 127, 61, -128, -51, 127, -128, -128, 127, -128, 126, 127, -128, -99, 112, 18, -128, 25, -56, -128, -36, 127, -128, -128, 127, 127, -128, -39, 73, 98, -128, 127, 26, -128, 75, -18, 57, -46, -128, 127, 127, -58, 127, -62, -128, -128, -128, -75, -128, -79, 127, 127, 74, 127, -128, -128, -115, -128, -128, -128, -128, 127, -128, -128, 34, -125, -99, -76, -128, 127, 97, -38, -125, 127, -128, -128, -43, 100, -128, -119, 127, -6, 66, 127, 54, -128, -14, 70, -35, 92, 79, 90, 77, -128, 71, -128, -13, 102, 110, -128, 127, 127, -128, 2, 127, 127, -128, 25, 127, 127, -128, -128, -128, -36, 114, -9, -31, 127, -117, -128, 8, 127, 127, 6, 127, -128, 127, 127, -128, 106, 127, 100, -128, 127, 127, -128, -77, 127, -41, -128, 127, 127, -128, -29, -55, -100, 105, -128, -43, 127, -128, -128, 127, -128, -95, 53, 127, 68, 17, 9, -60, 127, -128, -15, 127, 127, -128, 43, 70, -128, -128, 127, 106, -128, 6, -128, -74, 32, -126, 127, 127, 10, -38, -128, -105, -128, -128, 62, 127, 127, -69, 127, 127, -128, 89, 127, -128, -128, 127, 85, -128, -20, 127, -69, 97, 127, 66, 127, 76, -128, -128, 127, 127, 14, -128, -1, 127, 127, -63, 36, 127, -21, -128, 127, 127, -44, 127, 82, -48, 52, 127, -128, -107, -66, 52, -47, 127, 41, -45, 78, 127, -68, -76, 127, 127, -81, -128, 64, -36, -128, -17, 127, 127, 12, 66, -128, 127, -55, -128, 81, 87, 7, -128, 110, -100, 92, -128, 57, -128, 127, 117, 18, 127, -108, -128, 43, 127, -128, -128, 127, 127, 127, -9, -76, 127, -11, -128, 127, 112, 127, 127, 82, 126, 127, 77, -83, -128, 12, -46, -128, 127, 31, 127, -28, -19, -104, -107, -128, -28, 127, 99, -128, -46, 7, -65, -128, 59, 20, -128, 127, 127, -44, 127, 82, -128, -22, 127, -11, -99, -128, 127, -38, -128, 127, -20, -128, -128, 127, 43, -128, -26, 48, -128, 76, 37, -128, -128, 127, -128, -128, -88, 14, 64, 127, 127, 71, 107, -128, 0, -30, 77, -128, -128, -128, -27, 127, -63, -128, 127, 126, -128, 127, 127, 22, -20, -128, -128, 127, -81, -114, 127, -107, -40, 70, 127, -128, 127, 49, 56, -97, -110, -89, -45, -128, 19, 22, 127, -128, -128, 80, -88, 23, -128, -54, -68, -29, -62, -128, 127, 127, -128, -128, 127, -128, -93, 31, 79, -128, -128, -22, 127, 127, 8, 120, -124, -128, -88, 127, -128, 127, 127, -128, 116, 127, -62, -32, -128, 12, 65, -28, -128, -128, 125, -18, -128, 38, -128, -120, -46, -34, -108, -6, 127, -54, -65, -77, 127, 127, -128, 61, 127, 21, -54, 127, 127, -119, -13, -99, -76, 0, -128, -43, -128, -128, -83, -26, 127, 127, 37, 127, 127, -128, 127, 69, -128, 127, 45, -128, 83, -128, 110, 23, -57, 28, -95, -109, 108, -42, 127, 116, 127, -128, 127, 127, -128, 127, -117, -128, 127, -111, -128, 127, 93, -128, -45, 14, -128, 127, 14, -128, 127, 92, -98, 127, -128, -128, -93, 127, 32, 0, 99, -20, -128, -10, 127, -128, -23, 127, -128, 3, -128, 127, -66, -128, 127, 52, 79, 127, -128, 127, 114, -128, -128, 127, -19, -128, 98, -87, 127, 127, -112, -115, -128, 127, -94, -128, 127, 29, -29, 124, -128, 83, -128, -128, 48, -125, -128, 127, -52, 70, 127, 39, -113, -128, 127, 17, -66, -108, -128, 59, 127, 13, 34, 127, 42, 127, 127, -12, 120, -8, 68, -104, -39, 127, -103, 60, -38, -128, 40, -128, -79, 127, -90, -46, 13, 127, -66, -100, -22, 127, 127, -128, 127, 35, 110, -7, 31, -128, -128, 127, 29, -128, -128, 127, -128, -128, 127, 3, -128, 127, -104, -125, 127, -128, -43, 10, -27, 5, 127, -128, 127, -128, -128, -71, 104, 127, 34, -14, -35, -128, 53, -85, 127, -128, 17, 127, -128, 127, -43, 124, 6, 71, -93, 126, -128, -38, 76, -32, 127, 127, -104, 127, -128, -47, 127, -47, 127, -13, -106, 127, 127, 10, 94, 127, -128, 46, 21, -29, -128, 45, 127, -128, -128, 127, -128, 127, 127, -128, 25, 127, -128, 10, 127, -128, 72, -128, -21, 92, -59, 60, 116, 127, -128, -97, -49, -128, 127, -113, -128, 127, 102, -128, -25, 100, 114, -128, 127, 127, 26, -128, -128, 127, -128, -128, 85, 80, -121, 127, 72, -128, 127, 63, 76, -128, 127, 120, -128, 127, 61, 11, 127, -128, 95, 104, -22, -128, 92, -128, -31, -31, 100, 48, -29, -81, 127, -128, 127, 127, 123, -11, 46, -6, -128, 48, 53, 48, 127, -128, 5, 27, 19, 127, -111, -128, 24, 96, -128, -128, 56, 82, 127, -114, -128, 127, 127, -128, -128, -128, 127, -128, -128, 119, 64, 0, -128, 127, -24, -54, -128, -128, 127, 70, 23, 127, 127, 119, 37, 127, -36, -3, 127, 23, -128, 113, 105, -7, 127, -128, 51, -36, -128, -128, 127, -128, -128, 127, 124, -128, 127, 127, -128, 127, 127, -116, 13, -128, -128, 127, -128, -128, 68, -22, -128, -128, 127, 104, -19, -128, 45, 127, 0, -128, -34, -71, -128, 127, 127, 127, 127, -128, -89, 127, 90, 127, 112, -128, -22, 127, -128, -128, -56, -26, 99, 3, 127, 14, -102, 127, 127, -128, -26, -24, 127, -128, 102, 127, -128, 113, 20, -128, 6, 127, 76, -128, 127, 127, -105, 53, 19, -128, -14, -128, 127, -48, 43, 127, 55, -91, 127, 20, 80, 127, -105, 14, -128, 92, 127, -55, 127, -79, -41, 127, 127, -52, -128, 127, 127, -128, 71, 105, -22, -97, -128, 127, -128, -128, 127, 71, -40, -71, 127, -54, 29, -128, -128, 59, -128, -128, 127, 116, -128, -78, -128, 127, -13, -87, 47, 90, -128, 109, 127, -128, 127, -111, -128, 127, -77, -102, -110, -5, -59, -128, 127, -124, 31, 127, -128, 127, 127, -126, -42, -128, -128, -128, -13, 127, 100, -30, 127, -128, -128, 38, 82, -19, -57, -48, -14, -128, -30, 66, -124, 127, 127, 35, 60, -128, -128, 127, -15, -128, 127, 91, -128, 1, 64, 127, 89, -122, -52, -128, -113, 19, -46, -38, 39, -128, 127, -26, -120, -120, 127, 7, 38, 127, 39, 0, -128, -128, 23, -128, 127, -36, -64, 127, -128, 127, -78, -91, 127, 127, -39, 127, -70, 127, -128, -58, 127, -128, -99, 127, 127, -94, 4, 127, 61, -128, 21, 104, -128, -128, -128, -104, 56, -89, -128, 122, 127, -128, -128, -103, -128, -59, -30, 10, -1, -96, 96, -76, -52, -128, 127, 127, -128, -45, 127, -106, -44, 86, 51, 127, -128, 127, 117, -128, -128, 127, 127, 46, -123, 107, 127, 5, -62, -128, 127, 8, -85, 48, -81, 127, 127, -58, 127, 56, -93, 127, 96, -128, 127, 127, -128, 127, 88, 11, -128, -49, 127, -31, -128, 127, -128, -76, 127, 57, -128, 127, -128, -128, 105, -68, -68, 127, 127, -128, 40, 52, -128, -128, -104, -4, 127, 19, -124, 71, 14, -128, -128, -70, -55, -114, 127, -15, 102, 93, -128, 120, -114, -128, 36, -102, -128, 77, 126, 127, -128, -128, -128, 40, -34, -128, -6, 127, 55, -8, -128, -128, 66, 63, 98, -128, 17, 49, -128, 127, 127, -128, -121, 41, 122, 127, 25, 73, -116, -128, 53, 75, 11, -28, 127, -85, -96, -116, -128, 127, -128, -128, 127, 127, 23, -128, 47, 127, -128, -128, 127, -70, 127, -128, -44, 45, -74, 127, -128, 45, 0, 127, 127, -44, 127, -32, -74, -66, -39, 56, -128, -12, -128, -128, -128, -36, 76, 127, 127, 113, -100, 116, 69, -128, -128, 61, -63, -128, -96, -128, -82, 127, -97, -128, 127, -5, -128, 19, 127, -109, -128, 53, 127, 88, -128, 127, 127, -115, -128, 127, -71, -74, 127, -119, 127, -128, -128, -21, -128, 37, 106, 0, 127, -128, -49, -128, 127, 127, 109, 70, 110, -128, -128, 4, -128, -15, 10, 119, 127, -128, 127, -26, -128, 127, -128, -128, 124, -128, 42, -128, -107, 32, -6, -41, -94, -128, 75, -128, -128, 73, 127, -128, -128, 127, 38, 127, -128, 26, 127, 4, -79, 34, 127, 71, -100, -120, 127, 127, -91, 127, 127, 5, 127, 127, -55, 2, -8, 110, 127, -128, -128, 45, 97, -128, 24, 127, -128, 91, -46, -28, 127, 127, -17, 9, 38, 111, -128, -128, -128, 70, 127, 127, 81, 121, -128, 127, 127, -46, -81, 22, 127, -128, -128, 127, 72, 98, 127, -128, -128, 127, 127, 0, 127, 66, -128, 24, 127, -128, -31, 127, -128, -128, -22, -26, -128, -31, -26, -128, 127, 127, -10, 0, -128, -5, 127, 109, -89, -96, -128, 39, 9, 127, 72, 90, 125, 6, -128, 89, 64, -128, -128, -128, 127, 68, -128, 127, 127, 21, 127, -128, 28, 13, 31, 127, -128, 58, -128, -128, -126, -55, 75, 1, -78, 66, -128, 127, -128, 22, -128, 108, -41, -128, 123, 7, -63, -47, 127, 12, -57, 127, -128, 35, 111, -128, -128, 52, -128, 127, 127, -99, -128, -79, -83, -26, 3, -128, 127, 15, -128, 127, 127, 28, 127, 127, 127, 127, -128, -128, 28, 30, -48, 56, 73, 127, 127, -128, 53, 127, -78, -61, -76, 39, -128, 72, -74, -69, 127, 39, -11, -18, -128, 113, -128, 86, -128, 98, -128, 127, 31, -97, 89, 40, -128, 127, -128, 90, 89, 127, -128, -34, 127, 6, 127, 127, -128, 127, 127, -128, 44, -128, -128, -108, -30, 5, 94, -41, 127, 127, -128, -128, 51, 127, -128, 120, 127, -128, -12, 27, 127, -128, -128, 127, -65, -128, 42, -128, 0, -128, -128, -128, 68, 127, 127, 123, 127, 127, -1, -94, -88, 127, 54, -109, 127, 127, -128, -128, -88, -90, -18, 127, 38, 6, 127, -128, -128, 127, -128, 127, 56, -128, -128, -128, -71, -65, 19, 26, -87, 64, 127, -128, 49, 88, -108, 105, -128, 66, 127, -112, 127, 72, -128, -17, -35, -128, -128, -128, -54, -73, -2, 127, 127, 59, 127, -128, 127, 72, 91, 57, -128, -128, -42, -65, -73, 0, -23, -128, 127, -128, -128, -128, 127, 127, -126, -128, 127, -128, -128, 127, 40, 102, 22, 61, -79, 117, 100, -128, -128, 38, -128, 112, 111, -128, -34, 127, 127, 82, -31, 102, 104, 127, -128, 13, 14, -128, 114, 126, -128, 100, 127, 127, -128, -74, -116, -103, -113, -128, 57, -128, -128, 127, 92, 61, -102, 108, 69, -78, 127, -128, 127, -97, -128, 127, -97, 127, 21, -128, 127, 59, -128, 127, -128, 70, -11, -128, 127, 127, -128, 70, 127, -128, -25, 127, 22, -128, 103, 93, -128, 127, 127, -120, -65, 65, 127, -128, -128, 76, 127, 127, -128, -5, 127, 127, -128, -128, 108, 127, -128, 127, -30, -65, 127, -128, 127, 127, -128, -128, -93, -128, -61, -57, 75, 127, -105, 127, 127, -128, -76, 127, 68, -128, 127, 127, -86, 108, -128, 39, 127, -90, -108, 127, 127, -35, -17, -44, 10, 74, 88, -75, 127, 3, -87, -85, -128, 127, -128, -21, 127, -128, -128, 127, 0, -128, 93, 12, -128, 127, -128, -128, 127, 18, -128, -128, 127, -79, -128, 98, 90, -126, 127, -128, -91, -98, 127, 7, -128, 126, 127, -36, 120, 127, -83, -29, 32, -77, -128, 72, -106, 127, 127, 127, 18, 111, -18, -113, 127, 66, -128, -122, 127, 127, -127, 56, -7, 127, 20, 121, -114, 127, -51, -30, 60, 40, 36, -128, 21, -128, -5, -92, 85, 110, -128, 75, -112, -128, -111, 97, 4, -70, -128, 127, -106, -11, 127, -128, 99, -4, 5, 127, -128, 25, -128, 127, -74, -128, 127, 127, -128, -55, 127, 127, -128, 9, -14, -128, 30, -54, -24, -128, 127, 93, -128, 47, 35, -128, 127, -26, -128, 127, 119, -128, 99, -128, -128, -69, -128, 37, 127, 45, 8, -12, -128, 108, -95, -128, -69, -128, 127, 69, 127, 22, 0, 60, -128, 127, 127, -93, 127, -34, 93, -128, 127, 127, -128, 87, -128, -123, 127, -119, -128, 127, -104, 22, 127, -128, 102, -29, 26, -128, 127, 51, -128, 127, 127, 60, 40, 1, 51, 127, -5, -128, -102, -38, -23, 100, -128, 107, 91, -128, 127, -128, -128, 127, -128, -128, 127, 127, 43, -128, 127, 127, -128, 65, 26, -46, 127, 106, 51, -128, -128, 125, -38, -128, 48, 127, -100, 127, -54, 89, -94, -44, -5, -128, -43, -128, 127, 127, 8, 59, -128, 119, -128, -128, 127, 127, -128, -128, -104, -128, -128, -12, -17, 28, 127, -70, -128, 127, 36, -128, -128, -128, 96, -128, -70, 127, 49, -128, 127, 4, -128, 117, -128, -128, 61, -128, -55, 126, 20, -128, -12, 127, -128, -82, 127, 127, -128, -47, 91, 127, -102, -128, -8, 127, -128, -86, 74, -126, -13, 62, 31, -107, 127, 127, -128, 47, 113, -128, -128, 127, -59, -128, -128, -36, 127, -62, -128, 127, 127, -128, -40, -4, -128, 44, 70, 96, -124, 127, -47, 127, -128, 127, 17, -128, -128, 127, -128, -128, 88, 127, 127, -128, 127, 127, -128, 80, 127, -126, -128, -128, 24, 39, 38, 116, 127, -128, -128, -128, 127, 14, 127, -11, -24, 127, -62, -128, 127, -48, -128, 127, 102, -115, 29, -41, 21, 127, -91, -14, 127, -128, -128, -123, -128, -30, -27, -128, 127, 127, -39, -128, -4, 127, 60, -128, 57, -128, -128, 38, 127, 37, -128, 127, 103, -104, 36, -20, -128, -78, -90, -125, 59, -128, -113, 8, -108, -102, 126, 82, 127, -128, 127, -38, -128, 127, -128, -125, 51, -128, 37, 56, 127, -128, 92, -30, -128, 127, -128, -128, 124, -128, -128, 63, 127, -128, -128, 127, 127, -126, -128, 127, -89, -128, 6, 41, 127, 127, -113, 39, 12, -128, -89, -128, 0, -128, 103, 127, -86, 120, 107, 127, 127, -54, -128, -18, 127, -54, -128, -128, -12, 76, 76, -51, 127, -56, -63, 127, 28, -116, -128, 20, 117, -5, -128, 79, 127, -96, -128, 127, 127, -128, 97, -128, -128, 127, 127, -47, 127, -68, -128, -128, 125, -128, -128, 74, -34, 77, -128, -64, 127, -128, 0, 127, 77, 9, 127, 42, 86, -128, 47, 127, -128, -66, 127, 69, -87, -109, -128, -27, -6, 127, 127, 127, 127, -86, -128, -51, -128, -128, 127, 127, -128, 60, 13, 4, -128, -6, -114, -128, 127, 61, -128, 127, 127, -128, -37, 127, 11, -128, 127, -128, -128, 125, -8, 127, -11, 69, 127, 95, -128, -89, 127, -128, -7, 127, -114, 127, 70, -1, 74, -128, -128, 127, -128, 5, 127, 82, 71, 127, -54, -39, -119, -128, 127, -1, -128, 24, -36, -66, -128, -128, 85, 127, 7, -128, 127, 127, -128, 127, -128, -128, 70, -128, -128, -128, 127, 7, -91, -128, 85, -17, 62, -128, -78, -128, -93, 126, 127, -49, 53, 54, 2, 127, -7, -100, -128, 56, -128, -128, 127, 127, -23, 127, 127, -128, -93, -94, -128, 127, -69, 4, 127, -128, -57, -85, -98, 3, 127, -128, -2, 127, 127, 127, -40, -128, -116, -78, -128, -15, 127, 100, -71, -107, -8, 127, -52, -128, 76, -128, -128, 127, 91, -104, -12, 127, -59, 24, -96, 4, -128, 127, -21, -128, -112, -10, 108, 127, -128, -128, -80, -41, 127, -128, -81, 127, -71, 119, 127, -128, -120, 127, -112, -128, -126, -128, -128, 127, -14, -128, 127, 127, -128, -60, -106, -128, 108, 127, 88, -123, -41, -42, -128, 127, -35, 6, 127, 47, -1, -128, -76, 127, -128, 71, 127, -128, 45, -128, 52, -128, -128, -128, -30, 26, -15, 0, 127, 104, 91, 76, 78, 127, 127, 127, -128, -20, 127, 38, 127, 127, -128, -128, -45, -128, -128, -111, -66, -107, 127, -82, -128, 127, 127, -17, 49, -128, -65, 127, -75, -128, 127, 59, 59, 71, 0, 127, -95, -46, -20, 96, -128, -95, -128, 83, -25, -43, -3, 82, 66, 127, -128, 127, 127, 127, 127, 127, 127, 123, 23, -128, -128, 97, -128, 127, 127, -128, -128, -121, 65, 35, -27, 111, 127, -113, -43, 127, -128, -44, 127, -128, -128, 127, -41, -128, 90, -46, -128, -100, -128, -116, -128, -46, -126, 13, -91, -117, -112, 127, -128, -128, 127, -128, -128, 127, 127, -110, -128, 127, 127, 0, 122, -27, -3, -38, 48, 127, 127, -8, -81, 39, 127, 38, 127, 74, -128, 107, 119, -128, 51, 69, 127, -116, 17, 127, 42, -128, 127, 127, -128, -73, -63, 127, -28, -128, 127, 127, 28, -6, 26, -2, -128, -22, -78, -128, -89, 81, -37, 17, -18, -128, -91, 127, -128, 21, 127, -47, 127, 106, -128, -65, 127, 92, 127, -128, 127, -40, -128, 127, -38, -72, 110, -128, 48, -128, 127, -29, -128, 115, 40, -128, 127, 127, 127, 127, 126, -32, -128, -52, 119, 0, -103, -128, 127, -4, 47, 127, 127, 103, -24, 88, 127, -9, -57, -128, -68, 127, -75, -128, -128, -28, 49, -47, -3, 34, 127, 29, 127, 53, -128, -128, 3, 127, -23, -128, 0, 127, -8, 52, 127, -102, -128, 127, 17, -128, 127, 127, -128, 127, 127, -128, 127, 116, -69, 127, -128, 127, 127, -128, -41, 127, -73, 127, -104, -128, 127, 80, 102, 11, 105, -87, 127, -128, -128, 127, -54, 0, 93, -128, 127, -128, -83, 127, 23, 71, 105, -44, -66, 20, 97, -128, -55, 127, -127, 78, 127, -128, 38, 127, 127, -128, 127, 98, -128, -125, -65, -35, 127, -77, 127, 127, 62, 127, -27, 56, 127, 37, -128, 104, -98, -128, 127, 22, 112, -128, 127, 127, -128, 127, 127, -128, 122, 89, -17, -128, -9, 47, -128, -128, 127, -128, 127, 127, -128, 24, 127, 127, -49, 95, 104, -128, 57, 123, -73, -103, -128, -128, 127, 127, -128, 26, 127, -46, -128, -88, 4, -96, -128, 32, 14, -128, -69, 127, 127, -72, 127, 126, 127, 64, -128, 127, 45, -128, 109, -38, -14, -128, 63, -24, 127, 127, 13, 96, 127, 127, -27, -47, -92, 30, -128, -128, -61, -128, -81, 46, 70, -128, -128, 77, -128, -128, 127, 127, -37, 127, 68, 79, -128, -128, 127, 76, -128, -128, -128, -66, 34, 76, -34, 127, -18, -128, 127, 127, -14, -4, 127, 27, -128, 107, 127, -35, 78, 11, -128, 41, -128, -128, -65, 127, 46, 127, 124, 56, -128, -44, -34, 127, -53, 100, 127, 36, 70, -36, -20, -5, -128, -87, -92, 127, -18, -30, 127, 127, -128, -125, 86, -128, 13, 127, 106, -21, 127, 112, -48, -128, 34, 10, -128, -2, 127, -128, -128, -87, 10, -128, 39, 59, -80, -128, -22, -128, 31, -109, 82, 127, -128, -128, -20, 48, -100, -128, -128, 127, -128, -128, 127, 56, 13, 127, 127, 19, 27, -128, 42, -104, -85, 127, -128, -128, 127, -57, -128, 127, 127, 99, 127, -128, -36, 76, -128, 69, 110, -128, 127, 127, 42, 127, -128, -128, -128, -123, 113, 127, 121, -128, -128, -42, -128, -128, -128, -91, -126, 92, -19, 127, 127, 127, -26, 6, -25, 127, -128, -58, 127, 127, -128, -128, -58, -127, -128, 47, 127, -79, -128, 127, -128, 31, 127, -128, 102, 127, -128, -31, 127, 39, -128, -99, 127, -128, -95, 127, 31, -128, 29, -128, 127, 32, -68, -75, -128, 127, -128, -128, 100, 69, 127, 127, 40, -128, -128, 127, 106, -35, -128, -59, 127, 90, 89, -42, 49, 127, 48, 113, -128, -128, 127, -128, -128, 127, 127, 127, 109, 102, -66, 127, 77, -128, 119, -96, 19, 127, -128, -99, -128, 76, -99, 9, 127, 49, -85, 0, -2, -75, -128, 127, 127, 78, 127, 127, -128, -128, 47, 54, 127, -116, -128, -79, -128, -115, -21, -6, -48, 127, 34, 70, 1, -86, -128, -98, 64, -40, -65, -42, -128, 127, -80, -9, 116, -128, -80, -19, 127, 127, -128, 13, 127, 127, 127, -128, 127, 127, -128, -11, 95, -32, -128, 127, -98, 28, -7, 127, 81, -103, 97, 127, 79, -128, -128, -128, 85, -128, -73, -86, -128, 127, 124, -128, 69, 127, -128, -98, -128, 124, -46, -128, 4, 127, -113, -34, 127, -37, -128, 127, -73, -128, 92, 127, 116, -51, -128, -128, -128, -128, -128, 123, 127, -128, -128, 127, 2, 18, 127, -128, 127, 127, -128, -126, -102, 127, -52, -128, 127, 72, 52, -128, 30, -7, 87, -128, 127, 127, -3, 72, 127, 127, -128, -5, 127, -108, -7, 127, -128, 127, 127, -108, 127, 127, 57, 127, -21, 62, -128, -128, -88, 122, -87, -83, 127, 40, 127, -128, 42, 127, 32, -128, -128, -119, -25, 124, -128, -69, 127, -124, -128, 127, 127, -47, -116, 27, -128, -128, -27, 69, 36, 127, -36, -128, 64, -88, -96, -41, -13, 32, -128, 127, 102, -73, 119, -128, -128, 90, 36, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -95, -116, 116, -128, -128, 28, -128, -128, -128, 87, 127, -31, -115, 114, -27, -72, -51, -41, -128, 127, 127, 46, -128, -17, 127, -128, -128, 127, -51, 9, -115, 127, 36, -71, 127, 44, -128, 127, 127, -128, -98, 127, -1, -128, 127, 127, -128, 27, 102, -128, 17, 127, -29, -32, 127, 127, -128, -17, 123, 127, -2, 127, -125, -128, 46, -120, -71, -11, 44, 127, -128, 75, 4, -128, -128, 2, 94, 127, -123, -128, 48, -128, -128, 127, 127, 42, 127, 54, -128, -128, -128, -128, -128, -124, 127, 127, -46, 127, -128, -128, 87, -28, -97, -128, 127, -128, -128, 127, -86, 127, -59, -13, 127, -128, -128, 127, -78, -49, 8, -128, 71, 127, -82, 4, 93, -71, 127, -128, 127, 127, -15, -128, -34, -59, -128, 127, -54, -128, 76, 127, 127, -107, -73, 127, -8, -128, 127, -120, -128, 127, 88, 112, 127, 119, 127, 127, 127, -128, -75, -128, -2, 100, 22, 127, -128, -73, 97, -128, -128, 47, -44, 127, -128, -128, 111, 115, 127, 36, 127, -20, -128, -74, 17, 122, -128, -128, 127, -128, -128, 127, 127, -24, -128, -28, -48, -128, -38, -34, 58, -53, 75, -128, -128, 98, -71, -128, 81, 127, -128, -128, 127, 27, -128, -93, -35, -80, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -15, 127, -3, -75, 127, -128, 127, 58, 127, -128, 127, 127, 79, -29, -86, 14, -28, -128, 127, 49, -128, 21, 116, -86, 127, -30, 127, 127, -42, -128, -66, 114, -36, 116, 127, -92, -128, 127, 127, -128, 127, 127, -128, 127, -15, -128, -128, -53, 19, -128, -38, 127, -116, -18, -69, -11, -128, -128, -128, -29, 127, 127, -128, -77, -41, -128, 127, 127, -78, -128, 127, -79, -6, -128, 45, 127, -128, 120, 19, -57, -128, 22, -121, 6, -57, 65, -128, 74, 47, -128, 51, 127, -128, 102, -128, -41, 127, -128, -128, 127, -128, -128, 127, -12, 60, -128, 6, 65, 127, 111, -91, -53, 127, 74, -128, -128, 127, -22, 127, 13, -128, -128, -128, -126, -128, -128, 115, 127, 127, 127, 127, -122, -128, -128, -128, -69, 127, 127, -128, 127, -128, -128, 73, -128, -47, 95, 127, 106, -128, -128, -37, -128, -89, -128, 38, 127, 91, 28, 127, -78, 14, -128, 116, 127, -128, -128, 127, 91, -128, -48, 127, 79, -51, -76, 127, -74, -93, 72, 127, -128, -128, 127, -17, 114, 127, 22, 127, 127, -25, -3, -128, -128, 127, -3, 98, 127, -82, -128, 127, -71, -128, -4, -41, 127, 127, -46, -19, 127, -128, -128, -128, -45, 109, 127, 125, 127, 127, 45, 126, 127, -40, -128, 127, 127, -128, 127, 127, -128, -128, 127, 92, -128, -3, 127, 72, 62, -59, -30, 117, -104, 127, 81, -128, 127, 127, -128, -15, 127, -111, -128, 127, 127, -128, -128, 111, -22, -15, 44, -86, 127, -128, -128, 127, 71, -128, -103, 127, -109, -121, 51, -128, -85, -52, -102, 127, 127, -128, 75, 49, 127, 15, -78, 14, 46, -8, -128, -128, 127, -128, -82, -128, -128, 19, 69, 127, 61, 127, -128, 25, 104, -128, -128, 127, 127, -22, 60, -128, 114, 127, 81, -52, 127, 127, -61, -128, 127, 79, -43, -128, 19, -62, -128, 127, 75, -128, -7, 127, 127, -70, 127, -63, -87, -108, 127, -51, -41, 108, -115, -128, 34, -128, -128, -24, 127, 36, -115, 37, -103, 115, 86, -128, 127, 127, 34, -111, -35, 127, 21, -128, 93, -14, -128, 127, -128, 124, 127, -126, -126, 43, -65, -87, 127, -128, -9, 0, -123, 34, -32, 43, -128, 82, 121, -128, 1, -35, 127, -59, -109, -128, 15, 60, 73, -128, -97, -128, 127, -128, -128, 89, -128, -46, 127, -113, -115, 127, -128, 107, 127, -128, -128, -46, -128, 25, 127, -91, -120, 71, -128, -128, 48, 1, 49, -108, 59, 127, -102, -128, -128, 58, -128, -128, 127, 127, -105, 127, 127, -128, 127, 127, -112, -21, 113, -81, -12, 127, -128, 69, 116, -128, -105, 120, -31, 127, -6, 127, -4, -128, -30, -110, -128, 127, -8, -105, -22, 127, 82, 127, -21, 127, -128, -128, 104, -96, -76, -128, 127, 54, -128, -128, 119, 127, 99, 47, 127, -128, -128, 127, 115, 40, 77, -128, -53, -19, -103, -128, 62, -52, -128, 127, -29, -128, 91, 15, -128, -128, 37, -42, 127, 31, -128, 57, 96, -128, -128, 127, -128, -128, 127, 127, 65, 82, 127, 45, -128, -128, 127, -25, -128, 60, 127, 127, -128, 127, 127, -21, -124, -128, -128, -82, 86, -128, 81, 127, 61, 127, 127, -98, 123, 18, -128, 60, 127, -88, -128, 127, -18, -54, -81, 127, -128, -79, -6, 127, -128, -128, 127, -128, -128, 47, 127, 127, -62, 54, -20, 127, -13, 88, 11, 127, 127, -128, -128, 127, -106, 127, 32, -128, 127, -128, -128, -48, -128, 53, -42, -128, 127, 127, -112, -123, -128, 127, 127, 114, -34, 102, -128, -128, 21, -128, -30, 127, -128, -90, 127, -128, -128, 127, 127, 44, 13, -31, 127, 127, -128, -44, 57, 74, 5, -126, -128, 127, 127, 17, 127, -45, -17, -88, -128, 127, 127, -128, 63, 127, -102, -128, 127, 125, 35, -116, 126, 30, 127, 119, -29, 127, 89, -128, 117, 127, 3, 127, 127, 0, -128, -128, 127, -20, -128, 127, 51, -80, -106, -128, 127, -128, -48, 127, 15, -128, 127, 127, -32, -128, 127, 10, 113, 127, -128, -23, 26, -128, -128, 127, -128, -128, 127, 127, 4, -128, 4, 127, -128, -128, 127, 59, -128, 39, 48, -128, -128, 75, -128, -128, 127, 127, -128, -128, 127, -8, 103, 127, -128, 8, 127, 4, -119, -72, -128, 127, -128, -128, 73, -128, 127, 127, -125, 127, 110, -58, 105, -46, -88, -45, 93, 127, -79, 127, -7, 3, -128, 68, 21, -128, -77, 127, 87, -109, -75, -128, 127, 127, 39, 127, 127, 36, -76, -128, -35, 72, -128, -128, 127, 127, -128, 34, 127, 127, 127, -70, -128, -128, 2, -80, -128, -128, 109, 66, 127, -66, 32, 127, 92, -128, -128, 81, 120, -128, -105, 127, -128, -128, 102, 123, -128, -128, 106, 5, -47, -58, 127, 36, -128, -18, 127, -39, -64, 4, -128, 127, -61, -85, 127, -128, 127, -74, -60, 124, -128, -128, 127, 59, -128, 19, 127, 127, -128, 127, 127, -128, -128, 127, 127, -19, 54, 127, -21, 72, 48, 86, -128, -44, 127, 61, 5, 127, -22, -128, -29, 109, -110, -128, 127, -103, -128, 127, -60, 55, 127, 23, -54, -128, -55, -39, -94, 23, -91, 107, 127, -108, 23, 127, 127, 127, -128, 36, 92, -128, 62, 127, -117, -96, 127, 19, -128, -128, -53, -60, 105, 122, -107, 54, 13, -128, -20, -117, 38, 48, -90, 127, -26, 10, 127, -128, -87, 127, 87, -128, 127, 127, -76, 78, -36, 17, -64, -128, 72, 127, -43, -128, 61, -80, -128, -128, 127, 127, -114, 98, 93, -113, -128, 127, 127, -128, -73, 127, 14, 81, -17, -72, -128, 127, 115, 127, -128, 127, 26, -128, 127, -128, -35, 127, -17, -69, -44, 125, -128, 15, 35, 68, -95, -123, -128, -10, -53, -42, 80, 127, -82, 48, -128, 63, -128, -128, 127, 127, 10, -73, 95, -128, -128, 127, -128, -128, 127, -61, -20, 127, -128, 71, 39, -110, 127, -128, -128, 127, 39, -128, 127, 127, -128, -68, -128, -128, 10, 86, 69, -13, 127, -64, -128, 127, 127, -68, -47, 127, 57, -128, -112, 127, -5, -128, 127, 127, -128, 39, 61, 127, -64, 83, -4, -43, 29, 127, -128, -52, -128, 98, 66, 125, -108, 77, -59, 127, -66, -42, -128, -9, 48, -3, 127, -128, 54, 90, 71, -56, -128, 127, -128, -128, 21, 61, 127, -128, -124, 127, 127, 124, 127, 45, -128, 58, 127, -128, -128, 127, 127, -57, -11, 127, -76, -128, 62, -115, -128, 127, 54, -128, 127, -10, 14, 86, 127, -75, -128, -98, 127, 98, 15, 8, -65, -128, 127, 127, -128, 58, 2, 119, -35, -128, -128, -66, -128, 127, -71, -128, 127, 115, -128, -65, 127, -128, -128, -85, -64, 85, -128, -128, 127, 18, -119, 127, -9, -128, 127, 4, -55, -90, -128, -128, 127, -128, -93, 127, -128, 127, 127, -128, 127, 127, 0, -128, -86, 127, -13, 28, -110, -66, -128, -94, -23, 109, 127, -58, 64, 9, -128, 52, -128, 127, 35, -128, -128, 70, -87, -85, 127, 62, -64, 127, -31, -22, -128, -1, -128, -128, 127, -128, -128, 127, 58, -128, -73, -73, -71, 127, -128, -127, 127, 114, -128, -49, 66, 127, 65, -128, -54, 127, 40, -128, -128, 127, 127, -113, -93, -11, 127, 61, -91, -119, -125, -70, 6, -46, 108, -77, -128, 127, 127, -122, -128, 71, 127, 60, 127, 127, -128, -24, 127, 53, 96, -128, -128, 21, -119, 127, 127, -128, 8, 127, -128, -128, 127, -69, 11, 72, 127, -128, 127, 127, -4, 39, -128, -128, -61, -128, 88, -119, -122, 127, 77, -128, -4, 13, -128, 127, 54, 87, -3, 91, 60, -128, 127, -59, 127, 8, 127, 5, -128, -27, 91, 49, -128, -69, 0, -128, 127, 81, 127, 29, -128, -128, 25, -2, -52, -128, 107, -20, -128, -25, 127, -4, -128, 127, 127, 6, -128, -92, 127, 127, -128, 14, 18, 9, 127, -128, -69, 127, -94, -20, 54, 38, -128, 127, 102, -128, 127, 127, -128, -30, 127, -128, -128, -97, 127, -128, -124, 127, -30, 14, -14, 17, 127, -128, 127, 127, -128, 127, 35, -128, 115, -128, 52, 127, -68, -117, 127, 127, -19, 77, -117, -128, -10, -128, 127, -108, -24, 127, -128, 48, -98, -58, 127, 127, 8, 66, 127, 127, -21, 111, -128, -126, 6, -128, 127, -83, 66, 7, -74, -70, 127, 127, -128, -23, 127, -106, -126, 127, 127, 58, -128, -27, -70, -120, 127, 87, 127, -91, 119, 127, 127, 18, -128, -128, 3, -87, -128, 127, 127, -128, -128, 102, -87, -128, 13, 127, -128, -128, -44, 127, 7, 57, 127, -74, 25, 127, -128, -112, 127, -128, -128, 127, 127, 61, 75, -119, 103, 127, -128, -83, -114, 2, -13, 127, -13, 76, 127, -128, 111, -28, 108, 25, -128, -128, 28, 46, 127, 53, 127, -128, -128, -21, -106, 61, -128, -128, 127, -128, -53, 127, -128, -128, 127, -128, -12, -28, 127, -12, -128, -43, -128, 81, -128, 127, 127, -23, 127, 46, -128, 127, 18, -128, 127, 127, -128, 127, 127, -128, -127, -1, 77, 127, -128, -128, 57, 127, -66, -24, 127, -25, -9, 127, -128, -14, 27, -61, -18, 127, 127, 45, 115, 48, 93, -128, -128, 127, -106, 102, 127, 41, -128, -128, 127, -128, -23, 26, -17, 74, 91, -128, 127, -128, -45, 54, 127, 43, 95, -128, -44, 127, 45, -61, 127, 36, -128, -125, -124, -4, -11, -119, -20, -59, 124, 127, 98, -110, 127, 127, -128, -11, 127, -128, -56, 127, -128, -71, -77, 68, 15, 127, -128, 127, -71, -75, 127, -122, -128, 127, 88, 127, -128, 127, 127, -128, -64, -60, 43, -8, 100, 127, -128, -128, 75, 127, -128, -17, 3, -128, 127, -128, 127, 127, -128, 127, -73, -128, 64, -128, 86, 35, -128, -128, 32, -128, -102, 127, 21, 51, -9, 70, -119, -128, 127, -128, -128, 63, 52, -19, 77, 127, -128, 90, -128, 127, -40, -128, 127, 112, -128, 127, -15, -30, 127, 35, -128, 28, 121, -20, 48, -128, -128, -89, 104, -80, -125, 127, -15, -65, 127, -109, 127, -128, 5, 127, 90, -128, -66, 127, 100, -128, 127, -128, -128, -128, -128, -117, 25, 127, 97, -27, 127, 127, 127, -128, 5, 23, -58, -128, -128, 46, -128, 127, 23, 127, 127, -128, 127, 127, 73, 37, -15, 127, -63, -128, 127, 127, -128, -7, -89, 127, -128, -128, 127, 121, 91, 127, -43, -29, 57, -125, -128, 127, -38, -128, -128, 26, -121, 127, 66, -128, 127, 127, -128, 27, 44, -128, 94, 127, -71, -97, 127, -113, -128, 127, 71, 111, -128, 127, 127, -128, 88, 127, -128, -128, -111, 43, -128, -128, 99, 37, -127, 127, 127, -128, 85, -116, -75, 8, -23, -128, 127, -9, 127, 90, 127, -128, -55, -40, 18, 93, -128, -103, -10, 127, -128, -34, 127, -61, 68, 68, -109, 127, 127, -128, -45, 127, 127, -128, 112, -75, -128, -128, 127, -25, -128, 110, 127, -87, -128, -19, -128, -128, 127, 127, -41, -19, 127, 127, -128, -9, 127, -128, -128, 78, 6, -128, -128, -65, 69, -126, -128, 127, -128, -128, 127, 127, 108, -100, 123, 127, 53, -128, -128, 40, -38, -95, -74, 68, 127, -128, -10, 86, 20, -128, 127, -128, 127, -128, -128, 46, -71, -112, -128, -27, -128, -10, -73, -64, 127, 127, -128, -10, -32, 122, 127, -28, 102, -99, -128, 127, -18, 70, 127, -128, -128, 112, -128, -104, 127, 95, -7, -98, 127, -103, -128, 47, 105, -128, -122, 127, -24, 60, -128, -108, 127, -75, 127, -103, -94, 83, 2, 32, -128, 2, 115, -128, -58, -59, 127, -88, -128, 127, 47, 77, -111, -128, 54, 48, 115, 127, 98, -26, -113, 127, -43, -128, 127, 127, -52, 38, 20, 126, -103, 127, 127, -87, 119, -128, 59, -89, -128, 127, -44, -128, -40, -7, -54, 23, 127, 127, -128, 127, 127, 48, -128, -109, 127, 56, -128, 78, 127, -128, 90, 127, -128, -128, 17, 127, -60, -128, 127, -70, 34, 127, -128, -128, 127, 87, -30, -127, 127, 127, -128, 127, 127, -128, 5, 127, -128, -64, 127, 127, 83, 72, -15, 98, -128, -128, -6, -104, 127, -128, -79, 127, -54, 127, 95, -117, 96, 127, -55, 127, 125, -128, -128, -69, 127, 52, -128, -43, 71, -128, -128, 124, 105, -30, -128, -82, 5, 127, 127, 32, 127, -128, -128, 112, 127, -24, -128, 51, 127, -83, 70, 9, 69, -128, 34, 127, -128, -5, -79, -128, 127, 127, -27, 34, 127, 127, -123, 57, 109, -39, -128, -128, -128, 127, 127, -45, 127, -27, -52, 127, 127, -128, 127, 127, 25, 127, -97, 59, -83, 127, 127, -128, 54, 127, 127, -25, 127, 7, -76, -128, -128, -128, 112, 127, -62, 53, 48, 9, 127, -108, 59, 127, 73, -128, 97, 127, -128, -128, 127, 78, -19, -120, 60, -128, 127, 127, -128, 47, 127, -128, -128, -23, 127, 82, -58, 127, 127, -117, 127, 127, 87, 73, -46, 86, 77, -128, 17, 34, -34, 127, -94, 104, 71, -128, -128, -128, -116, -92, 127, 127, 119, 127, -23, -8, 120, 127, -70, 93, -128, 20, 114, -128, -103, 127, 127, -128, 65, 127, -128, -81, 127, -128, -128, 127, -128, -128, 127, -128, -128, 85, -43, 127, 127, 10, 127, -25, 15, -73, 127, -107, 19, -128, 79, -18, -24, 86, 6, 127, 127, -128, 127, -36, 93, 127, -97, 91, 127, -51, 41, -73, -128, 127, -12, 24, -14, 127, -128, -128, 10, 127, 114, 30, 94, 127, 127, 91, 15, -128, -122, 127, -128, -66, 127, 7, 127, 34, -128, -97, -128, -128, 110, 86, 127, 127, -128, 127, 127, -128, 92, 127, -82, -128, -47, -10, 127, 127, -106, 21, 127, 127, -128, 38, -128, -128, 65, 32, -128, -65, 82, -128, 127, 127, 46, 127, -128, -91, 120, 22, -128, 102, -128, -122, 127, 127, 47, 93, 127, -128, -128, -11, -128, -128, -59, 127, 127, -128, 85, 77, -112, -128, 106, -128, -128, 127, 127, 57, 110, 127, -1, -128, -4, 6, -105, 127, -128, 59, -128, -45, 97, -128, -128, 77, 127, 127, -128, 127, 127, 44, -128, 3, -83, -64, 3, -128, 127, -125, -128, 127, -108, -128, 127, -3, 66, 127, -128, 14, 127, -69, -89, -128, 122, 80, -22, -128, 127, 127, -128, 127, 127, -94, 127, -128, -117, -49, -128, -14, 127, -79, -128, 127, 127, -128, 114, 29, -128, 127, 56, -128, 123, 127, -32, -115, 127, -76, -128, 127, 127, 40, -22, -128, -100, 127, -29, -128, 127, 127, -128, 80, 127, -128, -93, -56, 122, 77, -128, 90, 20, 127, -81, 127, 127, -21, -128, -45, -128, -128, -25, 127, 127, 64, 127, -128, 26, 97, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -14, -111, -52, -94, -94, 127, 127, -108, -112, 127, 42, -119, 127, 5, 127, -128, -38, 13, 96, 126, -66, 1, 127, -128, -90, 127, -127, -128, 57, 10, -128, -128, 127, -128, 127, 30, -128, 127, -62, -128, 127, 127, 89, 127, 13, 36, -128, -128, 30, 127, -36, -91, 127, 110, -34, -128, -19, 127, -128, 127, 127, -128, -3, -126, -128, 78, 2, 64, 73, -27, -108, 121, -128, 127, 23, -42, 125, -128, 127, 35, -128, 127, 127, -110, 127, -128, -128, 127, 127, 127, 127, 102, -128, -128, -14, 127, -128, -128, 127, -9, -43, 127, -128, 127, -128, -11, -47, -128, 127, 91, 99, 120, -128, -35, 127, 107, -86, -122, -10, 127, -128, -128, 127, 2, -37, 127, 127, 13, 51, -128, -128, 127, -5, -128, -7, 122, -128, -28, -20, -41, -128, -69, 46, 78, -28, 127, 127, -15, -117, -128, -128, -44, -80, -128, 65, -78, 6, 40, 127, 104, 8, 98, -128, 127, -99, 21, -83, -128, 83, -128, -17, 47, -128, -34, 127, -11, -37, 127, 127, -128, -95, 14, -128, -128, 103, 60, 127, -109, -113, -128, 8, -128, -35, 127, -72, -128, 47, 127, 97, -79, 127, 127, -36, -128, 109, -3, -128, 20, -122, -128, -94, 127, -98, -128, 127, -128, -128, 127, -100, -78, -119, 127, 127, -128, -128, -128, -46, -128, -59, 61, 127, -85, 127, -18, 109, 125, -128, -7, 127, 106, -59, 127, 127, -63, -128, -66, 127, -54, -128, -30, 64, -128, -125, 76, -18, -111, 127, -128, -128, 127, 31, -128, -13, -111, -128, 127, 23, 73, -22, -29, 13, -128, -113, 62, 28, 127, 26, -32, 12, 127, 58, -128, -82, -64, -128, 61, 98, -111, 80, 127, -128, -128, 52, 96, -124, -128, -128, 43, 31, 127, 127, -17, 75, -20, 48, -87, 127, -128, 93, 18, -128, -128, 127, -43, -128, 81, 102, -128, 76, 127, -51, 127, 127, -128, -103, 117, 127, -128, -38, 127, 89, -128, -42, 31, -128, -128, -108, -109, 127, 127, -39, 49, 4, -128, 48, -91, -128, -128, -128, 117, 127, 127, -41, 127, 127, -128, 43, 127, -128, -128, 127, -87, -115, 127, 127, -128, 14, -128, -128, 48, 51, -93, 0, 127, 66, 39, 30, -63, -58, 69, 103, -120, -35, -128, 127, 26, -44, 127, -128, -19, 6, -128, 23, -128, 127, -68, -128, 83, 110, 9, 42, 66, 127, -128, 127, 45, -128, 52, -9, 6, 125, 3, 24, -128, -128, 127, -128, -128, 127, -128, -107, -100, -128, -69, 127, 127, 90, 127, -128, -15, 127, -14, 127, 108, 31, -31, 127, -63, -128, 127, 127, -128, 127, 99, -128, 45, -126, 127, -128, 0, 95, -128, 127, -72, 65, -63, 58, 127, 12, 1, 127, -81, -2, 127, -52, 27, 127, 127, -128, 127, 127, 0, 41, -49, 81, 6, -91, -116, -98, -64, -128, 106, 68, -80, -128, -76, 28, 127, 48, -12, 85, -128, 103, 82, -128, -128, 127, 25, 127, -128, -21, 127, 113, -128, -90, -128, 24, 47, 127, -98, -13, 127, -63, -128, -44, 53, -128, -128, 104, -128, 45, 74, 105, -128, 63, -128, 42, -128, -128, 35, -8, 127, 127, -128, 49, 13, -62, 19, -128, 127, 127, -30, -128, 96, 127, -128, -128, 127, -128, -128, -128, -4, -126, 98, 127, 15, 32, 37, 127, -128, -128, 91, 127, 86, -128, 127, 71, -128, 127, -128, -63, 127, -44, -128, -51, -100, 25, -128, 74, 127, -46, 127, 20, 127, 61, 35, 5, 18, 127, 111, 34, -128, -72, 64, -100, -128, 127, -23, -107, 127, -128, -128, 1, -90, 24, -119, -128, 125, 127, 38, 42, -128, -128, 47, 35, -128, -128, 66, 127, -94, -128, 86, 127, 6, -128, -97, 127, 110, -128, -115, 127, 127, -128, -35, 127, 119, -128, -61, -128, 127, -23, -128, -115, 127, 120, 35, -128, -73, -128, 97, 127, -128, 7, 127, -55, 66, 127, -74, -86, -128, -128, -41, 127, 127, -128, 22, 127, -128, -128, 127, 127, -26, 74, -35, -128, 127, -128, -128, 127, -52, 10, 59, -128, -128, -78, -128, 112, 127, 44, -96, -83, 127, -28, -128, 127, 127, -128, 127, -128, 102, 127, -128, 15, 127, -96, -112, 127, 86, -104, 127, 127, -117, -128, -128, 127, -55, -128, 127, 104, 23, 58, 127, -128, -68, -66, 127, -39, 37, -127, 127, 14, -128, 127, -4, -128, 127, 97, 9, 127, -49, 39, -97, -128, -126, 127, -128, -128, 127, 80, 127, -128, 63, -107, -128, -76, 127, 63, -128, 127, 127, -86, -64, 127, -95, -125, 127, 127, -128, -91, 127, 44, -128, -128, -128, -91, 89, -61, -128, -128, 108, -128, -90, 127, -19, -128, 112, -106, -69, -127, -87, 127, -30, 52, -35, 11, -68, -61, 1, -128, -128, 127, 40, 127, 127, -83, 36, 81, 127, 127, -128, 109, 127, 87, 2, -128, -128, 127, 0, 116, -76, 127, 127, -128, 127, 127, -116, 127, 127, 127, 127, 111, -128, -128, -13, -128, -128, 127, -128, -76, 127, -128, -128, 127, -89, -128, -128, -35, 127, 127, 45, 68, 109, 127, -128, -128, -93, -128, -15, 127, 127, 127, -99, -121, 80, 63, -76, -39, 127, -128, 127, -128, -73, 127, -128, 9, 127, 103, 83, -128, -128, 43, -57, -128, -43, -74, -128, -34, -128, -128, 43, -38, 127, -35, 127, 109, -17, 35, 49, 127, -128, -110, 127, -128, -11, -66, -103, 127, -128, 43, 127, -128, -128, 127, 18, -128, -128, 127, 17, -128, 76, -121, -128, 89, 127, 75, 124, 127, 58, -107, 127, -39, -128, -103, 127, -20, -34, 127, 127, -123, 127, 4, -89, 71, -49, 127, -128, 31, 127, -128, -128, 127, -96, -128, -68, 127, 109, -44, -128, -3, -128, -80, 127, 70, 53, 127, 127, 35, -128, -5, 0, -128, 10, 127, 127, 85, 127, 39, -128, -128, 3, 9, -124, 127, 47, -128, -128, 127, 65, 127, -71, -111, 127, -18, -128, 127, 127, -128, 127, 121, -115, -73, 93, -99, -82, -19, -128, 127, -128, -110, 9, -128, 127, -128, -55, 127, -128, -91, 127, -128, 7, 127, -128, -46, 14, 127, -70, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -10, -128, 80, 37, -128, 127, -56, 127, -128, 127, -41, -128, -59, 81, -128, -103, 127, -128, 73, -10, -25, -128, -128, 127, 34, -128, 3, 127, -128, -128, 87, 127, -128, -95, 123, 127, -128, 127, 127, -39, -128, -128, 107, 127, -128, -64, 127, -128, -128, 127, 127, -128, -122, 127, 127, 127, 23, 127, -19, -128, 100, 47, -128, 127, -46, 127, 127, -55, -32, -128, -61, -114, -128, 82, 20, 72, 127, 127, 127, 127, -127, -128, -26, 13, -24, -98, -128, 127, 119, -128, 127, 127, -128, 127, 127, -128, 6, 127, -128, -81, -25, 127, 18, -128, 39, 127, 1, -115, 127, 127, -128, 44, 99, -82, 103, 127, -121, 10, -79, -128, -99, -128, 127, -114, 64, 11, -75, -128, 64, 73, -93, 22, 42, -128, -76, 127, -45, -128, 86, 127, -128, -128, 127, -6, -53, 127, -65, 127, 0, -128, -94, 127, 51, -128, 58, 127, -128, 38, -128, -120, 127, -41, -41, 114, -98, 127, 35, 116, 127, -97, -128, -128, -128, 127, 127, 127, -25, 120, 51, -123, -79, 92, 127, 127, 116, -21, -125, 116, 127, 105, 2, -27, 102, -128, -128, 127, -82, -128, 127, -4, -128, 88, 127, 127, -128, -99, 127, 119, -3, -128, 59, 68, -128, -128, 21, 37, 34, 127, -128, 45, 103, 127, 43, -128, -128, 127, -128, -128, 127, 121, -128, 127, 127, 34, -36, -69, -128, 121, -128, 124, -42, -91, 53, -128, 79, -128, -128, 127, 92, -128, -128, 127, -37, -128, -22, 127, -128, 117, -41, -91, -128, 127, -103, 121, 85, 83, 27, 127, 0, 60, 114, 127, 127, -23, 34, 98, -96, -128, -13, -128, 97, 127, -61, -128, 117, -72, 115, 127, -128, 127, 127, -83, 104, -34, -55, -128, -128, 127, 30, -46, 113, 113, -128, 127, -75, -128, 127, 53, -91, 127, 24, 127, 127, 79, -128, -128, 35, -46, -27, 64, 52, 127, 127, -128, -18, -32, -41, 98, 127, -128, -95, 4, -128, -128, -128, 95, 127, -128, -128, 127, -128, -128, -106, 127, 127, 41, 17, 3, -128, -128, -59, -40, 127, -2, 2, -128, -54, 127, 127, -128, 124, 127, -87, -128, 35, 127, -128, 21, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 108, -128, 65, 17, 127, 124, 18, 127, 91, 46, -128, -61, 127, 103, -15, 127, 75, -128, 17, -128, -73, 127, 125, 127, 49, 23, -128, -55, 103, -128, -128, 127, -27, -128, 127, -128, 32, -128, 127, 126, -28, 6, 74, -121, 127, -128, 127, 2, -128, 127, -85, -128, 127, 8, 43, 127, 127, -88, 22, -128, 89, -15, 127, 127, -128, 40, 60, -128, 127, -57, -128, 6, -60, 127, -56, -128, 18, -45, -128, 127, 127, -109, 14, 120, -128, 10, -3, -98, 127, 112, -102, 127, -66, -128, 127, 58, 127, 127, -26, -55, 107, 80, -128, 71, -128, -44, 127, 9, 18, 127, -128, -128, 127, 127, -58, 127, 127, 75, -121, 119, 97, 82, 12, -128, 41, -48, -91, 127, -94, -128, 127, 127, -128, -61, 112, 52, -128, -128, 127, -128, -128, 127, -21, 53, 127, -128, 64, -5, -128, 127, 127, -128, -128, 127, 72, -125, 97, 127, 55, -128, 127, 1, -128, 2, 127, 15, -128, 127, 68, -81, 127, -86, -8, -48, -127, -74, 15, -10, -128, 12, 127, 103, -128, 127, 36, -79, -128, -128, 127, -128, -68, 104, -128, 97, 111, 127, 127, 127, -69, -58, -55, -97, -89, 127, 20, 53, 106, 93, -96, 13, -128, 127, -128, -114, 127, -90, -128, 32, -11, -36, 127, -128, -12, 127, -128, 127, 127, -128, 23, 127, -128, 63, 127, -128, -125, 1, -128, -52, -128, -128, 127, 127, -30, 127, 127, -128, 127, 17, -128, -128, 61, -49, -128, -128, 127, -128, 0, 127, 90, 13, 60, 127, -128, -128, 127, -128, -2, -22, 48, 127, -128, -128, 56, 119, -97, -128, 127, 127, -128, 40, 99, -128, -128, 127, 45, 77, -128, -123, 127, -128, 43, 127, -96, -48, 10, 127, 93, 116, -128, -89, -15, -128, 127, 28, -128, 11, 119, 40, -26, 119, 95, 12, -1, -128, 36, -110, -49, 127, 127, 42, 100, 39, 114, -55, -128, 83, -23, 127, 82, 127, -45, 44, -128, -128, 127, -57, -47, 127, -128, -128, 127, 105, -11, 38, 127, -119, -128, 127, -57, -65, 127, 93, -128, 31, 127, -119, -51, 127, -37, -24, -114, 97, -1, -77, 127, -24, -35, 127, -113, -128, 108, 12, -128, -34, -24, 127, 31, 45, -128, 127, 127, -108, 90, 110, -128, -128, 23, -29, -128, -24, -46, 99, -96, -19, -31, 127, -128, -128, 126, -128, 42, 36, -108, -102, -60, 71, 127, 77, 127, -86, -64, -8, 39, -128, -57, 127, 127, 127, 24, 65, -64, -63, -128, -128, 127, 13, 127, -92, -128, -128, 127, -128, -128, 127, 127, 48, 127, -81, 127, 127, -128, 127, 127, -128, 40, 1, 112, 127, 127, -128, -128, -57, -71, 127, -128, 48, 106, -128, 127, -9, -128, -128, 127, -128, -128, -128, -86, -128, -51, 127, 116, 127, 10, -90, 14, 127, 49, -61, 127, -128, -17, 42, 21, 127, -44, -111, 127, 127, -37, 127, -128, -36, 127, 30, 91, 83, -128, 3, -74, 112, 127, -128, 31, -25, 127, -128, -128, 127, 127, -128, -128, 127, -128, -49, 127, -82, -41, 127, 127, -128, 60, 127, 27, -128, 28, 127, -112, 30, 107, 127, -30, -128, 127, 42, -128, 127, 76, -128, 21, 25, -63, -128, 127, 10, -55, 127, 127, 31, -97, 60, -128, -128, -128, 87, 127, 78, -128, 127, 127, -128, -128, 127, -128, -128, 127, 59, -128, -126, 123, 127, -128, 127, 127, -128, -28, -5, 127, 127, -128, -128, 64, 127, 127, -12, 127, 127, 65, -128, 27, 127, -36, -117, -128, 22, -122, -128, -128, 127, -128, -128, 127, -78, -128, 127, 127, -128, 48, 113, -128, -128, 36, -14, -124, 74, 66, -128, 108, -128, 52, 127, -48, -1, -25, 21, -128, 46, 127, 15, -94, 17, 123, -88, 102, 127, -97, 127, 127, 86, 127, -128, -128, 127, 127, -128, -128, 127, 127, -61, 60, 15, -15, -128, 82, -128, -128, 127, -51, 63, 103, 77, -38, -128, -128, 127, 127, 66, 127, 127, -83, -128, -128, 127, -64, -128, 108, -73, -128, -44, 127, 127, -128, -88, -60, -65, 4, -113, -128, 26, -122, 127, 127, 127, 22, -18, 13, 127, 12, -28, -59, 35, 127, -128, -7, -128, 32, 58, -34, -65, 75, 127, -128, 65, 127, -62, -87, -19, 39, 127, 127, -128, 127, 127, 72, 66, 127, 108, 127, 111, -128, -7, 63, -70, 127, -128, 127, 127, -11, 127, 127, -128, -11, 106, -4, -19, 47, 127, -128, 104, 127, -19, 123, 127, -128, 106, 69, -128, 28, 127, -128, 40, 127, -128, 127, 127, -128, 127, 127, -128, 127, -41, 127, 127, -54, 122, -90, 51, -128, -128, 127, 127, -128, -128, -103, -128, 127, 23, -128, -128, 127, 42, -36, -128, 127, -128, -128, 127, -27, -128, 127, 127, -128, -49, 127, -128, -128, 127, -55, 39, 6, -44, 21, -21, 127, -128, 127, 47, -11, -57, -128, 127, 127, -128, 24, 94, 127, 127, -128, 127, 127, -128, -128, -128, -73, 58, 30, 99, 113, -69, 127, 96, -42, 127, 108, -128, -95, -128, -36, 22, -128, 127, 127, -128, 57, 122, -110, -128, 43, 127, -52, -128, 127, 9, -128, 127, -128, 109, 127, -128, 127, 127, -128, 127, 125, -111, -128, 64, 127, -32, -128, 127, 127, -110, 127, -58, 102, 127, -128, -128, 127, -128, -128, 127, -82, -128, -72, -89, -128, -54, 99, 22, 61, 74, 127, 127, 43, 127, 72, -56, -9, -128, 127, -4, 127, -128, -86, 127, -128, -128, -128, 127, 58, 127, -34, 127, 76, -128, -35, 127, -65, 17, 127, 8, 127, -17, 119, -128, 100, 100, -128, -128, -108, 127, -128, -128, -40, 72, -54, -128, -37, 127, -128, -128, 127, -56, -52, 127, -128, 127, 14, 89, 10, -128, 127, 13, -62, 127, -128, 71, 127, 127, -32, 90, -128, -25, -26, -96, 127, -128, 66, -62, -116, 57, -128, -111, 127, 127, -95, 127, 94, -128, -88, 127, -51, -128, 78, -128, 127, 127, -128, 83, 21, -128, 53, 127, -37, -128, 127, 127, -128, 127, -85, -121, 6, -128, 23, 105, -114, -38, 127, -104, -128, -40, -95, 127, 127, 127, 127, 127, 63, 89, 0, -83, -38, -3, 127, -90, -128, -58, 127, 27, 93, -128, 64, 99, 127, -25, -41, 127, 126, 127, -128, 80, 104, -128, -128, 127, -119, 48, 72, -21, 127, 127, -128, 15, 123, 14, -89, -49, -3, 48, 76, -128, -128, 127, -43, -128, -77, 127, -115, -9, 127, -1, -128, 127, 39, -128, -128, 127, -128, -77, 127, -128, -112, 127, -100, -107, 29, 24, 9, 127, -43, -124, -128, 109, -128, -128, 127, -46, -128, 127, 127, -128, -18, -42, -127, 127, -37, -128, 127, 90, -1, -115, -113, 10, -128, 126, -13, 51, -128, -128, 127, -128, 13, 127, -128, 115, 127, -128, 21, 127, -73, 127, -128, -128, -128, 88, -37, -128, 112, -82, -128, 127, -8, -128, 42, 127, -44, -128, -119, 127, -128, -102, 127, -44, -128, 127, -128, -128, 127, -82, -70, 25, -128, -70, 77, -128, -3, 127, 127, -128, -76, 127, 127, -29, 60, -128, -15, -128, -128, 127, 127, 108, -128, -93, 21, -14, 127, 127, 89, 24, -122, 127, 61, -117, 127, 46, -58, -5, 127, -128, 127, 127, 127, -128, -123, -54, -128, -19, 127, -17, 35, 102, -128, -73, -128, -128, 127, 127, -126, 127, 127, -128, -119, 127, 110, -128, 127, 91, -128, -37, -46, -128, 127, 127, 106, 127, -128, -128, -76, 127, 71, -128, 104, -58, 127, 127, -115, 120, -53, 127, 48, 49, 53, -128, 91, 127, -128, 127, 127, -46, 127, 127, 127, -128, 26, -35, -128, -70, 127, 78, 10, 113, 127, -128, -128, 14, -128, 127, 127, -24, -53, -128, -108, 56, 73, -128, -128, -128, 27, -94, 79, 127, -38, 127, -1, -128, -128, -128, 127, 127, -27, -125, -128, 87, 85, -30, -128, 127, -105, -5, 127, -128, 24, 6, 94, 127, -128, 127, 127, -128, -128, 113, -128, -128, 127, 127, -128, -10, 127, 127, 112, -49, -21, 112, 89, -103, -92, -128, 35, -128, -47, -74, 70, 10, 94, 8, 127, -128, -6, -66, -128, 63, 34, 119, 77, -49, 127, -60, -128, 127, 127, -128, -77, 127, 46, -128, -3, -99, 29, 20, -96, 48, 127, -128, 8, 10, 127, -128, 41, 36, -128, 110, -128, -63, -128, -128, 127, 5, -128, 23, 127, -128, 127, 119, -128, -63, -128, 127, -35, -128, 127, 21, -128, -74, -32, 24, -48, -128, 127, 127, -39, 127, -128, -124, 53, 60, -115, -128, -128, -128, -9, 127, 127, -128, 127, 127, 0, 5, 127, 65, -128, -128, -27, -18, -111, 52, 45, 127, 127, 127, 116, -128, -128, 127, -96, 20, 6, -128, 116, -122, -18, 127, 127, 127, 65, -19, 34, 115, -36, -128, 119, 127, -128, 114, 2, 22, -128, 127, 53, -105, -128, 39, 87, -78, 127, 127, -128, -128, -88, -128, -128, 104, 127, 24, 24, -128, 127, 6, -128, -10, -10, -128, -38, -128, 127, 76, -87, 127, 127, -128, 127, 127, -128, 127, 127, -10, 49, -40, 127, -128, -128, 25, 105, 42, 52, 127, 124, -128, 28, 127, -128, 49, -13, -128, 2, 127, -128, -24, 127, 9, -128, -128, 1, -112, -128, -72, -56, 127, 127, 127, 127, 14, -96, -63, 47, -11, -128, 121, -21, -44, -128, -75, 127, -128, -1, 127, -81, -93, -128, -4, -128, -128, -8, 48, -61, -128, -76, 127, 97, -116, 127, 127, -128, -82, 115, -38, -128, 127, 127, -30, 127, -41, 36, 13, 102, -128, -128, 120, -128, -76, 127, 43, 41, 127, 119, 73, 46, -100, 9, 93, 127, -128, 127, 127, -128, -42, 127, -39, -128, 121, 127, -128, 26, -128, -128, 127, -4, 68, 127, -128, -113, -128, -91, -128, 127, -128, -128, 30, -128, 54, 127, -47, -100, 127, -35, -128, 99, 127, 49, -128, -49, 127, -54, -128, 36, -128, 31, -78, 127, -49, -128, -128, 127, -111, 53, 127, -76, 127, -128, 65, 127, -128, 127, 127, -128, -128, -128, -128, 100, -128, -128, -41, 0, 54, 108, -3, 127, 127, -128, 81, 127, 127, -128, -128, -116, -74, -128, -92, -128, 127, 127, -55, -128, -128, -43, -58, -128, 77, 15, -128, 127, -128, 17, -128, -42, 127, -128, -85, 127, 127, 9, 95, -13, -5, 127, -128, -128, 36, 19, -128, 127, 66, -128, -128, 127, -47, -128, -128, 31, -128, -128, -59, -13, -128, -89, 127, 48, -122, 0, 127, -26, -128, 127, 13, -128, -10, 28, -128, 127, -45, 35, 112, 114, 127, -128, -128, 44, 61, -128, -128, 127, -85, -10, 127, -25, -60, -128, 69, -7, 0, -119, -41, -78, 127, 35, -13, -114, -79, 127, -105, -128, -91, -128, -22, 127, 109, -128, 106, 127, -128, -128, 127, 127, -95, -45, 8, -32, 72, 127, -61, 53, -128, -128, -128, -128, -128, -128, -128, -128, -30, 127, 51, -21, 127, -40, 127, -76, -74, 127, 99, -128, 90, 127, -128, 70, -128, 100, 96, -128, -47, -128, 86, 8, -105, 127, 127, -128, 79, -46, 108, -128, -128, 124, -46, -13, 5, 19, -2, -128, 53, -12, -128, 76, -128, 127, 79, -128, -128, 117, -128, -32, 127, 89, 127, 68, -62, 98, -68, 8, -31, 125, -128, -125, 127, 12, -78, 127, 114, 127, -128, 13, 127, -128, 74, 113, -128, 5, 127, -128, -3, 127, -128, -34, 40, -59, 55, 127, -97, -128, 127, -128, -128, 127, -128, -128, 81, -113, -128, 94, -85, 127, 92, -54, 127, 20, 127, 37, -5, -128, 127, -128, -128, 127, 127, 17, 127, 127, -7, 60, -104, 127, 127, -128, -39, 0, -34, -47, 127, -128, 0, 127, 86, -128, -107, 127, 5, -80, 127, -128, -128, 127, -40, 127, -128, 127, 127, -73, 127, -93, 127, 127, -120, 17, -106, 127, 4, -128, -87, 127, -80, 127, -126, 12, 127, -13, 2, 127, -128, 48, 127, -128, -128, 127, -104, -57, 127, 78, -128, 127, 127, -128, 127, 127, -128, 127, -60, -128, 60, -128, 79, 58, -128, -55, 127, -128, -128, 127, -81, -128, 117, -83, 100, -29, -128, 127, 42, 127, 48, 44, -121, -128, 106, 82, 127, 24, 127, 127, 105, 103, 48, -17, 19, -128, -128, -128, -128, 36, -128, -128, 127, -6, -91, 127, 127, -128, 82, 96, -128, -128, 127, -128, -93, -19, 119, 59, -128, 127, 0, 15, 35, 127, -128, -128, 59, 56, 127, -105, -128, 127, 127, -128, 4, 127, 127, 25, -107, -128, -58, 127, 127, 26, -17, -128, 127, 44, -128, 112, -61, -128, 127, 117, -128, -128, 127, -113, 127, 127, -128, 127, 7, -72, -59, -128, 127, 127, -56, 127, 127, -1, -51, -58, 77, -9, -128, 48, -128, 127, 127, -70, -97, 127, 127, 91, -46, 59, -41, 39, 127, 29, 127, 46, -54, 127, 104, -128, 42, -7, -128, -123, -108, 127, -115, -128, 102, 66, 127, -128, -128, 127, -128, -64, 127, 127, -128, -115, 93, -59, 127, 11, 0, -75, 127, 24, -128, 85, -48, -128, -64, -31, -128, -113, -57, 127, 127, -4, -128, -68, -48, -59, 127, 0, -128, 127, -39, 27, 58, -128, 127, 127, -128, -128, 115, 127, -128, -68, -93, -77, 127, -128, -90, 72, -46, -31, 21, 127, 127, -128, 127, 127, -128, -103, -23, -97, 127, -128, -128, 75, -128, 17, 97, 127, -61, 21, 127, 127, -38, 127, -128, -75, 127, -128, -128, 127, -55, -128, 127, 120, -62, 44, -64, -128, -23, 127, -18, -128, -34, 127, -128, -128, 121, -115, 38, -128, 116, 61, -64, -128, 127, 127, 95, -128, 0, -128, 127, 36, -128, -123, 127, -59, 127, -128, -128, 65, -14, -128, -128, 127, 127, -128, 102, -128, -21, -128, 127, 52, 127, 127, -128, 95, 123, -87, -128, -85, 108, 66, -128, 62, 90, -128, -92, -128, 39, -26, 48, 127, 127, 80, 104, -128, -128, 127, 82, 75, -39, 51, -39, 127, -128, -128, 95, -128, -128, -10, -128, -123, 116, 51, -128, -128, 127, -128, -37, 127, 7, -54, 19, 79, 127, -83, 127, 127, -128, -70, -128, -35, 0, 127, 125, 0, -8, -8, -102, -128, 45, 127, 2, -128, -128, -2, -128, 0, -72, -47, 127, -128, 69, 127, -128, 127, 94, -4, 80, -128, 90, 127, -128, 127, 127, -45, 127, -28, 17, -75, -127, -7, -128, 127, -45, 7, -18, -35, 64, -128, 49, 93, -97, 127, 17, 53, -72, -45, -105, -70, 23, 76, 35, 126, -107, -128, 78, 127, -51, -128, 0, 52, -128, -80, 53, 127, 127, -128, 23, 127, 127, -128, 127, 127, -128, -18, 127, -117, -66, 91, 24, 127, -95, -81, 127, -8, -128, 56, 127, -32, 127, -128, 45, -128, -8, -5, 127, -28, 75, 127, -87, -128, -27, -128, 77, 127, -128, -128, 127, 62, -128, -64, -69, -38, -5, 127, 14, -60, -117, -128, -128, 4, -68, -11, -49, 121, 65, 127, 29, 127, -97, 127, 59, -128, 127, 127, -128, -128, 115, 127, 127, -76, 86, 63, 14, -128, 87, -20, -128, 127, -128, -116, 127, -128, -128, 127, 127, -128, 64, -109, 21, -64, 82, -128, 94, -111, 0, 127, 114, -128, 111, 104, -128, 127, 94, -128, 127, 123, -128, 127, 116, -128, 20, 127, -122, -128, -110, 65, 22, -27, 95, -128, -128, 109, -128, -68, -15, -128, 127, -92, -83, 127, -128, -114, 127, -31, -128, -128, 127, 109, -93, 127, 127, -128, 57, 127, -128, -128, -56, -94, -121, 51, 127, -14, 127, 127, -128, -3, -114, -128, 127, 127, -17, 127, -39, -128, 14, 125, -81, 127, 127, -128, 127, 127, -54, 21, -128, -128, 127, -65, -128, 127, 127, -128, -70, 127, -104, -128, -13, 127, -128, 127, 127, -128, 9, 127, 117, -128, -128, 127, 127, 82, 127, 127, 127, 127, -43, -60, 46, 92, -128, 20, 127, -128, -119, 19, -128, 85, -45, -128, 127, 127, -128, 65, 10, 127, 127, -128, 127, 127, -128, 27, 127, 38, 77, 127, 102, 127, -128, -128, -107, -60, -121, -128, 66, 127, -89, -128, 127, 24, -128, -128, 127, -103, -128, 127, 127, -128, 62, 127, 18, -62, -128, 127, 127, -15, -128, 88, 127, -68, 121, -42, -41, 127, 127, -76, 127, -13, -62, 17, 3, -128, 127, -128, -128, 61, 125, 127, -128, 91, 127, -128, -128, 15, -128, 88, -69, -111, 46, 81, 8, 7, -128, 127, -128, -128, 10, -70, -94, 59, -128, -35, 127, -128, -36, 127, 47, 127, 127, -128, -128, 57, -79, -98, 127, -36, -128, 127, 34, -128, -86, -7, -128, 127, 3, -128, 127, 127, 127, -128, 6, 1, -128, 98, 127, -128, 127, 26, -87, -128, -128, 127, 127, -60, 93, 127, -128, -128, 42, 127, -20, -128, -69, 127, -128, -128, -82, 127, -128, -128, 127, -46, 88, 127, -128, 127, 120, -128, -128, 127, 125, 127, -128, -8, 127, 96, -128, -11, 127, 95, -128, 127, 127, 1, 13, 127, -95, -128, 127, 22, -128, 127, 95, -128, -128, 127, -3, -128, -128, 90, 37, 15, 21, 127, 15, 18, 37, 127, 28, -34, -128, -110, 127, -128, 26, 127, -128, 35, 127, -128, -114, 127, -121, -42, 127, -128, -128, 127, -102, 6, 127, -128, 96, -128, -128, 127, 81, -94, 26, 127, 127, -128, 127, 127, -13, -128, -128, -59, 127, -128, -128, 23, -42, -128, 18, 76, 127, -11, -128, 1, 52, 127, 64, -128, 86, 127, -128, -128, 127, 103, -128, -128, -72, -8, -109, -128, -70, 31, -36, 103, -128, -20, 127, 103, 27, 127, 88, -2, 97, -128, -128, 127, -111, -2, 127, 64, 126, -79, -92, 95, 127, 70, 94, 127, 68, -31, -128, 89, -128, -128, 127, -128, 127, 127, -128, 100, 27, -128, -44, -128, -128, -30, 124, 127, 63, -128, -7, 127, 56, -128, -114, 5, -79, -128, 37, -128, -128, 127, 54, -128, -52, -28, -128, 41, -128, -90, 9, -128, -24, 35, 127, 127, 81, 127, 75, -128, 107, 7, -128, 116, -128, -15, 127, 57, -128, -22, 127, 127, -62, 127, 127, -128, -9, 127, -128, 127, 127, -72, 10, -128, -44, -71, -97, -128, 106, 127, -122, 124, -19, 127, -128, 127, 127, 87, -128, -121, 127, 114, -105, -128, -66, 107, -46, 108, 88, 102, 127, -128, -128, 44, -100, 110, 14, -128, -7, 127, -104, -65, 113, -128, 127, -124, 57, -64, 47, 127, -128, -128, -81, -128, -25, -128, 30, 127, 28, -65, 80, -128, 35, 127, -54, -128, 127, 127, 38, -95, -128, -20, -128, -128, 31, 59, 127, -128, 127, 62, -128, 80, 127, 12, -128, -128, 127, -37, -128, 124, -32, -128, 127, -30, -128, -29, 127, -37, 21, 127, -65, -99, 91, -53, -128, 127, 110, 20, -54, -128, -128, -128, -109, -128, -128, -47, 23, 127, -128, -128, 127, -57, 57, -76, -128, 127, -11, -128, -43, 30, -128, -65, 34, -112, -128, 127, 25, -128, 27, -128, -128, -80, -14, -128, -128, 81, 39, -49, -109, 127, 127, -128, 127, 9, -128, 127, -128, -128, 113, 127, -128, 91, 127, -128, -109, 93, 3, -13, -66, 127, 127, -14, 77, 77, -128, 127, 0, -128, 122, -128, -2, -128, -128, 127, 127, -128, -80, 122, 127, -128, 18, 78, -128, -128, 127, -23, -128, 127, -119, -128, 127, -128, 127, 127, -128, -128, 0, 127, -128, -128, 127, 127, -128, -31, 127, 99, -128, 1, 127, -80, -128, 127, 127, -110, -128, 127, -71, -128, 52, 127, 53, 31, 127, 127, -128, -76, -105, 9, 25, 127, 21, -128, 127, 127, -128, 127, 127, -40, 98, 21, 29, -128, 57, 4, 78, 127, -65, -41, 127, -128, -128, 127, 66, -128, 103, -26, 48, -68, -128, -7, -128, 127, -97, -63, 127, -86, -128, 51, -2, -128, 24, 127, -128, -128, 127, 66, -128, 127, 127, 37, 127, -56, -52, -128, 127, -128, -128, 52, -106, -128, -48, 127, 127, -128, 69, 127, 127, -128, 127, 127, 44, 127, 91, 127, 52, 99, 127, -128, -54, 46, -128, -128, 83, 20, -65, -128, -60, -128, 127, 127, 53, 105, -75, -128, -113, 127, 37, -128, -128, -112, 41, 59, -15, 85, 127, -128, -128, -102, -3, 55, -2, -97, 13, 127, 24, -128, 28, 127, 127, 95, 127, -12, 127, 127, -106, -37, -128, -128, -128, -128, -71, 25, -32, 127, 79, -128, 127, 49, -14, 127, 127, 127, 127, 38, 27, 127, 127, -128, 29, 126, -124, -122, -128, 127, 127, 127, 28, 127, -65, -10, 62, 37, -128, 109, -76, -128, 0, -128, 45, -37, 127, -27, -54, 127, -128, 127, 127, -128, 14, 35, 127, 52, -6, -37, 52, 0, -47, 127, -128, 127, 61, -128, -128, -88, 127, -128, -128, 102, 127, -128, -128, 98, 127, 99, -128, 31, 48, 36, -128, -128, 127, 80, -21, -128, -128, 127, -51, -128, 4, 105, -70, 127, 13, -41, -64, 127, -128, -128, 119, 127, 18, -58, 83, -2, -88, -121, 127, 97, -128, 127, 127, -128, -128, -104, -128, 13, -128, -69, 127, -122, -128, 127, -128, -128, 127, 18, 75, 22, -128, 127, 127, -128, 87, 1, -128, 127, -95, 23, 127, 96, -128, 127, 127, -128, -21, 127, 127, -128, -55, 127, 127, -128, 111, 15, 8, -72, 17, -128, 55, 64, 32, -71, -86, 127, -128, -128, -125, -13, 54, 60, 112, 127, 76, 5, -74, -128, -128, 127, -128, -128, 127, 89, -128, -128, -56, 65, 127, -128, -111, 127, -83, -128, 57, 44, -128, 127, 111, -128, 1, 24, 4, -17, -128, 127, -30, 125, -54, 36, 47, -128, 52, -128, -128, 127, 127, 127, -128, -73, 127, 127, -128, -93, 127, 127, -128, 127, 127, -128, -13, -113, 127, -15, 73, 127, -40, -128, 127, 86, -127, -27, -128, 57, 93, -128, 127, 127, -128, -128, -128, -128, 7, 127, -128, -65, 127, -128, -128, -66, -128, 42, -39, 22, 127, 57, 127, 127, 121, 14, 127, -82, -128, -128, -128, 39, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -5, 56, 127, 89, -128, -128, 127, -112, 127, -47, 91, 127, -128, -29, 127, -128, -128, 127, 37, -95, -116, -36, 127, -52, -128, 24, 66, 96, -128, -128, 127, -81, -124, 127, 127, -44, 127, 122, 127, -128, 40, -53, -128, -30, 127, 127, -128, -23, 127, 127, -128, -128, -12, -128, -128, 4, 127, -116, -128, 127, -60, -128, 44, -74, -128, 7, 112, 99, -8, 91, 127, -21, 127, 127, -128, -128, -9, -91, 59, 90, 96, -17, -128, 127, 11, 127, 85, -128, 39, 127, -128, 36, 75, 13, 127, -128, 32, 127, -125, 103, 127, -92, 127, 44, -128, -128, -128, -35, -102, -128, 127, 127, -128, -17, 127, 57, 12, 127, -128, -128, 127, -107, 42, 112, -128, 46, 105, 44, -20, 79, 127, -128, 110, 127, -128, -128, -71, 8, -116, 58, -128, -128, 123, -128, -128, 124, -6, -128, -58, 127, -128, -75, 127, -11, -128, 10, -69, 127, 9, -128, 110, 127, -25, -128, 127, 127, 116, 127, 127, -128, -92, 127, 18, 112, -128, -128, 127, 24, -128, 127, 127, -35, 40, -3, -58, -128, 3, -128, -76, 115, -128, -128, -14, 127, -128, -128, 127, -128, -88, 115, -53, -48, 127, -29, -128, -128, 127, -128, -128, 127, -99, 127, 71, -108, 127, -95, -128, -31, -128, -128, 6, 127, 105, 63, 127, 27, -128, -128, 127, -128, -128, 47, -128, 127, -46, -104, 127, -98, 127, 46, -128, 45, 127, 124, -128, -10, 127, 127, -127, -1, 127, -103, -51, 127, -9, -128, -128, 127, -128, -128, 110, 75, -128, -64, 127, -128, 45, 127, 47, -128, -128, 29, -9, 31, 127, 127, -20, 127, 127, -17, -73, 111, 32, -128, -102, -92, -128, 17, -39, 127, 119, 127, -108, -128, 127, 127, -63, -72, 127, -31, -128, 40, 88, 95, -29, 81, -128, 127, 41, -2, 127, -83, 77, -128, -99, 127, -82, 127, 127, 127, 127, -128, -128, 127, 106, -128, -128, 5, 127, -80, -128, 85, 127, 11, -128, 127, 127, -88, -53, 14, 105, 36, 127, -46, 127, -128, -97, 127, -26, -128, 127, 127, -128, -80, 127, 127, -128, 117, 127, 81, 9, -128, 127, 2, -128, 127, -128, -128, 127, -128, 80, 127, -116, 127, 127, 79, 31, 127, 98, -128, 127, 125, -128, 62, -46, -128, 127, 59, -128, -128, 127, -95, 94, 127, -128, -42, 19, -53, 51, 127, -128, 100, -128, -90, -128, -128, 24, 97, -18, -128, 127, -128, 100, 127, -128, 127, 127, -106, 127, -128, -128, -58, 97, 79, -115, 127, 127, -4, 127, 48, -17, -128, -44, -91, 54, -64, -94, 127, -128, 127, 127, 110, 126, 96, 127, 124, -86, -93, -99, -128, 31, 127, 127, -77, 127, -3, -128, -35, -123, 122, -119, -115, -20, -121, 89, -128, 86, -59, -128, 127, 4, -128, -2, 18, -102, 127, -128, -24, 127, 127, -128, 127, 25, -128, 127, -94, 51, -99, -128, 127, -21, -40, 52, 47, 26, -22, -74, -28, -128, 127, -71, -108, 127, 127, -128, 127, 127, -71, -105, -76, 127, 107, -128, -19, 45, 59, -102, -54, -128, 127, -56, -128, -117, 127, -128, -128, 127, 75, -128, -128, 127, 29, -75, 98, -18, -128, 127, -128, -128, 127, -75, -128, 127, -128, -125, -128, 96, 127, -88, -128, 127, -6, -71, 127, -128, 9, 127, -75, -128, 127, 127, 55, 127, 11, 127, 127, -106, 82, -128, -128, 25, -58, -128, 4, 127, -128, 127, 127, -128, 127, 80, -112, 79, -109, -128, 122, 127, -128, -64, 127, -64, 4, 127, 127, -128, -34, 127, -128, -128, -23, -122, -128, -57, 127, 87, -111, -128, 82, -128, -107, -128, -128, -104, 127, 127, 127, 127, 92, -128, -74, -66, 88, 88, -128, 127, 127, 55, 127, -17, 127, 127, -18, -38, 52, -112, -128, 85, 20, 127, 28, 127, -128, 127, 127, -31, 3, -22, -128, -128, 0, -113, -128, -76, 127, -100, -128, -40, 70, -128, -128, 103, -103, -128, -38, -40, -128, 127, 29, -128, -128, -44, -128, -119, 61, 20, 108, 92, 127, -39, 10, -128, 65, 127, 65, -128, 127, 127, -114, 59, 42, -128, 127, 127, 63, -45, -35, 117, 127, -69, -128, -128, -87, -128, 127, 100, -128, 127, 108, 127, 127, 0, -125, 127, 127, -128, -93, 64, 34, -25, 127, -128, 116, 95, 26, 0, 90, 127, 89, -128, 127, 55, -128, 127, -128, 127, 127, -83, 42, -128, 94, 127, 35, -53, -107, 44, -128, -128, 127, -104, 11, 127, 64, 127, -31, -122, 127, -128, -128, 127, 95, -111, -26, 127, -66, -128, 127, 103, -128, 73, 10, -128, 87, -128, 95, 126, -128, -103, 127, 27, -128, 25, 127, -128, 23, 127, 127, 22, 3, -128, -73, 127, -63, -128, 74, 127, 127, -89, 42, 127, 76, -128, 127, 100, 127, 87, 17, -6, 127, 127, -10, 127, -128, -128, -110, -128, -122, 127, -128, -113, 127, -128, -75, 127, 40, 115, -12, 63, -45, -22, -128, -100, 127, 127, 55, 46, -47, -128, 127, 127, -128, -14, 127, -43, 5, -128, -128, 127, 127, -128, -7, 127, -128, -128, 115, -48, -128, 127, 40, -23, 127, -124, -126, 114, -128, 127, 127, -70, 79, -17, -103, -27, 127, -88, 127, -128, -52, -37, 127, 127, -70, -58, 127, 32, -128, 127, 127, -128, 113, -32, -128, 127, -47, -128, -69, 127, -128, -85, 127, -128, 122, -10, 113, -128, -128, 127, 103, -112, 127, 127, -128, 127, 126, 34, 127, 114, -128, 92, 68, -46, 127, -60, 41, -121, 20, -128, -128, 96, 127, 35, -91, 3, -128, 127, -128, -128, 124, -11, -128, 20, -128, 53, 127, -128, 57, 95, -128, -54, 127, -45, -66, 62, 119, -128, -29, 127, -128, 103, 127, -128, -128, 127, -128, -128, 110, 79, 30, 127, 110, -128, -69, -128, 64, 79, -119, -15, 37, -128, -128, -42, -128, -65, 127, 42, -128, -27, -28, -5, 127, 74, 127, -128, -92, 47, -17, 46, -102, 23, -109, 20, -17, -128, -128, 127, -1, 26, 127, 70, 7, -128, 127, -110, -128, -41, 126, 47, -128, 127, 99, -121, -81, -128, 127, 127, -53, -61, -111, -56, -39, 127, -128, -68, 127, 64, -128, 127, 127, -13, -96, -128, 127, -79, -63, 126, -128, 127, 127, -94, 127, 120, 46, -12, -128, 127, -128, -128, 127, -128, -128, -128, 99, 54, -13, -81, 127, 80, 97, 127, -88, 127, -128, -128, 38, 81, 127, 31, 35, 28, 115, 127, -90, 127, -128, 2, 71, -128, -99, 127, 127, 127, -114, -68, -128, -27, 77, -53, 85, 127, -39, -128, 72, 96, -128, 127, 15, -128, 127, -8, -128, -54, -89, -128, -128, 127, -128, 119, 127, -128, 48, 127, 115, -128, -68, -85, 22, 53, -8, -9, 127, -128, -128, -77, -46, -98, -123, 127, 127, 127, -128, 62, 86, 127, 45, -128, -128, -128, 127, 127, -87, 34, 127, -98, -128, -97, -8, -53, -122, -95, -18, 127, -128, -128, 127, -99, -128, 127, 47, -128, 5, -55, -128, 127, -95, -20, 40, -71, -128, -128, 96, 127, 127, 127, 127, -71, 94, 127, -128, 25, -128, 71, 8, -128, 127, -19, -122, 124, -128, -54, -15, -95, 19, 127, -53, 59, 127, 8, -128, -106, 127, -128, -128, 127, 127, 127, -128, -128, 127, -95, -128, 127, 127, -100, 127, 108, -128, 127, 127, -102, 48, 127, -121, -128, -56, -72, -39, -128, -128, 127, -128, -128, 127, 83, -54, -128, -128, 127, -128, -59, -78, -128, 127, -128, -71, 127, -94, -21, -54, 124, -128, -128, 76, 51, 127, 1, -10, 127, 127, -128, 127, 35, -128, 127, -23, -128, 127, -74, -128, 127, 60, -128, 127, 127, 127, -128, -51, 91, 22, 97, 127, -128, -18, 127, -128, -128, 99, -128, 127, 1, 127, 127, -37, 45, -128, -42, 114, 120, 127, -128, 123, 127, 40, -108, -54, 127, 38, -75, 127, -128, 97, -10, 34, 127, -128, 69, 127, -128, -128, 73, -128, 36, 127, 127, -78, 127, 73, -128, -116, -8, -128, -128, 97, -128, -128, 6, -30, 127, -42, -128, 127, 47, -86, 120, 127, -128, 56, -30, -38, -128, 127, 127, 100, 127, 108, 46, -128, -128, -40, 11, 48, -116, 127, 127, -128, -128, 127, 127, -128, 74, 10, 127, 127, -4, -23, -128, 28, 127, 127, -123, 22, 127, 32, -90, 127, 19, 99, 5, 127, -128, 108, 70, -51, 43, -128, 4, 96, -128, 24, -38, -128, 127, -106, -128, -124, 8, -128, 30, 4, -102, 127, 19, 127, -45, -25, 127, -11, -128, 25, 127, -92, 127, 73, -128, -128, -54, -128, 26, 127, 127, 70, 127, -5, -123, 127, 127, -128, 116, 23, 32, 127, -43, -37, -128, -105, -128, -128, -128, -128, 18, 127, -15, -128, 64, 127, -4, -128, 52, 127, -121, -128, 78, -128, 72, -7, -58, 127, 46, 127, 1, -128, 127, 127, -39, 52, 99, -128, -128, 127, -30, -128, 127, 105, -128, 127, -128, -128, 17, -128, 127, 43, 63, 74, 18, 127, -128, 127, -128, -128, 127, -55, -77, 14, -128, -47, 127, -28, -128, 127, 127, -79, -22, 127, 127, 6, 127, 127, 19, 93, 112, -82, -36, 127, 94, -128, -128, 34, -128, -128, 127, -45, -79, -73, -41, 51, 65, -128, 127, 127, -128, 77, 127, 100, 25, 98, -97, -105, -128, 89, 127, 57, 57, 25, -24, -51, 127, -128, -128, -42, 17, -128, 127, -10, -128, 1, 127, -38, -128, 127, -128, -102, 127, -94, -128, -123, 43, -128, 83, -60, -128, 81, 77, 127, 120, 97, -128, -128, -128, -110, 82, 119, -85, -94, 122, -99, -128, 127, -13, 18, -11, -93, 127, -48, 21, 121, 69, -24, 127, -128, -128, -128, -65, -21, -128, -128, 24, 80, 18, -128, 127, 127, -128, 98, 127, -21, 59, 123, -34, 127, -114, -28, -128, -128, 127, 127, -128, 2, 115, -128, -128, -45, 110, 127, 48, 69, 127, -123, 127, -128, -128, -128, -6, 127, -96, -128, 127, -19, -128, -61, 93, 127, 111, -83, 127, 80, -128, -128, 127, 32, 109, 127, 127, -95, -128, 127, 69, -128, 127, 127, -128, 127, 127, -128, -128, -51, -128, -128, 70, 115, 127, 72, -128, 85, -29, -128, 127, 127, -128, 127, 127, -128, 107, 127, 24, -100, -128, -128, 127, 46, -128, 127, 127, -128, -83, 127, 127, -128, 127, 70, -128, 127, 6, -128, -111, 23, -89, -128, 119, 127, -128, 115, 127, -128, -119, 98, -128, 127, 54, -128, -79, 95, 77, 46, -128, 125, 127, -128, -66, 57, -73, -128, 127, -128, -128, 46, -128, 127, 127, -128, 127, 72, 79, 14, -128, 127, -58, -128, -128, 0, 58, -128, -128, 127, 46, -128, 127, 127, -18, -111, -128, 58, 127, -95, -128, 0, 4, 127, 105, -128, -80, 127, 127, -89, -128, 0, 127, -128, -128, 127, 82, -128, -128, 127, 62, -128, -68, 127, -63, -40, 9, -128, 127, -128, -59, 77, 9, -86, 87, 92, -128, 127, 127, -128, -39, -113, 127, -128, -128, 54, 127, -11, 53, 127, -128, -24, -112, 38, 127, 65, -28, -128, -128, -46, 42, 49, -114, 20, -76, 1, 39, -128, 127, 121, -61, 127, -128, 1, 82, 127, -128, -128, 45, -128, -128, 77, -128, -128, 66, -65, 13, 127, -88, 127, 127, -114, 127, 24, -128, 127, 48, -128, 127, 64, 127, 127, -128, 127, 127, -48, -31, -15, 127, 127, 127, -2, 127, 36, -128, -44, 18, -112, -114, -128, 83, -128, -45, 127, 80, 127, 127, 127, 99, 79, 31, -17, 81, -128, 17, 127, -128, 92, 127, -128, 127, 96, -128, -56, 127, -123, -58, 91, -111, 127, -128, -35, 127, -128, -92, -47, 127, 127, -128, -5, 127, -128, -128, 127, 127, -83, 127, 127, -128, -90, 127, -128, -128, -126, 127, -128, -128, 127, -18, -128, -1, 119, -128, 111, 127, -77, -124, -37, 127, 92, 69, 76, 127, 100, -128, 6, 127, -22, 127, 127, -108, 127, 127, -128, 127, 42, -64, 80, -128, 127, 127, -128, 127, 127, -20, 57, 89, -69, -128, -128, 127, 2, -128, 127, -69, -128, 99, -125, 127, -128, -128, 66, -127, 46, 127, -128, -128, 127, -128, -128, 127, -125, 97, 127, -128, 28, 75, -128, -128, 20, -128, 127, 36, -128, 20, -41, -128, 127, 24, 127, 81, -76, 123, 127, -128, -128, 127, -66, -128, 127, 62, 127, 26, -38, 43, -69, -128, 64, 127, 127, -104, 127, 127, 127, 104, 127, 88, -112, -27, 5, -128, 5, -128, 48, 127, -128, 127, 127, -128, -128, -128, 103, 127, -128, -128, 127, -6, -69, 127, -1, -80, -61, -128, -97, -86, 127, 87, -128, 127, -128, -68, 127, -128, -128, -5, 3, 113, -128, 79, 127, -11, 127, 15, -128, -19, 127, 56, 100, -128, -87, 115, 65, -128, -128, -122, -34, 127, 15, -128, 127, 49, -128, 41, 127, -128, -128, 85, 30, -128, -120, 103, -119, 53, 102, -125, 127, -128, -128, 13, -128, 56, 127, -56, -104, 127, 127, -75, -128, -36, 40, -128, -19, -66, 95, 38, 2, 127, 127, -20, 22, -128, -128, 127, 110, -128, -70, 127, 23, -128, 83, 68, -128, -128, -128, -75, -128, 66, 47, 78, 41, 127, -128, -128, 127, -100, -57, 127, 127, -128, -128, 74, 127, 13, -72, 127, 127, -128, 127, 46, -128, -89, 3, -65, 127, -128, -12, 127, -128, -128, 127, 127, -128, -36, 127, 127, -128, -72, -2, 127, -128, 102, 127, 14, -128, 4, -56, 30, -54, -23, -128, -128, 127, -128, -128, 127, 127, 127, -72, -100, -1, -69, 127, 106, -128, 127, -128, -128, 127, 29, 41, -77, -59, 127, 127, -98, -128, -83, -103, -128, 127, -79, -92, 87, 0, 127, -128, -128, 127, 127, -31, -128, -128, 100, -104, -111, 71, 127, -127, 127, 127, -128, -71, -128, -66, -86, -15, 127, -97, -1, -128, 82, 127, -128, -128, 45, 127, 65, -128, 115, -114, 113, 71, 83, -128, -14, -86, -128, -128, 75, 51, 90, -49, -128, 127, -128, 90, 127, -128, 127, 60, -108, -85, -128, 127, 71, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 24, 121, 119, -128, -128, -39, -128, -15, 127, 66, 81, 59, -128, -79, -128, -128, -15, 127, 127, 54, 72, 120, -128, -128, 127, 32, 66, 127, 123, 81, -128, -103, -128, -128, 47, 103, 127, 127, -128, 127, 127, -128, 91, 127, -123, 37, -44, -128, 21, -128, 69, -128, -10, -128, -128, 31, -82, -128, 127, 127, -79, -128, 88, -128, -128, 127, 127, 31, -40, 127, -128, -128, -100, 127, 40, -128, 81, -73, -128, -128, 91, 127, 62, -86, 110, 97, -128, 127, -128, -128, 127, 90, -38, -69, -128, 59, -128, -128, 127, -52, -125, 127, 127, -128, -94, 77, -128, -128, -28, 127, 119, -128, -128, 54, 31, 127, -128, -128, 127, -31, -107, 127, -128, -128, 30, -128, -120, -54, 5, -68, -128, 45, -76, -29, -41, 127, 127, -128, -6, 127, 123, 76, 29, -31, 127, -115, -120, 127, 127, -128, 127, 127, -55, -29, -128, 127, 18, -128, -32, 127, -128, -124, 127, -128, 53, 0, -128, 3, -128, 69, 103, 92, -102, 127, 127, 3, -128, -102, 120, -96, -128, -93, -128, 120, 107, -86, 51, 127, -128, -79, -90, 36, -128, 127, -128, -105, 127, 127, -128, 127, 127, -128, 0, 127, 127, -128, -69, 27, -128, -128, 127, 99, -27, 127, 73, 127, 127, 41, 6, -80, -128, -128, -128, -128, -79, -32, 80, 116, -51, -60, -128, 60, 127, -73, -128, 127, 71, -121, 127, 13, 127, -41, -128, 127, -40, -92, 127, -128, 127, 127, -128, -109, 9, -128, -128, 127, -36, -128, 127, 89, -128, 127, 38, -76, 127, -128, 127, -128, -128, 127, -128, -128, -22, 12, -128, -96, -128, 71, 103, 91, -128, -128, 127, -128, -128, 95, 74, 127, 127, 29, 103, 40, 87, -128, -68, 127, 60, -98, 127, -36, -114, 31, -128, 127, 127, 127, 105, 127, -58, -128, 57, 47, -17, -128, -11, -128, -128, 61, -14, -12, 43, 127, 127, -43, 127, -8, -103, -116, -11, -4, -128, 127, -124, -76, -39, 127, 127, -108, 36, 105, -92, -106, 127, -128, -128, -128, 127, 79, -128, -81, 127, 127, -128, -128, 127, 45, 35, 108, 127, 13, 68, 25, 127, -128, -128, 127, -128, -62, 87, -89, -53, 127, -128, 89, -128, -128, 127, 127, 127, -128, -66, 126, -128, -94, 23, -85, 100, 127, 127, 127, 46, -128, 58, 117, -128, 80, 127, -128, 127, 127, -128, 44, -128, -68, 98, -57, 127, 37, -128, -128, 73, 12, 127, -128, 83, -12, 127, 56, 127, -128, 127, 127, -128, 98, 127, 127, -86, 68, -11, -128, 127, -77, -117, 127, -52, 13, -128, 127, -34, -8, -46, 12, -107, -128, 127, 38, -128, -128, 127, 12, -128, -128, 127, -109, -100, 127, 15, -128, -53, -128, 127, 3, -128, 127, 127, -39, 127, 46, -32, 2, 127, -78, -90, 127, -128, -128, 92, 119, 81, -71, 19, -128, -127, -15, 127, 69, 17, 127, -128, 12, 39, -128, -128, 127, 17, 47, -5, -128, 86, 127, -128, -128, 109, -115, 123, 12, 43, -63, 127, -128, -128, -25, -22, -21, -128, -128, 47, -128, 93, 72, -21, 127, 14, -31, -128, 127, 4, 73, -59, -128, 127, 127, 76, 127, 9, -128, 108, 121, -111, 127, 127, 127, 109, 76, 116, 127, -128, -128, 127, -37, -20, 18, -128, -95, 8, 78, 127, -44, -128, -128, 41, 127, 127, -109, 14, 127, 127, -128, -128, -21, 127, 25, -128, 79, 127, -128, 25, -7, -111, 31, 127, 62, -128, 127, -38, -128, 127, -128, -56, 127, 110, -128, 127, 127, -128, 95, 127, -128, -61, 119, 122, -108, 72, 32, 104, -128, 73, 127, 114, -128, 127, 127, -65, -21, -9, 64, -128, -128, -19, 119, -128, -40, 127, -45, -100, 0, 127, 127, -128, 127, 81, -56, 127, -39, 26, -128, -72, 74, -111, 58, 127, 127, 38, -128, -98, 127, -86, 46, 127, -128, -128, -32, -128, -128, -128, 107, 108, -74, -120, 127, 38, 49, 127, -39, 127, -15, -128, 95, 37, -128, 66, 1, -90, 127, 26, -43, 76, -26, -128, 21, 127, -107, 38, 127, -49, -79, 127, 21, 127, 23, -27, -41, -12, -128, 127, -71, -128, -103, -128, -44, -37, 41, 99, -128, -128, 56, -12, -128, -128, 127, -128, -128, 127, -128, -128, 127, -111, -35, 127, 30, -62, 31, -128, -90, 127, -83, -15, 127, 117, 127, 87, -128, -128, -92, -128, 30, 117, -86, 127, 127, -57, 127, 43, 127, -128, -111, -77, -128, 127, 44, 127, -18, 82, 127, 6, -98, 127, 127, -77, 91, 76, -73, 127, 127, -128, -128, -24, -128, -128, -90, 30, 127, -34, -128, 81, 127, 47, -128, 127, -18, 61, 28, 111, 127, -75, -128, -30, 14, -128, -128, -31, -128, 127, 54, -100, -128, 127, -128, -128, -58, -128, 127, -2, -128, 127, 60, -117, 127, -120, 98, -128, -128, 127, 127, 73, -128, -60, 65, -128, 127, 95, 60, 127, -24, 100, 127, -66, -128, 127, -68, -88, 106, -128, 127, 68, -128, -31, 127, 2, -81, 127, 83, 127, -27, -128, 8, 70, -56, -107, 127, 37, 127, 127, 127, -23, -128, -128, 127, 77, -57, 55, 127, 88, 127, 54, 127, 127, -127, -128, -115, 29, 6, -128, 32, 89, 30, 58, 0, -128, -128, 127, -128, -11, 127, -128, 12, -82, 127, -111, -128, 18, 127, -128, 127, 127, -128, -128, 127, 25, 70, -128, 127, 127, -128, 0, -128, 127, 127, -90, 115, 127, -74, -128, 112, 127, -48, -30, 127, -116, 127, 127, -3, -127, 58, 127, -87, -128, 127, 127, -128, -128, 29, 127, -128, -128, 127, -19, 127, 98, -30, -49, 126, 124, -31, 6, 100, -37, 127, -128, -128, -128, 127, -128, -128, 89, -116, 127, 104, -128, 127, 127, -31, 127, -121, 77, 52, -128, 127, -128, -17, -128, 127, 127, -128, 18, 127, -37, 127, 73, -128, 24, 127, 77, -128, -60, 127, -88, -19, 127, -128, -128, -128, -128, 126, -69, -128, 54, 127, 127, -128, -1, 127, -5, -128, 127, -128, -128, 127, -1, 127, 8, -128, 127, 127, -63, 53, 127, -38, -128, 127, 127, -111, 66, 11, -82, -96, -128, -128, 61, 127, 127, 126, 127, -128, -128, -6, -128, 22, 45, -128, 127, -72, 124, 127, -128, 127, -44, -128, 71, 126, 127, 10, -128, 42, 127, -108, 75, 127, -37, 124, 127, 127, -128, -43, 127, -128, -128, 127, 100, -128, -128, 127, 37, -128, 86, 127, 5, -8, 127, 97, -128, 127, 127, -128, -128, -40, -125, -128, 127, 95, -128, -128, -74, -128, -91, 55, 127, -36, -25, 127, 22, 71, 104, -128, 90, -128, 127, 68, -128, 127, 127, -121, -60, 127, 113, -107, -69, 80, -95, -128, 127, -128, -112, -73, -19, 127, -128, 81, 127, -128, 127, 127, -128, -70, 96, -25, 127, -128, -2, 127, -47, -128, 127, -3, -128, 127, 127, -93, -128, 9, 127, -53, 127, -30, 108, -35, -65, 127, -128, 127, 127, 123, -128, -29, 127, 80, -128, 127, 13, -128, 127, 95, -128, 18, 127, -108, 127, -128, 45, 5, -128, -111, 127, -128, -128, 127, 6, -128, 127, 127, -128, 122, 94, 127, 57, -15, 25, 108, 49, -57, -128, -128, 127, 64, -49, 127, 127, -52, -128, 34, 127, -128, 11, -72, -49, -128, 127, 127, 127, -128, -48, -97, -12, 23, -128, -125, -99, 127, -128, -128, 127, -128, 99, 86, -108, -91, 94, 72, -35, -128, 17, -75, -125, -128, -46, 127, 24, 18, 127, 42, 127, 102, 83, -73, 127, -34, -68, 127, -70, -128, 75, 127, 14, -128, 4, 79, 127, -128, -128, 127, 127, -128, -128, 127, -128, -112, -128, 127, -26, 23, -92, 43, -128, -128, 71, 127, 109, -126, 53, -105, -46, -110, 127, 9, 61, 39, -3, 127, 127, -29, 6, -37, -85, -128, 0, -128, 55, 127, 2, -87, -117, -71, 32, 52, 14, 127, 1, -128, -14, 127, -89, 127, 1, 127, 127, -27, -128, -128, -128, -128, 3, -8, 127, 127, -128, 127, 76, -128, 127, 106, -128, -104, -128, 127, 0, 45, 54, 15, 86, -119, -86, 127, -128, -8, -57, -80, 23, -128, 31, 127, 127, -120, 127, 127, -128, 127, 62, -128, 106, -25, -128, -73, 49, 109, -128, 53, 127, -126, -128, -13, 46, 115, -75, -128, 127, 109, -128, -128, -45, 127, -128, -128, 127, 110, -128, -111, 127, -120, -128, 55, 97, -128, -106, 127, -85, 127, 127, -128, -48, 91, -128, -128, -128, 127, -128, -121, 127, 14, 4, 127, -128, 102, 105, -128, 127, 127, -108, -128, 2, 80, -128, 127, 127, -14, 127, 109, 127, 87, 127, 127, -42, 1, 127, -46, -128, 127, -128, -128, -102, -128, 79, -128, -128, 127, 127, -108, -128, -30, 127, -80, -128, 127, 127, -91, 116, 127, 127, -116, 127, 127, -46, 127, -128, 25, 127, -128, -124, -23, -128, -47, 108, -128, -54, 127, 6, 127, -128, -9, 127, -128, -128, 102, 127, -41, -14, 49, -128, -8, 80, 80, 127, -128, -2, 127, -82, -47, -81, -128, 127, -128, -106, 48, -128, -73, -128, 120, 127, 51, 79, 1, -128, -2, 127, 111, -28, 127, 4, 127, -2, -128, -34, -8, -128, 127, 42, -96, -114, 88, -128, -128, -48, 22, 13, 24, 127, -128, 127, -10, 18, 123, -127, -89, 43, -49, -15, -61, 127, 127, -128, 106, 62, -128, -11, 127, -128, -128, 127, 127, -52, -128, -54, 7, 116, -73, -49, -98, 127, 65, -104, -128, 127, 127, -123, -102, -98, -6, -61, 127, -40, 127, 127, -88, 127, 127, 5, 90, 127, 127, -1, -128, -128, 111, 127, 127, -128, -92, -51, -128, -58, -98, 13, 127, 22, 127, 55, -128, -21, -120, -128, 127, 14, 87, 127, -78, 127, -128, -90, 74, 2, 127, -87, 2, 35, -62, -128, 127, -128, -63, 100, -119, 78, 127, -87, -34, -32, -95, 117, -128, 127, 127, 63, -128, -128, -12, -113, -93, 127, 127, 15, 96, -45, -128, -128, -128, -128, 95, 127, 74, -128, 19, 127, -128, -128, 127, -96, -128, 127, 127, 56, 63, 89, -89, -2, 97, -128, 127, 59, 127, 127, 127, 38, -51, -70, 127, -128, -128, -64, 38, 103, -128, 121, 9, -128, 73, -128, -128, -40, 127, 127, 59, 54, 121, -128, -128, -128, -24, -128, -88, 105, 81, 92, 89, 110, 127, -128, -47, 127, -128, -128, 127, 127, -72, -41, 36, -128, 127, 89, 127, -15, -128, -105, 127, -128, -128, 17, -105, 30, 108, 127, -75, 32, 23, -19, -105, 127, -61, -79, 127, -125, -128, -40, 127, -128, -11, 17, -128, 127, -12, -86, -56, 127, -128, 127, 127, -128, -20, -66, -128, 127, -11, -128, -128, 88, 103, 91, -128, -9, 127, -128, -1, 19, -11, -128, -128, 127, -59, -52, -7, 127, -36, -104, 127, 127, -128, 43, -128, 127, -128, -98, 127, -103, -78, 127, -128, 98, 127, 127, -128, 11, 127, -128, 5, 127, -127, -74, 106, 99, -72, 127, 93, -128, 34, -128, -123, 86, 21, -128, 127, 127, -83, 107, -128, 127, 127, -128, -72, 127, -127, -68, 127, -128, -128, 66, -66, -128, 127, 55, -18, -86, -128, -13, -128, -128, 121, 127, 72, 41, -8, -128, -128, 127, -125, 2, 98, -128, -128, 127, 127, 127, 46, 27, -128, 110, 73, -128, -7, -18, -128, -128, -86, -128, 35, 78, 110, 127, -126, -36, -26, -128, 127, -128, -60, 127, 127, -128, -77, 18, 127, -128, 107, 127, -128, -99, 102, -29, -128, 20, -128, -128, 127, -106, -128, 20, 127, 127, 104, -114, -128, 127, 57, -128, -82, 20, 23, -52, 127, -128, -4, 127, 127, -88, 83, 48, 127, 127, -128, -128, -29, -122, -4, -48, 127, 27, 9, -128, -127, 127, -128, -120, -53, 115, 90, 55, -82, -11, -123, -128, 127, -128, -128, 60, 11, 32, 20, 127, -128, 56, 127, -128, -128, 1, 103, 113, -128, -128, -128, 127, 127, 127, 68, 124, -128, -127, 98, 11, 127, 64, -110, -128, -5, -17, -128, -128, 127, -128, -128, -74, -41, 127, 20, 19, -14, 119, 94, -74, 127, -128, -128, 35, 35, -128, -128, 123, -86, -128, 127, -32, -128, 64, -18, -128, -10, 127, -128, -128, -24, 21, -15, -128, 127, 93, 0, 127, 18, 127, -44, -128, -112, 58, -128, -128, -41, -128, 82, 21, -128, 127, 127, -4, -128, 48, 30, -128, 104, -128, 127, 127, 21, -60, -28, -25, -10, 83, 127, 34, 35, 127, -79, -128, 18, -128, -128, 127, -22, -24, 114, 127, 100, -103, -122, 127, 99, -63, 14, -41, 127, -128, -55, 112, -125, -36, 28, -128, 127, -127, 127, 120, 6, -128, -82, -40, -128, 127, -51, 97, 127, -57, 117, -128, -96, 127, -128, -128, 127, 127, -128, 76, 127, 9, 89, 127, -1, -85, 104, -110, -90, 100, -128, 127, -70, -128, 127, 127, -128, 113, 58, -94, 26, -53, -128, -128, 127, 21, -85, 127, -64, 82, 97, 73, -128, 38, -41, -128, 96, 88, -7, -128, 127, 127, 41, 98, -128, 25, 127, 110, -20, 127, -128, -128, 96, -102, -128, -104, 127, 113, -128, 3, 127, -89, -120, 127, 60, -95, -128, 57, -128, 127, -128, 40, 127, 71, -128, 127, -45, -128, -8, 37, -43, -128, 89, 70, -128, 127, 127, -128, 127, 95, -128, 49, 29, 59, -128, -7, 127, -26, 127, -128, -128, 127, -13, -128, 127, 25, -128, 70, 127, 127, -73, -56, -97, -128, -125, 69, -128, 15, 127, -69, 127, 127, -7, 45, -8, -13, -128, -128, 30, -128, -10, 88, -128, -128, 121, 26, 43, -79, 81, -128, 127, 62, -128, 127, 127, -128, 127, -42, 5, -15, -71, 20, 127, 22, 127, 8, 127, 127, -54, -76, 43, 100, 89, -5, 30, -128, -4, 127, 98, 22, -128, 127, 127, -94, -128, -62, 127, -116, -128, -128, 77, -128, 65, 124, -128, -88, 6, 94, 43, -128, 123, 127, -128, -119, 127, -128, -123, 127, -66, 45, 127, -54, -110, 127, 127, -128, 127, 34, -128, 91, -77, -128, -24, 8, 24, 127, 127, 127, 88, 17, -48, -55, -127, 41, 127, -128, 127, 127, 70, 10, -109, -65, 127, 1, 127, 58, 56, 29, -90, -120, -36, -128, 45, 12, 39, 127, -51, 127, -128, -61, -83, 48, 47, -86, 127, 127, 0, -128, 127, 127, -128, 4, -95, -128, 29, 42, -78, -36, 35, 61, 127, -128, 91, 127, -128, -128, -128, 4, 42, 127, 14, -79, 17, 127, -81, -128, 127, 127, -128, -90, 127, -10, -128, -3, -13, 127, -128, -128, 127, -128, -63, 127, -128, 127, 127, -128, 127, 70, -108, 127, -128, -128, 55, -126, -98, 127, 127, 78, 127, 127, -53, 22, 78, -128, 78, -20, -128, 127, -128, -17, 127, -128, 62, 127, -128, -54, 99, -60, -128, 123, -128, 112, 127, 127, -128, -51, -9, -128, -114, 127, -121, -128, 54, -14, -128, 127, 126, -128, 127, 127, -128, -47, -60, 127, -77, -128, 83, -128, -73, 109, 127, -76, 127, 110, 127, 127, 127, 78, 78, -128, 8, 29, 80, -26, 79, -128, -45, 127, -55, 113, -128, -99, -128, -5, 32, -128, -115, 120, -128, 30, -111, -122, 1, 23, 8, 127, 127, -128, 124, -35, -38, -1, 123, 116, -128, 111, 122, 127, -86, 69, -48, 119, -128, -128, 127, -128, 115, 127, -48, 105, 53, -128, -119, 127, -128, -94, 127, 127, -128, -30, -88, -128, -2, 127, 127, 127, 127, 123, -128, -72, 127, -92, 0, -46, -128, 95, -91, 115, 127, -95, -128, -42, 127, -34, -11, 127, -122, -19, -22, 8, 127, -128, 127, 127, -128, -2, 127, 26, -128, -110, 127, 127, -128, 12, -12, -128, 127, -128, -128, 127, 127, 127, 106, -123, 127, 29, -128, 123, -103, -128, -125, 127, 127, -8, 127, 54, -128, 60, -113, -93, 127, -3, -128, -96, -128, -63, -128, 127, 127, -128, 127, 127, -128, 60, 59, -128, -108, -128, 127, -128, -128, 127, -128, -23, 105, 127, 127, -128, 39, 34, -42, -9, -128, 127, -128, 81, -30, 127, 13, 127, -19, 36, -128, -128, 93, -6, -128, -128, 127, 127, 74, 11, 7, -128, 127, 93, -87, -15, 127, 127, -128, -28, 127, -37, 127, -115, -59, -32, -42, 127, -128, -111, 98, -128, 127, 127, -128, -66, 127, 127, -128, 127, 88, 127, -128, -96, 10, 125, -128, -128, 127, -128, -128, -29, 61, -128, -8, 108, -128, -30, 127, -17, 127, -56, -124, 40, -60, 25, 1, -69, 127, 127, -128, 73, 1, 117, 127, 120, 4, 127, 127, -128, -128, 108, -86, -38, -77, 111, -59, 127, -128, -32, -94, 127, 31, 21, 127, -95, 27, -110, 61, 127, 127, 4, -22, -128, 64, 34, 82, -128, -3, -56, -128, 127, 127, -46, 55, 127, -128, -128, 127, 127, -128, 44, 127, -128, -128, -128, 90, 0, -125, 127, 35, -128, 95, 127, -18, 110, -73, -120, 127, 98, 23, -128, 79, 127, -128, -128, 127, 51, -128, 125, 127, -104, -128, 54, -128, 47, -128, -128, 127, -108, 127, 127, -128, -128, 57, 0, -111, 69, 112, -58, 127, -128, -98, 127, -128, 127, 38, -19, -128, -110, 126, 122, -128, 106, 127, -128, 93, 127, -113, -128, -121, 37, -107, 88, -128, 18, 127, -65, 127, 127, -128, -55, 127, 102, -128, 127, 127, 54, -103, -31, -128, -128, -122, 127, -128, -128, 127, -128, -128, 127, 54, -18, 73, 127, 127, 38, 42, -78, 127, 127, -128, -127, 0, 106, 83, 69, -128, -43, 19, -128, -28, -128, 66, 127, -128, 127, 124, -128, 127, 43, 68, -128, 127, 98, 127, 127, 49, 127, -22, -128, -79, 103, -128, -128, -22, -128, -128, -128, -6, 127, 127, -24, -113, 57, 127, -128, -21, 127, -128, 127, -56, 3, 127, 127, -128, 127, 3, -128, 116, 127, -24, 127, -22, 64, 76, -128, 116, 127, -128, 45, 105, -59, 127, 127, 127, 75, 5, -128, -128, 127, 79, -128, -128, 127, 127, 127, 61, -76, -25, 39, -106, 97, -128, 127, -98, -90, -128, -57, -128, 3, 11, 127, 62, -128, -56, -12, 127, 127, -65, 70, 127, -2, -128, -17, 127, 127, -93, 127, 127, -128, -128, -62, 127, -52, -128, 30, -70, -63, 127, 102, -128, 127, -128, -128, 127, -55, -128, -117, 127, -128, -62, 127, 93, -32, -56, -98, -26, -85, 26, -128, 127, 48, -119, -76, 112, -80, -128, 127, -128, -128, 20, -59, -128, -128, -128, 11, 39, 107, 35, -109, 127, 46, 23, 127, -128, 82, 1, -128, -57, 127, -87, -109, 127, 14, 55, -128, 22, -49, -128, 4, -111, -69, 114, 24, -68, 127, -128, 28, 56, 114, -128, 108, 127, -128, -12, 127, 127, -128, -128, -55, -10, -62, 21, -77, 127, 127, -54, -22, -128, -107, -36, -122, -128, 113, -128, -81, 127, -128, -128, 127, -70, 24, 127, -128, -128, -56, 62, -128, -128, 56, -128, 127, -54, 127, 127, -55, 109, 48, -41, -128, -32, 97, -120, -88, 127, -128, 127, -63, -80, 121, -128, 127, 32, 8, -75, 127, 88, -128, 127, 78, -128, -23, 127, -114, 74, 127, -128, 127, 29, -128, -128, 127, 55, 127, 127, 66, 42, -120, 127, 127, -128, 127, -25, -128, 127, 127, -128, 127, 120, -128, 127, 127, -128, -92, 39, -113, -28, 127, -128, -128, 127, 127, -75, 125, -59, -128, -128, 127, -32, -128, 127, 13, -54, 127, 19, -128, 127, 9, -128, 127, -128, -13, -39, 127, 127, -47, 74, -47, 122, 127, -121, -128, 70, -65, -128, -35, 66, 127, 115, -128, -21, -49, -128, -121, 92, -14, -94, 127, -128, -112, 127, -9, -128, -19, 24, 127, 44, 127, -128, 74, -77, -128, 127, -128, -128, 127, -128, 124, -15, -6, -128, 79, 98, 126, -8, 127, -128, 53, 127, 127, -128, 58, -81, 108, 39, -128, -11, -64, -27, 127, 2, -95, -97, 105, 36, -65, 127, -48, -128, 37, 6, 127, 127, 23, 49, -102, 127, 91, -128, 127, 127, -128, 127, 70, -128, -128, -128, 20, 68, -15, 110, 45, -121, 127, -128, -91, 127, -10, 127, -117, 127, 27, -128, -90, -85, 127, 127, -90, -34, 5, -82, -15, -123, 108, -24, 127, -128, -88, 127, -120, -128, -12, 37, 127, 79, 87, -128, -3, 127, 31, 127, -128, -58, -128, -38, 121, 127, 89, 127, 127, -128, -128, 127, 127, -128, -19, 61, -128, -128, -12, -128, 127, 65, 23, 127, -72, 127, -128, 105, 127, -128, -128, 87, 121, 113, 25, 127, 127, -128, -97, 127, -13, 127, -23, -124, 127, -128, -128, 54, 71, -51, -128, 78, 127, -128, -128, 44, 127, -82, -30, 127, 127, 43, 127, -128, 32, -49, -128, 127, 91, 127, -30, 127, 45, -128, -62, -128, 12, 127, 127, 127, -27, -128, -95, 94, 26, 39, 127, 127, 0, 108, -105, -64, -128, -128, -15, 18, -128, -85, 127, -128, -128, 127, -126, -40, -100, 127, 127, 102, 127, -128, -96, 127, -128, 5, 122, -128, 41, 127, 127, -128, -24, -17, -77, 127, 127, 127, 127, 127, 65, -128, -56, 127, 36, 127, -128, -128, 127, -86, 63, 127, -128, 110, 1, -128, 127, -128, -128, 25, 127, -128, 21, 65, -128, 127, -14, -128, 103, 127, -83, -128, 109, 127, 44, -123, 88, -128, -96, -128, 127, 88, -128, 97, 127, -128, -128, 127, 0, 127, 127, -128, 127, 127, -128, 105, 127, -128, 127, 73, -128, -65, -128, -128, -128, -96, 103, -58, 66, 127, -128, -128, -13, -60, -128, -128, -34, 122, 127, -56, -128, -13, 26, 85, 47, -128, 26, 127, 49, -128, 99, 127, -5, -18, 127, -27, 99, 77, -8, 127, -128, -128, 45, 127, 94, -128, 12, 127, 106, 22, -128, -52, -128, -128, -21, -128, -68, 25, -29, 110, 127, -128, 127, 127, -121, 127, -128, -128, 14, 64, -92, -38, -125, 127, -128, 0, -102, -128, 108, 127, 127, -34, -72, -113, -25, -128, -127, -83, 127, -30, -5, -37, -128, -114, 37, -128, 58, 127, -128, 127, 127, -128, -128, 64, 86, -23, 76, 127, 54, 127, -128, 42, -107, -128, 127, -7, -128, 127, -46, -128, 127, 73, 127, -128, -56, 52, 99, -128, 69, 127, -34, 11, -128, -128, -2, -128, -69, -62, 97, 127, 127, 89, 127, 3, 127, 126, -128, 127, 36, -128, 127, 127, -128, -128, 37, -128, 11, 127, -19, 24, 127, 115, -128, -8, 127, 54, -128, -76, -54, -128, -41, -10, 62, -128, -128, -44, -128, 127, 46, -64, 116, -128, -1, 127, -79, -128, 127, 3, -114, 127, -102, 127, 127, -24, -128, 21, 17, -128, -71, 127, -128, 89, 127, 127, 127, 37, 127, -13, -128, -128, 127, 127, -45, -12, 127, 127, -128, -38, -65, -128, 127, 127, -128, 2, -8, -128, -128, -128, 32, 90, 102, -65, -62, 127, 41, -128, 127, 28, -128, 127, 59, 127, 126, -3, -128, -128, -25, -128, -128, 127, 127, 34, -128, -74, 127, -8, 1, 127, 60, -55, -53, -128, 127, -128, -123, -128, -27, 116, 64, 111, 127, 1, -28, -96, 51, -85, -36, 4, -128, 0, -56, 1, -61, -128, 35, -128, 127, -128, -128, 127, 127, -6, 127, 13, -128, 14, -66, -128, 127, 127, -128, 1, 127, 126, -28, 127, 30, 94, 39, -128, 56, 127, -3, -104, 71, -128, -128, -128, -20, 45, -128, -128, 127, -41, -128, 57, 127, 73, 12, -17, -128, -76, -38, 5, -128, 77, -128, -128, -128, -60, 127, -9, -128, 127, 119, -128, -128, 127, 127, -128, -59, -128, 57, -127, 32, 91, -128, 127, 127, -38, 7, -122, 87, 87, -128, -100, 60, 127, 31, -124, -102, 100, -122, -7, 127, 106, -128, 73, 36, -128, -128, -128, -128, 73, -23, 122, 0, -128, 88, -8, -55, 70, 90, 59, 34, 60, -88, 17, -128, 120, 8, 43, -94, -122, 127, -128, -117, -128, 39, 74, 73, -82, 26, 127, -15, 59, -128, 127, 4, -108, 127, -119, -91, 127, 18, -128, 127, 127, -128, 58, 127, 63, -128, 26, 85, -128, 83, 127, 56, 35, -128, 99, 127, -83, 72, 112, -128, -128, 119, -128, -116, 127, -128, -128, 92, -128, 66, 127, 48, -128, -46, -72, -123, 127, 127, 56, 23, -51, 127, -99, -128, 93, 127, 127, -128, -2, -56, 127, 97, -128, 11, 127, -75, -128, -3, -122, -128, 78, 127, 30, 127, 127, -128, 12, 127, -99, -128, -32, -59, 127, 127, 12, 127, -128, -97, 127, 8, -28, 78, -128, -78, -98, -97, -3, -128, 127, 127, -41, 127, 127, 21, 75, 52, -128, 5, -128, 63, 80, -128, 82, 127, -123, 127, 11, -6, 127, -63, -128, 127, 127, -128, 94, 127, -95, -79, 127, 29, -55, 127, 23, 63, -128, 89, -54, 68, 127, -128, 127, 60, -92, 30, -128, 36, 127, 127, -24, -1, -128, 127, -128, -128, 127, 127, -68, -128, 127, 127, -58, 127, 127, -35, -17, 122, 127, -128, 127, 56, 127, -56, 127, 63, -128, -128, 97, -128, -128, 127, 127, -128, -9, 62, -128, -128, 127, -128, 78, 127, 3, 11, 52, -128, -128, -68, 10, 122, 73, -12, 127, -128, 19, 127, -128, -61, 127, -11, 127, -64, 127, 94, -59, -1, 119, -128, 24, -128, -116, 127, 127, -128, 127, 127, -41, 13, 99, 60, -128, -107, 127, 96, 6, -128, -128, 127, -128, -24, 127, -76, 117, 22, -58, -128, 8, 125, 127, -128, 45, 127, 127, -128, -72, -6, -128, 87, 116, 127, 14, 56, 127, 127, -128, -105, 40, -128, -128, 127, -86, -128, 94, -128, -128, -88, -79, 15, 99, -128, -128, 127, 127, 78, -29, 6, -128, -128, 127, -34, -28, 107, 127, 126, -128, -94, 127, 3, -1, -2, -128, 127, -14, -128, -128, 127, -128, -128, 28, -128, 127, 127, 127, 116, 52, -128, -128, -128, 127, 127, 79, -91, 127, 76, -128, 127, 127, -128, 4, 127, -128, -128, 127, -110, 93, -128, 105, 127, -128, 29, 122, 29, 12, -74, -90, -85, 127, 30, -128, -44, -128, -128, 86, 127, -100, -74, 81, 62, 127, 53, 127, 127, -95, 116, 127, -128, 127, 127, -128, 127, 127, -128, 47, 127, -128, -128, -11, -128, -128, -20, 127, 82, -44, 127, -94, 127, 127, -53, -128, -62, -128, -128, -128, 125, 18, -28, -31, 127, -128, -128, -115, -75, -74, -104, 127, 127, -128, -122, -128, -128, 80, -128, -128, -2, -57, -128, 12, -115, -1, 127, -128, -128, 127, -128, -128, 127, -49, -128, -128, 127, 65, 13, 127, -89, 99, -128, -115, 127, -128, -104, 127, -128, 92, 127, -128, -87, -105, 127, 69, -128, -26, 87, 65, 89, -128, 127, -123, -10, 127, -128, -128, 127, -28, 51, 127, 87, 127, 28, -41, -128, -63, -128, -128, 28, 22, 127, -11, -128, -107, -128, -32, -128, -128, -41, -46, -128, -128, 127, 127, 127, 57, -25, 5, 127, 47, 127, -128, -37, 127, -86, -128, -56, 127, 17, -120, 127, 127, -128, 115, -11, 0, -119, 127, -32, 30, 127, 127, -64, -128, -48, 127, 127, 18, -128, -128, -72, -128, 24, -128, -128, 127, 104, 74, -128, -61, 52, -128, -128, -54, 38, -104, -30, 87, -128, 127, -128, -128, 127, 127, -70, -128, 40, 127, -63, -4, -37, 35, 127, -128, -20, -128, -56, -128, -128, 127, 102, -128, 127, 127, -128, -82, 127, -39, 40, 127, -128, -128, 127, 74, -128, 127, 127, -97, -107, -93, -128, 90, -1, 81, 127, -68, -128, 127, 127, -128, 127, 127, -128, -128, 57, 66, -128, -127, -92, 122, -91, 127, 127, -128, -36, 103, -128, -128, 127, 127, 68, 0, 121, 127, 127, -93, 127, 127, 59, 22, -128, -20, 117, -92, -128, 127, -103, 30, 127, -128, 108, 127, -128, -128, 100, -128, -128, 127, -128, 127, 127, -26, 127, -106, 119, 53, -82, -128, 127, 127, -38, 8, -66, 127, 83, -117, -7, -73, -90, 127, -128, -128, 127, -85, -25, -128, -128, 30, -128, -128, 19, -128, -128, -24, -47, -17, 11, 105, -32, -128, 127, 127, -128, -4, 97, -121, 45, -128, -128, 102, 127, -108, 114, 127, 9, -20, 127, -128, -128, 127, -18, -128, 127, 127, -128, -78, 121, 127, 93, -20, 127, -44, 127, 9, -128, 24, 74, 127, -17, 127, 57, 127, 15, -128, -128, 127, 25, -123, -128, -43, -10, 23, 25, -75, 47, 43, -128, 127, 82, -128, -102, 127, -70, -126, 87, 95, 127, -128, 127, 91, -66, 87, 127, -128, -108, -128, -13, -44, -117, 127, -102, -117, 127, 102, -120, -128, 110, 127, -128, -128, 9, 127, -128, -128, 127, -128, -128, 110, -128, 93, -112, -128, 120, -124, -128, 11, -38, 127, 127, 81, 112, -128, -128, 42, -117, -128, 127, 87, -128, -62, 127, 24, -128, 127, 58, -128, -40, 124, -128, -128, 46, -128, -128, 127, 3, 127, 127, -121, 127, 86, -74, 102, -128, 13, 127, -54, 127, 127, 24, -128, -107, -114, 127, 127, -128, -2, 127, 21, -128, 114, 127, -40, -128, 127, 127, -128, -8, 127, -128, -120, 112, -123, -128, 81, -13, 65, 127, -128, -98, 127, -128, -128, 127, -128, 19, -2, 127, -128, -128, 127, 44, -119, -128, 47, 127, -128, 40, 88, -128, 127, -128, -119, 92, 63, -128, 106, -87, -17, -128, 127, 127, 46, 104, -60, 48, -128, -128, 18, -128, -111, 0, 127, 88, -128, 127, 127, -91, -103, 127, -43, -128, 127, -21, -128, 127, 85, -128, 127, 56, 17, -64, -7, -128, 127, 58, -128, 127, -24, -128, -71, -128, -128, -100, -128, 36, -128, -128, 102, 127, -128, -128, 126, -128, 42, 127, -125, -23, 64, 64, 127, -128, -81, 127, 11, -128, -128, 46, -128, -79, 65, 35, 117, 99, -128, 127, -128, -21, -5, 3, 123, -108, -14, 127, -128, -128, 114, -128, 70, 127, -105, -114, 127, 127, 65, 2, -63, 127, 127, -128, 60, 127, 26, 41, -128, -9, 70, -51, -128, 127, 12, 27, -88, 103, 5, -128, 82, 55, -117, 127, 5, -128, 99, -3, 35, 68, 127, 127, 127, -128, 20, 71, 127, 113, -128, -9, 127, 127, -128, 127, 127, 40, -88, 127, -128, -128, 114, -128, 116, 127, -128, -128, 100, -128, -128, -21, -128, -30, 127, 60, -78, 127, -128, -128, -21, -128, -128, 127, -128, -128, 78, -128, 127, 127, 54, -128, 127, 79, -128, 127, 127, -36, -128, 70, 127, -128, -128, 12, 127, -55, -128, 127, 127, -128, -99, -128, 127, 60, 25, 127, -24, 112, 34, 45, -128, -10, 127, -128, -13, -113, -111, 127, -86, -38, 127, 3, 127, 104, -43, 99, 127, -7, 25, 40, 52, 127, -126, 127, 53, -128, 127, -55, 96, 127, -105, -122, -65, -128, -128, 25, 96, -98, 48, 40, 127, -82, -29, 127, -111, 127, -128, -128, -128, -4, -44, 18, -78, -19, 127, 120, -128, 127, 76, -18, 83, -5, -128, -76, -128, 74, 108, -128, -97, 1, -128, 127, 108, 110, 127, 65, -54, 26, -18, -128, -66, 127, 69, 127, 127, -128, 15, 31, -128, -85, 127, 82, -48, 99, 127, -43, -128, -94, 121, -117, 127, -9, 54, 87, -128, 19, -128, 127, 106, 127, 42, 20, 127, 127, -128, 31, 127, 98, -128, -128, -61, -128, -128, 34, -17, -128, -47, 57, 78, 127, -128, -83, 127, 127, -128, -128, -46, 127, -128, -128, 39, 43, 127, 83, 127, -128, -128, 127, 27, -128, -128, -128, 7, -128, -128, -97, 127, -55, -128, 24, 5, 95, 127, -128, 57, 99, -47, 81, -32, 127, 83, 108, 127, -128, 127, 98, -128, 127, 127, -128, -128, -78, -46, -103, 43, 127, 127, 102, 116, -17, -51, -74, -128, -95, 127, 114, -65, -128, 25, -46, 54, -76, 127, 109, 127, 100, 85, 20, -32, 89, 48, 88, -128, 6, 127, -82, -128, 59, 127, 3, -85, -128, 127, 127, -128, -128, 127, 79, -128, -27, 127, 88, -85, -53, -44, -18, 111, 120, 106, -69, 127, 70, -128, 103, 27, 127, -128, 127, 94, -128, -40, 127, 68, -14, 127, -8, 45, 74, -128, 78, -119, -112, 127, 127, -128, 127, 127, -128, -128, -128, 127, 26, -95, -49, 127, -74, 18, 82, -128, -60, -128, 13, 1, -41, -83, 127, -20, -68, 54, 127, -4, 42, 127, -100, -128, 124, -128, -72, 127, 127, -60, 79, 127, -128, -49, 127, -128, -78, 127, -116, -128, 95, -128, -77, 30, -74, -128, -107, 127, -59, -128, 127, 127, -128, 12, 7, 17, 66, 127, -128, 127, 26, -128, -128, 15, 29, 127, 104, 124, -128, 21, 127, 85, 126, -7, 95, 73, -128, -23, 127, 127, -128, 15, -39, -128, 127, 127, -31, 127, -17, -83, -18, 27, -128, 127, -128, -128, 69, -69, -40, 127, -128, 127, 127, -128, 127, 18, -24, 6, 18, 127, -128, 127, -82, 96, 43, 127, 70, 127, 127, -28, -32, -104, -128, 8, -128, -103, 127, -128, 127, 91, -128, 77, 127, 63, -128, -128, 54, -128, -128, 24, 127, 75, -79, 127, 127, -128, 28, -128, 127, 127, 19, -29, -44, 127, 127, 127, 127, 127, 113, -52, 111, 127, -121, 113, 78, -26, -128, -128, -58, 127, 52, -128, -128, -128, -76, 4, 127, -71, 127, 127, -128, 69, -128, 46, 78, -128, 91, -60, -18, 71, 53, -76, 127, -128, -128, 127, 127, 4, -72, 15, 127, -99, 127, 107, -128, -128, 105, -128, -128, -128, -71, -128, -92, 127, 127, 125, -120, -41, 127, 127, 58, 127, -3, 127, 36, -128, 112, -42, -21, -82, -108, -106, 127, -128, 127, 127, -128, -44, -17, -91, -12, 59, -128, 127, -128, 127, 25, -128, -128, -76, -128, 81, -81, -128, -34, 127, -24, 30, 127, -57, -128, -128, 127, -128, -128, -15, 100, 127, 22, 66, -104, -72, -83, -31, -22, 27, 3, 127, 127, -128, -3, 6, 126, -128, -128, -5, -128, 127, 127, -128, -73, -1, -128, -128, 127, 127, -58, 127, 127, -128, -99, 94, -128, -128, 64, -126, 127, -92, -49, -17, 34, 127, -128, -128, -45, -128, 79, -128, 59, 127, -128, -73, 86, -128, -41, -43, -55, 127, -128, -35, -77, 127, -59, -128, 127, 127, -100, -66, 127, 94, 127, -128, 127, 27, -128, -123, 127, -128, -94, 127, 127, -51, 127, 127, -128, 127, 105, -128, 12, 99, -128, 115, -35, -128, -25, -128, -128, 52, 127, 127, 41, 92, -128, 127, -53, -128, 127, 29, -128, -72, 37, 127, 127, -128, 127, 125, -128, -128, -66, 127, 83, -128, -95, 127, -128, -128, 46, 127, 79, 55, -68, 127, 127, -128, 127, -128, -128, 127, 28, -128, 127, 127, -128, -79, 127, -128, -128, 34, 52, 74, -65, 44, 127, -128, -128, 83, -42, -104, 41, -7, 127, -128, -128, 127, -7, -5, 127, -128, -128, 127, -93, -128, 127, -31, -68, 127, 127, -58, -128, -40, 127, -128, -128, 57, 37, -128, 127, 127, -128, -32, 127, -46, -128, -2, 17, -128, -128, 127, 0, 64, -128, -128, 75, -128, 127, 110, -128, 47, 13, 64, -110, 44, -83, -128, 127, 54, 85, -128, 127, 127, 82, -92, -121, 25, 113, -119, 127, -23, -41, -128, 127, 105, 127, -122, 127, 34, -128, 66, 41, -96, -94, 98, -128, 59, -128, 74, -128, -128, -128, 69, -39, -128, -88, 100, -85, 124, 127, -61, 127, -116, 127, -87, -61, 59, -128, 127, -114, 18, 127, 9, 127, -2, -128, -128, -125, 87, -128, -128, 127, -1, -25, 94, -128, 110, -128, 127, 75, -111, 127, 127, -128, 11, -126, -128, 127, 127, 96, -107, -25, 26, -12, -27, 127, -88, 36, 75, 127, -128, 127, -15, -119, 127, -128, -51, 127, -24, -128, 127, 43, -128, 32, 77, 125, 127, -128, -85, -2, -95, -104, -62, 127, 108, -57, -128, 127, -90, -121, -128, 78, -105, -128, -128, 127, -2, -96, 127, 42, 127, 127, 36, 82, -128, -128, -75, -30, -106, -128, -7, -13, -6, 127, 3, 127, 127, -39, 127, -128, -128, -117, -75, 97, -23, -107, -128, -17, 127, -128, -128, 127, -128, -128, 127, -13, 24, 127, 127, 86, -109, -128, 75, 61, -128, 127, 49, -128, -128, -128, 127, 127, -91, -49, 59, 127, -128, -128, 127, 127, 127, 45, 127, 98, 19, 127, -127, -71, -128, 104, 127, -128, 15, 127, -104, -128, -104, 127, -57, -86, 127, 127, -48, -52, -123, -115, -128, -114, -56, -72, 5, 63, -43, 49, 127, -128, -47, 98, -128, 125, 65, -128, -128, 83, -128, -59, 127, 127, 29, 95, -128, -128, 49, -112, 127, -128, -128, 127, -128, -128, 71, -128, -106, -112, 127, 91, -2, -22, 127, -85, -128, 127, 127, -128, -29, 55, -32, 127, -15, -45, 112, 127, -128, 35, 100, -106, -60, -38, -128, 127, 127, -128, 24, 127, -82, 127, -128, -1, -2, -128, -128, 127, 127, -128, 34, -128, -128, -114, 120, 127, -104, -128, 6, 127, -116, -128, 127, -42, -128, -27, 12, -114, -128, -128, -128, 12, 127, 10, -66, 9, -128, 9, -128, -128, 93, 36, 127, 127, -128, -95, 127, 20, -128, -24, 73, -128, 87, 87, -37, 127, -128, -90, 127, 127, 24, 82, 51, 127, -72, -128, 127, 127, -128, -128, 22, 127, 10, -128, 127, 127, -128, -128, -6, -128, 75, 127, 96, -117, -61, 11, -11, 9, -128, 127, 41, -104, -128, 127, -2, -66, -71, -61, 127, 36, -128, 127, 127, -70, 124, 85, -59, -35, 127, -128, 127, 56, -93, 127, -37, -128, -49, 127, -31, 22, -128, 24, 127, -121, -128, -128, 127, -128, 87, 127, -128, -23, 46, -45, -128, -69, 127, -26, -128, 13, 127, -60, 127, -128, 82, 122, 90, 56, 127, 127, -128, -128, 102, 127, -128, 127, 127, -128, -13, 127, -40, -128, -9, 127, -128, 125, 127, -40, -128, -128, 127, 127, 1, -128, -128, 27, -128, 127, 127, 19, 127, 127, -128, -103, 124, -128, -128, 127, -42, -128, 127, 127, -103, 127, -128, -115, 49, -128, 127, 127, 70, -128, -37, 127, -128, -76, 74, 106, -128, -65, -122, -128, 69, 49, -27, -27, -128, 102, 127, -128, -128, 127, -128, 127, 120, -94, 127, -73, 127, -128, -128, 127, 62, -90, 56, -128, 22, 127, -122, -128, 127, 36, -128, 14, 127, -128, -128, 37, -24, 127, -68, -128, 11, 127, 55, 36, 93, -56, 44, -47, 122, -128, 37, -128, -36, -26, 127, -57, -128, 90, 127, -126, -128, 82, 127, 92, 29, 9, 14, 71, -121, -128, 91, 91, 123, -128, -48, 127, 51, -87, -109, 104, 26, -128, -128, 127, -2, -128, -14, 127, -105, -128, -85, -78, 96, -128, -115, -8, -128, 75, 127, 127, -64, 127, 127, -128, -128, 68, 47, -128, -74, 127, 74, -121, -120, -112, 127, -109, -37, 9, 15, -100, -22, 54, -128, -44, -55, 127, 10, -14, 94, -128, 127, -90, -126, 1, 21, 127, -24, -128, 127, 127, -128, 75, -63, -128, 127, -64, -128, 114, 127, -128, -112, 127, -128, -91, -34, -128, 127, -128, -36, 24, -128, 127, -47, -95, -58, -58, -2, -58, -20, 127, -128, -128, 87, -128, -128, 127, 28, -125, 127, 127, -103, 78, 127, 66, -128, -128, 112, -128, -76, 127, -125, 11, 127, -70, -128, -128, 127, -23, 74, 127, -96, 127, -76, -128, -108, -128, 55, -128, -128, 127, -128, 10, 127, -58, 127, 127, -15, 14, -128, -128, -35, -128, -87, -128, 127, 127, -68, -111, 27, 55, -128, 58, -61, 127, -128, -90, 127, -59, -128, -18, -31, -128, -128, 127, 46, -128, 92, 127, -34, 127, 89, 41, 97, 7, -22, 64, -128, -128, 127, 38, 68, 59, 127, -6, -128, -114, 29, -128, 127, 106, -128, 86, 127, 127, 79, -128, 23, -128, -128, 127, -97, -128, 127, -128, -128, -19, 20, -42, -128, 112, -128, -76, 127, 81, -128, -7, -81, -66, -128, -21, 127, -128, -128, 122, -128, -128, -128, 59, 127, 56, -128, 127, 127, -128, 62, -43, -128, 127, -109, 39, -128, -87, 127, -128, 127, 127, -128, 127, 127, -58, 127, -128, 127, 127, -128, -45, 127, -32, -63, 1, -128, 75, -4, -128, -51, -128, 73, -69, -128, 127, 82, -128, 127, -82, -77, 46, -128, 127, -128, -128, -72, 127, 5, 127, 127, 106, 60, -70, -25, 127, 127, 127, -30, -128, 4, 127, -128, -128, 127, 83, 44, 127, 127, 82, -128, 100, 127, -128, -128, 93, -128, -128, 78, 127, -128, -128, 127, -77, 127, 127, -35, 127, 127, 127, -49, -128, -128, -51, -85, -128, 127, 127, -128, 64, -128, -128, 127, 115, -29, -45, 105, 20, -11, -128, 127, -82, -37, 127, -128, -128, 127, 127, -61, 108, -46, 47, 127, -128, -116, -14, -128, -96, 127, 127, -99, -97, -128, 89, -38, 95, -128, -128, 127, -128, -128, 47, 127, -128, -72, 23, -105, 43, 127, -128, -112, 127, -128, -42, -5, -128, -61, -26, -128, 90, -128, -102, 127, -21, 58, 127, -86, 127, 127, 4, -42, 127, 127, -128, 122, -128, -128, 127, 127, -6, -41, 13, 127, -113, -128, 8, 53, -85, 107, 127, -128, 127, 127, 7, -128, -21, 27, -128, -128, 127, 78, 79, 77, 122, -55, -128, -68, 127, 77, 102, -73, -128, 104, 127, -94, -53, 127, -81, -128, 127, 127, -128, -12, 127, -128, -51, 86, 127, -128, -128, 77, -128, -128, -79, 119, 43, 127, -99, -128, 123, 111, 18, 98, 127, -125, 40, 127, -128, -128, 127, 127, 59, -128, -21, 49, -6, -87, -30, -128, 127, 58, 94, 127, 7, 59, 3, -128, -128, 38, -128, -128, 29, 127, 127, 120, 10, 37, -41, -128, 48, -12, -128, 96, -90, 127, 65, 75, -128, 127, 127, -128, 127, 127, -128, -128, -110, -128, -52, 26, -128, -65, 127, 127, -81, 63, 27, 127, -128, -97, -73, -77, -103, -100, 127, -123, 5, -52, -128, 47, -29, -128, -22, 127, 92, 104, 127, 38, 70, -30, -128, -128, -128, 36, 127, -12, -2, 127, 37, -23, 0, 127, -128, 86, 127, -121, -21, 127, -108, -89, -128, 127, 106, -128, 19, 127, -49, 127, -128, 127, 110, -40, -128, 127, 102, -128, -9, 127, 0, -128, -52, 127, 58, -128, -113, -11, 127, 127, -110, 127, 127, -128, -128, -39, -128, -7, 127, -91, -123, 25, -57, 127, -128, -49, 32, -128, 59, -128, -128, 3, -128, 90, -49, -113, 85, 30, -60, -44, -128, 36, -44, 127, 127, -35, 44, -5, -127, -128, 125, -10, 127, -128, -40, 23, 127, 2, -89, -128, -120, -128, -10, 93, -31, 91, 127, -128, 127, -65, -128, 113, 69, -128, 26, 0, -128, -77, 127, -116, -40, 24, -11, -41, 119, -128, -94, 115, -128, -14, 127, -116, 9, 127, -128, 97, 4, -128, 41, -128, 127, -71, -128, 94, 126, -128, 53, 93, -128, -128, 127, 90, -128, 108, 127, 6, 39, 36, -128, 91, 127, 76, -93, 127, 127, -128, -128, 69, -29, -128, -128, 126, -128, -15, -66, -128, -128, 61, -88, -102, 127, 127, -66, -83, -128, 94, 127, 127, -124, -3, 127, 127, -128, -128, 68, 127, -26, -19, 127, 113, -128, -128, 127, -128, -128, -87, 94, 55, -128, -128, 127, -128, 19, 97, -106, 127, -52, -128, 52, 96, 127, 127, -128, 83, 127, -128, 39, 86, 72, 65, -128, -7, 127, -10, 75, 97, 24, -49, -128, 127, 127, -21, 36, 127, 127, 37, 77, -28, -18, -123, -128, 127, -128, -128, 127, 127, -58, -128, -35, 127, -128, -128, 3, -128, -91, 66, 127, -32, -128, 127, -31, -128, 27, 127, -125, 14, 127, 75, 26, -13, 127, -128, -128, -128, -1, -76, -88, -81, 87, 83, 8, -127, -128, 127, -3, 98, -57, 55, -45, -80, -128, -128, 45, 49, -53, -128, -7, -128, 127, 110, -117, 2, -128, 91, 127, -128, -15, 127, -128, -128, 61, 125, 57, -128, 127, 127, -128, -116, 127, 90, -128, -74, 109, 75, -47, -11, -105, 35, -128, 127, -128, -68, 127, -104, -23, 114, -122, -120, 127, -99, -128, -103, -113, -128, -128, -3, 113, 127, -128, -1, 122, -125, 127, -128, -24, 127, 49, 77, -25, 59, 127, -51, -128, -42, 127, -128, -24, 127, -128, 29, -107, 127, -116, -128, 23, -65, -41, -72, -128, -56, -128, -39, 39, -128, 127, 127, -128, 127, 127, -54, 1, 125, 127, -85, 71, -128, -128, 127, 45, 30, 45, 127, -8, 117, 127, -64, 127, -128, -112, -109, -128, 127, 76, -61, 62, 127, -128, -128, 127, -29, -102, -3, -97, 127, 127, 106, -128, 78, 127, -128, -128, 127, 103, -128, -128, 88, -41, 88, -128, 41, 95, -128, -128, 127, -128, 88, 97, -128, 127, -128, 91, 127, -128, -27, -128, 77, -21, 17, 127, -128, 49, 127, -128, -128, 81, 71, -71, -128, 32, 89, -75, -114, 127, -128, 15, -128, -128, 0, -128, 47, 60, -82, -128, 127, -128, -4, -58, -128, 127, -35, 72, 127, 110, 127, 34, -128, -46, -92, -106, 127, 72, -46, 64, 127, -41, -128, 30, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 21 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
