-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
            -13, -13, -3, -2, 2, -3, -9, 17, -1, 14, 2, -20, -20, 14     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( 41, 36, 66, -33, 119, -21, -55, -6, 75, 76, 14, 84, -90, 54, 17, -24, 105, -34, -79, 42, -90, -19, -32, 101, 9, 81, -20, 51, -124, 84, 18, -52, 98, 28, 57, 110, -19, -99, -84, -119, 33, 5, 119, 17, -44, -3, -16, -119, -61, -56, 124, 19, 71, -52, 110, 26, 105, 67, 124, -18, 42, 22, 51, -99, 79, 114, -62, -56, 25, -80, -88, 75, 68, -36, 49, 31, 60, 67, -12, 118, 9, 75, 111, 65, 15, -2, 37, -27, 15, 36, -99, 77, -88, 91, 13, -32, 2, 56, -45, 44, -100, -52, -109, 38, -114, 6, 0, -127, -117, -99, -26, 88, 110, -83, -110, 104, 70, 15, 114, 80, -6, -123, -87, -49, -77, 16, -74, 19, 95, 59, -74, 78, -61, 100, -117, -110, -115, -16, -90, -106, 80, -43, -36, 35, -81, -51, 31, 52, -18, 17, 111, 121, 107, 62, -123, -100, 111, 92, 45, 56, 105, 84, -52, -26, -74, 68, -69, 31, 60, -4, 55, 49, 107, 85, -51, 16, 54, 99, 92, 99, -40, 124, 19, -14, 19, -25, -101, 107, -4, 41, 88, -109, 7, 112, -13, -40, 103, -37, 127, -119, -76, -56, -75, -77, -127, 57, -36, -20, -23, 95, 91, 90, 47, -107, -117, -101, -52, -2, -77, 85, 7, -113, 43, 31, -82, 119, 105, 35, -104, -119, -19, 86, 55, -57, 76, 57, 33, 70, -22, 48, -29, -126, 91, 76, 29, -61, 14, 27, -25, 29, 119, 60, 112, 79, 80, -94, 90, -92, 48, -113, -88, 117, -21, -41, 74, -18, 101, 1, -79, 9, -36, 6, -73, 38, -113, 8, 37, -121, -24, 28, -39, 29, 64, -44, -65, -17, 72, 36, -55, -25, -95, 115, -54, 108, 21, 43, -87, -74, 10, -58, -62, 95, 28, 65, -116, 59, 53, 6, 47, -17, 48, -2, 3, -50, 9, 15, 74, 122, 107, -74, -85, -60, 103, 121, -61, 105, -42, -49, -115, -38, 109, -88, 28, -53, -116, -103, 81, 49, 98, 120, 71, 46, 88, -92, 28, -92, -83, 62, 108, 42, 99, -85, -92, 6, 80, -13, -12, -76, -14, 54, 103, -87, -72, 124, 61, -62, 33, 22, 67, 27, -36, 59, -10, -38, -21, 6, 89, 1, 40, 71, 79, -68, 1, -72, 9, -100, 89, -128, 9, 113, 20, 95, -4, -1, -61, -61, 35, 44, 95, 0, 51, -1, -23, 65, 67, -25, 2, -90, -6, 53, -61, 66, 81, -121, 3, 43, -94, 69, -95, 29, -109, 123, -4, 106, 44, 2, -76, 56, 97, -3, -5, -52, 110, 103, -121, -91, -59, 91, 9, 120, -69, -97, -42, -108, -69, -33, -87, 53, -3, -112, 87, -101, -50, -22, -95, 73, 97, 35, 74, 124, -39, 88, -16, -96, -125, -81, 49, 88, -56, 111, 59, 10, 64, -70, 46, -39, 60, 104, -24, -125, 70, -28, -122, 66, 125, -109, 104, 104, 62, 61, -125, 18, -121, 78, -77, -124, 114, -72, -69, -96, -110, -23, 2, 11, 75, -50, -63, 103, 111, 93, 45, 26, 45, 118, -4, -1, -115, 45, 112, 66, -90, -18, -86, -2, 26, 7, -43, 25, 63, 67, -122, 13, 113, 95, 126, -9, 85, -108, -52, -59, 59, 91, 127, 28, 40, -48, -99, 63, 46, -122, 10, 113, 61, 57, -109, -92, 13, 103, 76, -52, -35, -67, 93, -14, 2, -22, -43, 8, 4, 37, 37, -88, 94, 70, -77, -87, 127, 39, -45, 115, -78, 110, -105, -46, 51, 2, -29, -63, -122, 22, 40, 84, 127, -16, 9, 49, 25, -96, -89, -50, 29, -106, -8, 126, -13, 125, 88, 48, 56, -30, 104, -13, 118, -95, 125, -81, 69, -128, -100, -48, 85, -21, 75, -60, 63, 112, 79, 37, 105, 105, -79, 75, -128, 102, -35, -98, 19, -97, -121, 72, -32, 77, 95, -74, -26, 77, -83, 111, 36, 5, -75, 110, 118, 51, -44, -86, -122, 39, 88, 78, 55, 102, 32, -64, -97, 120, -89, -16, 58, -15, -22, -81, -10, 85, 121, 70, -14, 57, 21, -112, -43, 101, 58, -86, 88, -121, 55, -9, 12, 68, 25, 116, 55, -104, 121, 70, 19, 43, -103, 60, 95, -111, 93, 111, 32, 127, 8, -14, 16, 83, -48, -125, 111, 105, 95, -107, 48, 57, 17, 100, 32, 5, -119, -65, -98, -75, 56, -106, -43, 68, -93, 5, 88, -62, 22, -48, -96, 106, -14, -67, 126, 52, -103, -3, -61, 87, -70, 89, 102, 67, 127, -15, -36, 37, -106, 76, -6, -30, 68, -113, -60, -58, -79, -2, -6, 38, -64, -77, 98, 103, -108, -56, 53, -78, 58, 107, 79, -53, -30, -90, -20, 56, 79, -77, -75, -17, 5, 116, -12, 92, 63, -12, -17, 8, -109, -40, 56, -32, -31, 33, -86, 67, 57, -50, 60, 41, 75, 93, 61, 117, 38, 104, 36, 44, 11, 19, -21, -123, 17, 3, 12, 4, -61, -62, 65, -8, 37, 36, -20, -12, -80, 115, 103, -111, 103, 43, 123, -65, -95, -31, -63, 11, 7, 125, 62, 110, 101, 74, 109, 120, 94, -117, 26, 12, 40, 70, -1, -89, -27, -112, -82, 110, -101, -27, -126, -35, 67, 69, 32, -22, 70, -114, -107, 56, 19, 12, -57, -28, -48, 99, -48, 65, -77, 5, 102, 50, -116, 77, -4, 107, -87, 62, -87, 83, -66, -67, 118, -14, -40, 78, 94, 33, -7, 8, -127, 102, 30, 113, 17, 29, -21, -120, 43, -114, -36, -99, -83, 59, 94, -95, -122, 46, -82, 50, -61, 58, -54, -111, -49, -117, -4, -56, -30, 71, 113, 93, -20, 112, -51, 57, 26, 121, -113, 122, 91, 36, 65, -27, -46, 28, -60, 31, -105, 23, 19, -12, -1, 52, 37, -69, 11, -106, -81, -93, 19, -85, 6, 11, 55, -20, -68, 6, 53, 119, -106, -116, -13, 37, 44, -106, -36, 41, 113, 126, -73, 22, -86, 23, 46, -108, 27, -8, 54, -48, 82, -22, 15, 85, -3, -99, 77, -103, 51, -46, -85, 66, -11, 107, -116, 13, 57, -53, -93, 121, -128, -19, -20, 68, -88, -35, -87, 104, 19, 5, -94, 52, 4, 68, 81, 10, -24, 112, -45, 35, 76, 9, -90, 18, -34, -58, 85, -43, 81, -33, -120, -112, 49, -6, 81, -64, -81, 96, -37, 97, 41, 96, -22, 40, -85, 0, 20, -60, 101, -49, -99, 33, -68, -10, 33, -59, -112, 86, 86, -17, -4, 116, 83, 10, 111, 96, 77, -54, -67, -19, 83, 44, -53, -128, 39, -17, 64, -58, -63, 127, 101, -29, -64, -98, -33, -57, -127, 122, -8, -113, 112, -41, 48, -76, -85, 4, 58, -20, 26, -12, -120, 60, 115, 87, -24, 125, 108, -118, 9, -6, -103, 85, -111, 117, 10, 90, 31, -69, -66, 80, 117, 112, 57, 103, -57, -67, -126, -60, -17, 111, 40, -101, 90, 99, -12, -112, -34, -87, -48, -67, -127, 25, -121, 67, 23, 114, 62, 113, 104, 102, 126, -101, -106, 60, -108, 54, -116, 114, 93, -50, -110, 20, -105, -45, -84, 60, -57, 41, 126, 110, -110, -5, 72, -42, -8, -126, -50, 110, 106, 64, 44, -53, -16, 106, -15, -111, 64, 94, -25, 32, -104, -63, 20, 65, -23, -69, -117, 101, -20, -70, -17, 97, 43, -84, 101, 10, -2, 56, 61, 126, -25, -72, -77, -55, 102, -66, 15, -106, 123, 107, 34, -47, 15, 17, 84, -116, 48, -48, 94, 20, 69, -51, -125, -51, -120, -95, -4, -115, -46, -115, 64, 30, -105, -79, -9, -93, 45, 95, -106, -54, -5, -96, 41, 44, -88, 84, -100, -83, 123, 28, -105, 4, -111, -123, 42, -15, 28, 22, -91, -38, -74, 35, 2, 1, -109, 41, 12, -79, -105, 57, 74, -122, 8, -118, -90, 104, 57, -48, 51, 52, -68, 10, 122, -70, 79, -24, 113, 55, 120, -109, -70, 81, 80, 12, -4, 76, -99, -106, -82, 68, -105, -3, 5, 4, 121, 52, -30, -88, -118, -121, -88, -20, 1, -59, -103, 108, 42, 111, -23, -118, -15, -65, -18, 75, -63, -63, -64, -117, 47, 31, -111, -85, -117, 99, 47, 37, -37, -6, 102, -98, 127, 67, -105, -90, -95, -40, -64, 101, 39, 127, 124, -26, 41, 36, -75, -9, 99, -54, 2, -115, 45, 15, -60, -70, -39, -32, 121, -40, 79, 105, -39, 26, 106, -121, -56, -82, 92, 48, 17, -105, 12, -83, -73, 85, -8, -74, 34, -43, -13, -86, 16, -17, -96, 49, -110, 78, -57, -89, -28, 57, 19, -115, 72, 74, 111, 84, -51, -37, -83, 101, -77, 45, -42, 61, -56, -86, -65, 80, 107, -41, 16, -105, -103, 16, -77, -75, 43, 118, -85, -71, -28, 36, -52, -76, 116, 81, -102, -105, 96, -126, -126, 94, -101, 38, -1, -12, 66, -107, -117, -87, -101, 10, -122, 57, -52, -25, -70, 70, 26, -72, 59, 32, 56, 114, -58, 101, 63, -116, -92, -95, -66, -69, 99, 27, 80, 73, 84, 76, -85, -39, 40, 51, -98, 17, 111, -78, -38, -23, 61, -102, 28, -101, -69, -40, -14, -103, -98, -12, -112, 55, 103, 50, 44, 24, 4, -25, -28, 26, -104, 109, -6, -50, -62, -72, -37, 69, -3, -84, 32, -88, -29, -40, -105, -15, 115, 52, 5, 34, -41, 122, 61, 60, -29, -114, -89, -85, -17, 59, 74, -67, -29, 40, 19, -44, 62, -72, 63, 3, -44, -117, -73, -58, 64, 24, -56, -10, 115, -105, 91, 42, 5, -121, -84, -64, 6, 49, 20, 65, 69, -11, -57, 115, 91, -93, 91, 89, 116, 64, -62, -2, -89, -100, -118, -92, 79, -81, -34, 91, -77, 106, -61, -60, -110, -45, 75, -23, 52, 11, 105, 104, -75, -27, -18, 110, -1, 87, 76, -39, 70, 119, 70, 32, -66, -64, 103, -12, 40, 81, -22, 46, 76, 80, -59, 47, -36, -98, -100, 28, 104, -32, 98, 110, 123, -100, 37, 41, -50, 92, 22, -20, 65, -99, 94, 49, 72, 0, 54, -42, -74, -32, -39, 125, 66, 112, -44, 118, -112, 61, -60, 68, 73, 112, -99, -99, 89, -38, -17, 108, 10, 26, -76, -75, 78, -10, 64, 91, -1, 39, -24, 53, -124, 45, 113, 13, 77, 46, 60, -19, 72, 78, 25, 40, 0, 45, -119, 16, 16, -128, 75, -115, 11, -15, -45, -81, -122, 61, 18, 100, 47, 95, -1, -100, 78, 20, -101, -50, 86, 63, -122, 103, 35, 70, -11, 101, -41, -67, 62, 36, 32, 122, -35, 55, 78, 59, -48, 118, -103, -66, -112, -13, -47, -12, 108, -76, 57, -42, 125, -37, 36, 60, -112, -115, -41, 125, -109, -65, 96, -85, -29, 43, -87, 32, 35, 76, -102, 46, 124, 26, 111, 70, 47, -51, -91, 20, -65, 99, -23, 76, -123, 43, 77, -63, -40, -56, 87, 43, -81, -126, -124, 104, -127, 124, -104, 94, 48, -20, -32, -1, 8, 73, 114, 22, 88, -78, -85, 71, 85, 71, 75, -73, -107, -21, 124, -13, 24, -31, 98, 8, -50, -27, -102, 123, 117, 87, 80, 64, 74, 59, -73, -1, -69, 34, 23, -112, -81, -109, 95, -33, -50, -109, 22, 120, 19, 47, -123, -108, -63, 32, 10, 12, -26, 74, -99, -23, -11, 118, -66, -34, -46, -68, 119, -46, -3, 118, 90, 95, -61, -2, -63, 121, -10, 55, -27, -113, 87, 71, 16, 44, 82, 99, -64, -22, 117, -5, -39, -114, 7, 79, -122, -122, 104, -74, -15, 9, -113, 53, 30, 61, 114, 59, -23, -7, -10, -97, -97, -55, 118, -7, 3, 85, -87, 92, 127, 110, -14, -37, 83, -45, 16, -29, 34, -81, -64, -89, 44, -70, -54, 29, 12, -89, 98, -27, 15, -31, -25, -16, -101, -52, -90, -71, -47, 18, -62, 47, -18, -13, -102, 54, -65, 62, 32, -62, -41, 50, -77, -81, -32, -54, 38, -59, -91, 113, 87, -12, -72, -14, -47, -128, 63, 50, 99, 14, 40, -68, -103, 91, -19, 81, 88, 115, 28, -71, -21, 32, -52, 116, 11, 40, -115, -24, -127, 86, -60, 120, -82, 127, 35, -31, -110, 29, 124, -66, 28, 118, 17, -3, -12, -47, -36, -102, -31, 68, 27, -111, 48, -93, 29, -76, -15, -40, 111, -82, -119, 97, 61, 51, -47, -51, 106, -40, -76, 87, 112, -62, 32, -46, -16, -109, -119, 31, -103, 25, -19, -126, -68, -58, -88, -75, 28, 106, -108, -107, 71, 5, 58, 36, 16, 35, -70, 24, 66, -60, -26, 78, 41, 36, -87, 124, 31, 68, -9, -125, 42, 62, -95, -57, -96, 13, 114, -46, -22, -111, -50, -115, -51, -55, 110, 78, -122, -97, -6, 46, -21, -80, 89, 53, 35, -82, 126, -113, -109, -33, 91, 64, 38, -18, 98, -92, -69, -78, 17, 124, -30, 120, -61, -91, -89, -63, 43, -103, 3, 36, 49, -32, 96, 121, 44, 27, -7, -10, -47, -22, -123, -67, -65, -58, -121, -118, 42, 94, 32, 122, 111, -107, -41, 121, 1, 46, 126, 45, -77, -94, -17, 87, 53, 61, 8, -50, -82, -26, 121, 19, 9, -54, -51, -96, -70, -41, 44, 88, 70, -20, -1, -120, 3, -88, 19, 17, -100, -54, -60, -119, -17, -5, 76, -79, -28, -53, 48, 85, -93, 10, -115, -64, -125, -120, 110, 57, 21, -83, -51, 91, -3, 14, 26, -66, -12, -29, 121, -9, 115, 7, -65, 35, 117, -57, 91, -36, 40, -117, 49, -65, 120, 20, -39, -15, 83, -68, 7, -46, 111, 115, -95, 112, -67, 127, -58, -92, 32, 101, 16, -115, -125, 28, -110, 96, 99, -47, -36, 61, 60, 31, 90, -83, -113, 2, 46, 6, 83, 17, -58, 99, 82, 93, 36, -78, 108, 58, 110, -60, 79, 5, 59, 92, 41, 83, 103, -95, 41, -21, -47, 31, -67, -126, 40, 54, -17, 50, 39, 8, 106, -56, -13, -41, 77, -78, 124, 97, -113, 47, 101, 71, -9, -42, 29, -76, 103, 95, -91, -75, 102, -128, 62, 30, -80, 72, 6, 104, 113, 23, 47, 55, 122, -18, -84, 62, 21, -31, 116, -54, -111, 36, 20, 4, -69, 120, 118, -88, -41, 29, 59, 53, 89, -67, 3, -9, -29, 24, -31, -111, -88, 18, -100, 33, -60, -32, -117, 98, -42, 123, -73, 112, -87, -93, 72, -83, 109, -87, -40, -27, 21, 34, -110, 23, 87, 62, 88, -68, -36, 26, 82, -2, 102, 25, 41, -11, 7, -112, -53, 34, -17, -66, -47, 4, 18, -53, 122, -87, 19, -118, 73, 108, 3, 55, -96, -112, 56, -66, -30, 102, 112, 62, 35, 80, -56, -27, 109, 52, -111, -13, 36, -117, 50, -122, 76, -114, 21, -49, 5, 79, -113, -91, -30, -72, -56, -117, -87, -116, -108, -26, 22, -48, 1, 43, 58, 92, 31, -124, 57, -67, 102, -29, -28, 30, 17, 96, -53, -87, -1, 98, -80, -5, -109, 30, 122, 127, 124, -33, -38, -91, 13, 101, 56, -111, -75, 85, -117, -58, -100, 20, -56, -21, 90, 99, 118, -60, 72, -91, -86, -48, -123, 55, 111, -26, -45, 29, 17, 45, -12, -44, -6, -63, 94, -51, 94, 27, -109, -79, -81, 44, 6, 49, 125, -112, 4, -31, -37, 9, -35, -47, 101, -90, 105, -117, -127, -13, 116, 90, -25, 38, 73, -22, 54, 51, 37, -26, 108, 17, -119, -97, 87, 124, 5, -94, 8, 41, -109, -105, 126, 100, -76, 17, -27, 33, -7, -7, 46, -87, -57, -92, 14, 63, 109, -8, 64, -106, 115, -86, -82, -43, -91, 85, -117, -13, 77, 0, 10, 86, -37, -1, -107, -26, -27, 10, -27, 11, -38, -95, 44, -48, 52, -123, 9, 106, 73, 9, 78, 100, 51, 78, -58, 65, -21, -31, -99, -123, -46, 66, -122, -19, -117, -11, -7, 126, -33, -111, 44, 127, 42, -94, -59, -95, -105, -9, -114, 121, -3, 3, -56, 125, -120, 48, -74, -45, 36, -40, 38, 27, 0, -51, -38, 69, 78, -14, -88, 83, 97, -42, 65, -42, 106, 108, -126, -64, 49, -119, -49, 50, 93, 38, 66, -120, 84, 101, -101, -58, 0, 27, 98, -72, 55, 91, 108, 110, -119, -124, 76, -29, -112, -91, -120, -36, -124, -128, 93, 19, -89, -27, -33, 126, 85, 46, 54, 105, 73, -104, 122, -107, 71, -22, -27, -84, 39, -52, -84, -49, -27, 105, -87, 67, 114, -124, 47, 33, -14, -12, 126, -107, -121, 126, 71, -76, -80, 2, -96, -41, -63, 37, -117, 30, 18, 10, 60, -116, -72, 46, -42, 24, -92, 28, 4, 81, 70, 21, 69, -16, -71, -53, 111, 27, -31, -92, 35, 62, 95, -112, -106, 57, 8, -125, 21, 113, -128, -1, 53, 77, -1, -5, 103, 24, -63, 38, -52, -54, -118, 12, -111, 79, -24, -80, -6, 63, 6, -82, -70, 91, -67, -79, 39, 88, -49, -10, -71, -23, -47, -67, 22, 11, 21, 73, -112, -73, -50, -94, 93, -96, 97, -85, -25, -57, -128, 97, 104, -122, -74, 84, 118, -77, 39, 42, 95, 118, -5, 59, 126, 49, -107, 70, 22, 102, 17, -74, -7, 78, -87, 105, -32, -74, 103, -11, 95, -112, -46, -51, -2, 83, 65, -86, 48, -45, -36, 3, -87, 101, -64, -72, 76, 53, 39, 69, -7, -112, -60, 80, 78, 8, 60, -89, 2, 57, -84, 127, 107, -101, -70, -124, 114, -55, 118, -16, -29, 101, -16, 26, -12, -96, -89, 61, -75, -18, -23, -5, 100, -31, 119, 15, -99, 104, 59, -29, 5, 59, 4, -81, 89, 83, 39, -28, -98, 32, 25, 71, -52, 27, 40, 54, 49, 10, -97, -92, -103, 73, -118, -101, -100, 36, 5, -101, -24, -30, 61, 32, -87, -38, -95, 11, -69, -114, 21, 16, 56, -87, -107, -29, -17, 46, 118, 88, 19, 69, 92, 75, -107, 108, -12, -123, -89, -94, -16, 72, 111, -53, -77, -116, -48, 70, 5, 96, -17, -120, 20, -26, 91, 70, -39, 4, -121, 22, -82, -88, -102, -67, 118, -70, 98, -28, -37, -113, 16, 58, -119, -92, 121, -44, 57, 85, 126, 0, -67, 59, -1, 4, -123, 55, 65, 117, 90, -116, 113, 66, -96, -88, -23, -107, 49, -85, 54, -73, -33, -66, -18, -12, 0, 39, 4, 5, 109, 114, 73, -89, 101, 121, -112, -107, -116, 100, -12, 22, -93, -69, 92, 98, 21, 48, -4, 19, 110, 65, 73, 58, -86, -19, 66, 102, 99, 119, 76, -102, 65, 79, -116, -7, -120, -4, 111, 104, -73, 76, -110, 10, 93, 0, -106, 8, -61, -122, -51, 35, 12, 69, 102, -34, 46, -126, -92, -115, 89, -37, 20, -112, -57, -113, 57, -68, 34, -73, -124, -89, -32, -81, -30, 28, -91, 23, -119, 6, -73, 103, -70, 67, -115, 89, 53, 45, 33, -117, 30, 63, 14, -41, -114, 80, 47, -86, -49, -89, 41, -95, -71, 101, 110, -42, 119, -107, 118, -110, 107, 19, -25, 52, 88, -112, -47, -42, -94, -125, 110, 75, -79, -112, 25, 106, 20, -111, 35, 41, -101, 83, -115, 20, -126, -71, 42, 8, -5, -128, -92, -6, -104, -82, 45, 122, -12, 25, 82, 74, -10, 6, -60, 21, 105, 31, 115, 111, 57, 99, -1, 66, -16, -119, 19, 65, -78, 46, -79, 108, -77, 26, -83, -16, -25, -6, 33, 67, -115, -34, -118, 13, 21, 20, -47, -72, 123, -70, 32, -78, -22, 8, -29, 39, -1, 20, -2, 7, -67, 25, -69, 126, -5, -87, -75, 56, -87, -106, 31, 95, -117, 41, 110, -90, 81, -70, -56, 73, -119, -79, -126, -45, 111, 45, -79, 37, -59, -88, -80, 85, -112, 26, 79, -106, 71, 82, 115, -76, 104, 99, -41, -10, 56, 114, 33, -19, 70, -25, 47, -57, 109, -21, -32, -122, -61, -90, 56, -25, 12, 127, 75, 113, 17, 31, 26, -9, 107, 95, -16, 125, -16, -29, -10, 32, 7, -57, -36, 1, -44, -57, -82, -58, -96, -56, -73, -116, 98, -127, 122, -104, -12, -80, -112, -5, 51, -98, 80, -63, 107, 51, 67, 36, 89, -16, 23, 101, -79, -30, 56, 49, 38, -115, -121, 121, 85, -91, -86, 123, -96, -43, 53, 101, 46, -35, 85, 101, 7, 121, -12, 49, -66, 75, 5, 57, -124, 98, -86, -87, -47, -75, 93, 7, -18, 34, 60, -79, 78, 24, -66, -58, -54, 51, 21, 115, -54, 38, 113, -53, -107, 45, 22, -96, -128, 123, 45, 48, 45, 109, 92, -89, -74, 89, 91, -112, -96, 4, 105, -94, 126, -109, 82, -119, 36, 124, 126, 115, -16, -60, 1, 52, 83, -96, 61, 7, -106, 94, 91, -77, -75, 110, -51, 16, 38, -14, 55, -72, 75, -41, -16, 58, -37, 80, -61, 41, -42, -114, -116, -2, -32, 108, -99, -58, -12, -53, -44, -70, -45, -34, -111, -104, -47, 29, 15, -81, 44, -13, 118, -58, 78, -47, 77, -100, -18, 14, -83, 81, -52, 83, -91, 86, -19, -27, -64, 18, -12, -112, 93, 92, 110, -24, 93, -93, 5, -83, -75, -116, 105, 111, -120, 114, 44, -77, 91, -22, -98, 112, -73, 84, -39, -2, -10, 29, -53, 30, 10, 103, 20, -70, -89, 84, 58, -84, 17, 25, -12, -120, 106, -67, -125, 58, -25, 6, 36, -116, 80, 24, 22, -56, 48, 102, 50, 51, -23, -126, 75, -94, -88, 118, 36, 23, 69, -125, -121, -1, -99, 11, 59, -79, 96, 85, 105, -61, 110, -82, 6, -17, -77, -87, 10, 116, 7, 123, -70, -70, 55, -9, -81, 15, -23, 80, -19, 38, 6, -93, -79, -104, -82, -80, -74, 65, 108, -53, 82, 48, -78, -57, 17, 103, 77, 62, 99, 125, -4, 108, -14, 101, -78, -70, -110, -103, 89, 86, 108, -125, 98, -76, 110, -121, 108, -87, 36, 38, 0, -41, -126, 80, 85, -83, 29, 113, 118, -99, -114, 75, 41, 96, -59, -35, 7, -109, -121, 21, -55, -104, -58, 3, -116, -44, -78, 117, 77, -23, -22, -33, 0, 55, 124, 118, 93, -64, -41, 64, 53, -58, 40, 25, 51, -14, -12, 31, -121, -109, 17, 89, 73, 23, 9, -57, 66, 28, 116, -80, -101, -24, 87, 1, -109, -51, 19, -30, 75, -56, -89, -67, 14, -84, -53, -115, 12, 91, -112, 107, -14, -3, 112, 50, -51, -74, -119, -124, -95, 26, 38, -116, 65, 32, 6, -70, -128, 89, 94, 55, -84, -82, 23, 113, -25, 74, -86, -76, 45, 66, 88, 71, 78, -104, 33, -124, 22, 119, -89, -43, -4, 98, -6, 121, -122, -40, -25, 85, 99, -128, 34, 114, 88, -77, 105, 85, 36, -10, -72, -102, -10, -48, -57, -46, 125, 98, -59, -1, -86, 78, -19, 73, -4, -34, -26, -16, 124, 38, -4, 98, -102, 72, -52, 53, -88, -110, 4, -64, -9, -109, 62, 101, -75, 12, 13, 18, 112, 59, 80, -12, 124, 91, -46, -9, 51, 99, 108, -69, -20, -36, 121, 52, 21, -83, 12, 42, -77, 108, -22, 120, 59, 16, -13, 39, 91, -120, 85, -41, -78, -87, 2, 119, 77, 22, 103, 71, -51, -24, -86, 31, 63, 38, -98, 51, 1, -37, -7, -1, 105, -45, 51, 120, 87, 30, -23, 98, -48, -113, -124, -28, 92, -69, -107, -71, -88, -52, -32, -65, -78, -32, -127, -11, -103, -101, -11, 10, -15, -70, -9, -28, -87, -10, -90, 51, 5, 104, -101, -50, -42, -52, 110, -117, 60, 31, -112, -14, 102, 86, -18, 90, -97, -7, 61, 125, -54, -72, 35, -67, -103, 111, 35, 64, 21, 7, 6, -66, -29, -79, 18, 9, -3, 119, 99, -124, 83, -46, 15, -21, 55, 53, 31, 111, -87, 81, -53, 99, 115, -62, 115, -104, -72, 16, 79, -85, 83, -26, -11, 125, 51, 25, 126, 107, -90, -101, -65, 86, 121, -105, 94, 93, 125, -125, 104, 80, 91, -73, 73, -51, -25, 78, -77, -83, -33, -68, 2, -107, -97, -19, 84, 63, 4, -46, 86, -17, -128, -79, 96, 22, -74, -12, 121, 80, -33, -17, -45, -28, 120, -63, 1, -54, 41, 1, 95, -55, 54, -43, 66, 10, -109, -128, -122, 113, -83, 126, -31, 105, -9, -97, 54, -112, 108, 69, 38, -47, -90, 107, 89, -31, -43, -99, -105, -85, -16, 95, -38, 124, -28, -115, 57, 126, 110, -45, -5, 27, 107, -12, 74, -52, -108, 60, -14, 32, -69, -84, -84, 49, 33, -54, -59, 63, 86, 108, -23, -48, -72, 82, -26, 100, 114, 51, -5, 120, -79, 12, 44, -90, 31, 39, 105, -54, -126, -29, -40, 110, 98, 84, 28, 35, -29, -6, 12, 38, 21, 37, -72, 123, -125, 42, -109, 56, -44, -15, -37, -125, -18, -90, -77, -32, 74, -16, -27, -36, -51, 79, 67, -62, -68, 79, -123, 31, 55, 105, 12, 53, 34, -30, -36, 85, -61, -96, -95, 105, -2, 49, -87, 105, -50, -78, 127, 89, -80, -50, 31, 68, -7, 39, -21, 37, -87, 25, 92, 87, -3, 40, 88, -44, 66, 47, -9, 37, -36, 12, -118, 5, -119, 66, 79, 70, -40, -49, -82, 0, -6, -58, 112, -78, 29, 108, -94, -109, 39, 127, 79, 7, -42, 13, -77, 38, -107, 98, -103, -91, -60, 90, -39, 45, 124, -80, 90, -121, -99, -10, 31, 59, -18, -23, -32, -4, 64, 90, -27, 116, -83, -47, -119, -96, -44, -25, 21, 19, 56, -118, -54, -35, -58, -68, -12, -64, 14, -86, 17, -111, 26, -23, 14, -79, 45, -50, 22, 79, -125, -126, -104, -115, -77, -99, -128, -80, 0, -105, -30, -78, 92, 30, -62, 12, -26, 0, 57, -6, 54, 65, -128, -30, -126, -103, -14, 39, 21, -38, 87, -103, -115, -73, 54, -20, -61, 101, 106, -84, 10, -119, 116, -7, -37, -14, 105, 70, 52, -52, -9, -109, -47, 0, 124, 77, -27, 30, 74, -61, 19, -86, -113, -4, 97, 78, 5, 15, -31, 4, 73, 30, 60, 11, -115, -128, -14, 51, 113, 105, 88, -30, -63, 44, 73, 103, 119, -86, -60, 10, -54, 1, -92, -40, -39, 64, -3, -32, -87, -109, -63, 12, 30, -69, 100, 120, -14, 11, -42, 82, -38, -56, -38, 61, 17, -114, 38, 104, -50, -108, -46, 117, 76, -24, -3, 8, -9, -62, -107, -42, 82, -61, 116, 70, -103, -61, -21, -79, 36, 62, -44, 61, 77, -109, 13, -16, -44, -72, 81, -1, -75, 63, -82, -88, 18, -10, -108, -52, 9, 70, -82, -28, -35, 33, 47, -97, 122, 31, -79, 37, 28, -89, -61, 59, 123, 95, 68, 14, -64, 72, -122, -45, 60, 9, 82, 80, 75, -44, 93, -99, -111, -84, 35, -55, 14, -98, -93, 12, -61, 8, -40, 106, 125, -47, -25, -77, -89, -111, -47, 9, 116, 16, -64, 96, -92, 53, 120, -41, -39, 14, 25, 122, -43, -71, -53, 13, -94, -114, -24, 69, 77, -15, -52, -92, -88, 107, 3, 115, -46, 8, 41, -1, -27, -28, -115, -12, -106, 100, -24, 3, -43, -23, 92, 95, 3, 47, 30, 42, 18, 34, -122, -85, 83, -49, 81, 21, -100, 11, -43, -120, 121, -80, 82, -119, -95, 111, -100, -95, -126, 52, -82, 82, 117, 87, -3, 13, -127, 19, 57, -70, 98, -89, -20, -92, -85, -100, 23, 5, -107, -18, 121, -126, 123, -118, 52, 14, -58, 106, 15, 16, -2, 121, -87, 93, -16, 12, 101, 62, 92, 38, 30, -31, 44, -37, 107, -43, 26, -2, 101, -2, 40, -5, -33, -97, -50, -101, -11, -23, -48, -26, 109, 52, -84, -97, -107, 77, 99, 68, 105, -108, 88, 39, -1, 71, 85, 111, 50, -4, 20, 90, 95, -71, 77, 29, -125, 29, -81, -46, -26, -84, 48, -113, -34, -23, -21, -2, 45, -18, -106, -77, -39, -62, -79, 96, -23, -36, 28, -85, -19, -16, -86, -3, -95, -127, 123, 17, 47, 122, -88, 102, -83, 42, -44, -68, -31, -69, -109, -78, 70, 101, 88, -41, -119, 103, 26, -75, 42, -124, 68, 36, -37, -41, -59, 44, 85, -75, -70, 77, 106, 118, -128, -97, -121, 71, -23, 124, -71, 27, -5, -16, 99, 127, -23, 90, 38, -51, 42, -90, -57, -33, -6, 91, 1, 109, 11, -35, -40, 88, 26, 33, -14, -75, -22, -1, 59, 51, 114, -65, 89, -79, -15, -79, -55, 0, 26, 108, -49, 45, 23, 15, -22, -94, -27, -24, 76, 110, 79, 35, -82, 95, -102, -88, -16, 81, 103, -3, -113, 64, 71, 77, 36, 126, -9, 51, 85, 53, -87, -55, -34, 23, 46, -54, -87, -114, -36, -124, -42, 68, -45, 104, 113, 59, 75, -9, 15, -74, -122, 50, 112, -103, -1, -126, 55, -88, -114, 27, -70, -74, -36, -52, 107, -11, -29, 72, 17, 45, -117, 81, -48, -51, 39, -45, 43, -127, -87, -6, -39, -67, -8, -9, -99, -74, 53, 89, -71, 96, 22, -115, -3, 42, 94, -84, 32, -62, -100, -94, 95, 59, 127, -5, 10, 80, -61, -19, -75, -14, 115, 83, -8, 13, -7, 127, -104, 73, 5, 47, -9, -102, -44, -79, -49, -5, -10, -41, 20, -122, 124, -3, 112, -54, -125, 91, 51, -30, 30, 115, 32, 60, -57, 14, 64, 87, -103, 35, 104, -39, -2, 5, 91, -32, -21, 27, 12, -75, -87, -12, 62, -25, -114, 71, 11, 76, 0, -86, 2, 35, -80, -86, -56, -108, 124, 1, -84, 75, 69, -6, -110, 71, -76, 18, -15, -15, -87, 108, -106, 114, -72, -97, 68, 87, -128, 45, 74, -5, 57, -77, -77, 125, 54, 74, 108, -53, 40, -26, 10, -93, 2, -36, -72, -74, -80, 15, 75, 0, 83, -11, 43, 71, -12, -105, -100, 109, -4, 18, -34, -102, -104, 2, 71, -24, 62, -91, 16, 47, 101, 125, -67, -117, -11, -44, -114, -46, -80, -113, 34, 70, 64, 94, 21, -93, 69, -74, 33, 25, -119, 103, -95, -111, 62, -25, 28, 21, 11, -52, -22, -117, 23, -42, 33, -41, -11, 88, 59, -12, -13, -13, 23, -91, 48, 56, -21, -70, -107, 48, 65, 24, -97, -101, -63, -12, 100, -44, -70, 110, -127, -66, 102, -91, 117, -52, -118, 79, 29, -123, 93, -35, -109, 106, -4, -61, 58, 98, -49, 102, -128, -19, -8, -34, -38, -123, 39, -80, 66, -126, 0, -12, 60, -88, 35, -82, -27, -5, -54, 25, 45, -44, 87, -25, 2, 36, -109, 112, 22, -50, 11, -91, 84, -39, -78, -61, 26, -49, -27, 71, -67, -89, 87, -45, 34, 100, -38, 59, -24, -79, 57, 59, 12, 27, 9, -96, -120, 23, -126, 54, -115, 63, 51, 89, -80, -43, 66, -109, -109, 50, 70, -64, -31, -40, 100, 48, -74, 118, 110, 86, 90, 107, 67, 103, 9, -78, 92, 115, 19, -124, 84, 29, 16, 65, 2, 29, 6, 115, -47, 56, 105, 83, 98, -123, 4, 119, -21, 122, 120, -98, -114, -15, 70, 93, -64, -27, -85, -26, 92, -113, -24, 53, 37, -127, 17, 60, -114, 94, 58, -9, 19, -8, 66, -70, 82, 25, -55, 71, 90, -29, -122, 15, 10, -16, 108, -15, 26, -90, -81, 93, -10, -123, 106, 108, 68, -2, 120, 36, 92, -105, 21, -32, -1, -116, 40, -102, 80, 96, -99, -111, 71, -101, -89, -90, -49, -16, -55, -10, 121, -24, 29, -113, -13, 68, -83, 67, -61, 74, 39, -29, 84, -9, -17, -95, -16, 13, 104, 18, 98, 38, -15, 19, 26, -86, 99, 30, 107, -30, -98, 74, 34, -55, 54, 97, 2, 10, -33, 54, 101, 101, 55, -66, 88, -21, -35, -23, 119, -108, 20, -112, -24, 109, 24, 100, 30, -51, -20, 118, -74, -76, -94, -78, 117, 70, -100, 73, 82, -26, 22, -79, 32, -108, 126, 105, 106, -9, 68, 11, 68, 1, -116, -55, -116, 55, 53, -101, 81, -47, 111, 72, -120, -73, -23, 121, 30, -24, -95, -5, -89, 107, 37, 89, -124, -84, 93, -94, -101, -49, 70, -77, -38, -51, 26, -123, -8, 73, 42, 59, -79, -15, 0, -100, 19, 1, -104, -15, 54, -128, 81, 110, 98, 49, -128, -10, -79, 123, -92, 5, -2, 72, 93, -45, -13, -55, 126, 21, -56, 84, 4, -81, -124, -115, 125, 83, -88, 117, 11, 15, -96, -122, -25, 74, -60, 83, 111, 15, -26, 123, -10, 73, -51, 34, -97, -120, 23, 0, 106, 101, 1, -96, -49, -93, -17, -32, -102, -92, -120, 41, 118, -10, -74, -59, -87, -102, 75, 118, -99, 21, -67, 120, 92, -67, -32, -117, 59, -47, -41, 61, 123, -87, 47, -81, -87, 16, -124, 93, -11, -17, -42, -18, 98, 41, 38, 72, -61, 121, 35, -39, 55, -11, 73, 125, 104, 7, 0, 41, 13, 62, 18, 10, 47, 81, 46, -45, -11, -60, -125, 36, 7, -46, 58, -20, 14, -51, 25, 67, -74, -82, 122, 79, -72, -122, -44, -6, -110, 2, -52, 113, -128, -55, 40, -6, -82, 70, -44, 20, -43, -91, 22, -18, -78, 73, 29, 2, 27, -98, 72, -36, -84, 84, 12, -97, -105, 8, -74, -12, 99, -124, 89, -22, 9, -19, 50, -48, 121, 0, 88, 66, -67, 89, 122, -99, -59, 1, 31, -75, -40, -64, 31, -9, 41, 31, -43, -6, 50, -56, 79, 26, 42, -30, 95, -75, 29, -66, -124, -67, -121, 52, -2, -101, -40, 3, -20, -77, 88, 29, 116, -66, -50, 36, -50, -81, -9, 107, 31, 82, 72, -60, 46, -11, -69, 52, 26, 116, -49, -26, -94, 76, -12, -120, 33, 13, -91, 6, -32, 116, -29, -55, 105, -107, 42, -53, 26, -69, -28, -26, -97, 6, -87, 24, -107, -56, -30, -4, -63, 68, 77, 55, 68, -41, -80, 77, 37, -99, 88, 35, -69, 12, -22, 75, 82, -34, 112, 3, -78, 92, 30, 15, -115, 55, 84, 98, 109, 75, 31, 85, -59, -38, -22, 126, -60, -55, 24, -16, -84, 32, -19, 89, 38, -1, 19, -30, -67, -3, -74, 17, 85, 25, 24, -59, -65, -120, 114, -106, -34, -124, -98, 81, -127, -121, 11, -119, 76, -76, -109, 119, -11, -81, 53, 71, -30, 107, 123, 79, -85, 40, 106, 109, -120, -91, -105, 3, 39, 41, 105, -5, -81, -7, 30, -27, 0, 4, -35, -98, -116, 117, -109, -48, 22, -21, -67, 37, -12, 50, -117, 117, 42, -102, -126, -52, -12, -92, 59, -47, 124, 106, 63, -23, -1, 36, 98, -113, 27, -128, -104, 105, 76, -112, 127, 75, 35, 37, -42, -46, -80, 18, -123, 38, 113, -84, -39, -118, 26, 7, 55, 81, -113, 23, -53, -75, -120, 38, 120, 74, 25, -21, -2, 85, -11, 91, -101, 47, 101, -32, 36, 85, -74, 0, 49, 15, 51, -76, -61, -108, 106, 43, 22, -18, -41, 82, -106, -46, 96, 0, 121, -77, 27, 49, -128, 96, -86, 83, 65, 119, -87, -122, -100, -67, 81, -53, -114, 42, -2, 82, -3, 6, -47, 63, 83, 122, -124, -46, -81, -45, 116, -37, -117, -40, -87, -11, 11, -126, -118, -88, -59, 16, 125, 86, -99, -79, 119, -127, -37, 50, 116, -124, -46, -62, -94, -46, 124, 85, 110, 39, 29, -21, -38, 106, 37, -17, -103, 69, -43, -8, -15, 0, -92, -63, 26, -34, 50, -61, -125, -121, -128, 43, 63, -95, -78, -85, 109, 101, -62, -12, -117, -99, 94, -80, -52, 3, 55, 127, -18, 63, -101, 35, 27, 121, 95, 118, -25, -122, -2, -38, 71, 62, -58, -28, -9, 117, 65, 50, 69, 111, -41, 127, -40, -83, -45, -67, 117, 86, -60, -94, 108, 99, 18, -118, 60, 83, 119, 32, 1, -54, -55, 75, 7, -13, -90, -67, -4, 23, 34, -110, 121, -60, 62, 50, -11, 97, 76, -115, -50, 38, 108, -11, -125, -48, 35, 95, 45, -74, 39, 94, 29, -71, -117, -2, -75, 103, -90, -47, -29, -70, -73, -85, -89, -31, -40, 120, -122, -55, -79, 33, -39, 22, 77, 19, -89, 108, 66, -23, -128, -116, -68, -93, 68, 13, 99, 125, 39, -86, -123, 44, -120, 13, 75, 105, -26, 72, -77, -121, 101, -54, 80, 43, 69, 116, 68, -58, -58, -18, -120, 75, -91, -20, 121, -84, 94, 48, 74, 47, 65, -68, 16, -23, 82, 63, 110, -46, -123, -80, -23, 99, -120, 109, -32, 20, 65, -127, 59, 69, -110, -92, -102, -103, 115, -46, -45, -6, -19, 44, -61, 110, 21, -28, -22, -93, 7, -116, -87, -45, -70, -68, -76, -31, 62, 7, 65, 118, 93, -63, -87, 101, -127, 108, -26, -32, 47, 31, -88, -62, 42, 37, 15, -47, 99, -64, 121, 83, -59, -82, -127, -35, 35, -51, 85, -30, 12, 62, 80, 94, -52, 119, -106, -78, 117, -18, 39, 25, -24, -75, -42, 45, -77, 100, -29, 116, 74, 60, 112, 7, -47, 69, -88, -28, -27, -101, -76, 48, 64, 42, -119, -12, -42, -4, 121, 90, 14, 83, -89, -113, -44, -57, 17, 113, -88, 77, 42, -106, -111, -106, 74, -127, 119, 16, -34, 94, -52, 64, 102, 5, -83, -33, 100, -3, -60, -18, 55, -101, -96, -50, -8, -93, 17, -13, -41, 97, -48, 66, -126, 36, 110, 77, 101, 70, 79, -6, -81, -35, 88, 97, -56, 70, -82, 61, 5, -74, 56, 21, -58, -114, -22, 73, 104, -98, 4, -93, -68, 18, 15, -14, 15, -64, -52, 63, 67, -36, 76, 105, 127, -54, -41, 20, -8, -77, -41, -34, 51, -37, 100, 57, 74, 47, -123, -113, -10, -29, 86, -124, -109, 89, -44, -65, 22, -89, -55, -115, -12, -95, -114, -75, -126, -53, -119, -100, -13, 47, -75, -50, 127, 0, 82, -31, 73, -67, -18, -105, -108, -60, -51, 104, 56, -12, -37, 15, -113, -97, -70, -96, -48, -127, -47, -33, 78, 8, -54, -55, -125, -3, 90, -124, -91, 107, -57, -115, -97, 108, 95, 30, -123, -97, 35, -13, 114, -18, 90, -61, -117, -127, -73, 69, 84, 116, 25, 6, 83, -45, 118, 20, -114, 106, 41, -125, -50, 15, -41, -9, -81, 21, -125, 28, -100, -110, 42, 98, -94, 50, 126, -104, -4, 22, 65, -40, -100, -27, -91, 30, -39, -18, 23, -70, -13, -48, 57, 118, -49, 61, 101, 2, -19, 61, 3, 49, -49, -72, 29, -122, -124, -91, -39, 113, 38, 64, -96, 22, 2, 13, 64, 18, -92, -35, -60, -45, -107, -50, -105, 64, -73, 51, 76, -7, 93, -48, -126, -79, 53, -25, 8, -1, 69, 8, -8, -62, 56, -29, -81, -114, -88, 99, 29, -6, 64, -27, -105, -6, -110, -12, 109, 4, -95, 121, -83, 95, -25, 23, -58, 121, 59, -77, 116, 17, 55, -62, -83, -2, -69, -15, 107, 82, -62, -79, 43, -68, 90, -86, 121, -7, 119, 11, -43, -127, 105, -62, 76, 5, -36, -34, -80, -22, 80, 63, -86, -119, 30, -74, 20, -106, -110, 116, 77, 91, -108, 44, -55, 105, 26, 99, -48, -99, 28, 88, 99, 51, 70, -1, -117, 127, -30, 126, 110, -34, -64, 11, 74, -37, 50, -101, 56, -73, 89, 51, -36, -56, 79, 87, -110, 21, 43, -47, -88, -60, 14, 108, -82, -42, -29, -80, 25, 15, 114, -12, 15, -34, 117, 85, -13, -117, -86, -69, -121, -43, -80, 59, 46, -17, -42, 111, 67, -55, -125, -44, 55, 102, 20, -126, -118, -42, -57, -115, 49, 19, -67, 25, 1, 16, 76, -25, -103, -47, -102, -101, -36, -98, -103, 100, 39, -5, -118, 73, -69, -9, 37, 92, 78, 68, -128, 95, -23, -121, -89, 114, 113, 84, 10, 100, 30, 73, -104, -97, 126, -25, -15, 71, -71, -2, 84, 82, 27, -70, -33, 34, -26, -26, 44, 78, -1, 121, 60, 33, 113, 46, -70, -53, 19, 81, 120, 78, -112, 88, -7, 33, -24, -30, 71, 31, -115, 22, -106, -35, -39, -93, -54, 124, 90, -25, -70, -128, -65, 121, -64, -88, -92, -16, 105, 61, 84, -85, 8, -69, -120, -29, 100, -64, 5, -93, 77, -97, -113, -66, -16, 122, -16, 56, -80, 51, 17, -46, -104, 32, 37, -91, 76, -24, -3, 82, 41, 58, -102, 18, -104, -21, -39, -99, -103, -114, 127, 56, -42, -27, -107, -36, 29, 23, 54, -81, 104, 81, -84, -59, -32, -127, -55, -26, 93, 76, -78, -122, 17, -56, 31, 73, -13, -70, -41, -74, -67, 80, 93, -46, 100, -72, 124, 3, -126, 86, -80, -110, 45, 115, 1, -41, 1, 35, 80, -73, -127, -37, -35, 104, -89, 66, 125, 114, -38, 106, -124, -59, -52, -91, -45, 82, 61, 37, -57, 40, 11, -23, -8, -79, 112, -10, -20, -93, -104, 72, 92, 68, 26, -72, 11, 31, -40, -51, 71, -100, -9, -93, 42, -109, -31, -87, -30, 17, -63, 106, -1, -65, 93, 85, -59, -119, -109, -26, 51, -54, 39, -65, -102, 64, 4, 109, -81, 103, 60, -25, -32, 53, -7, -33, -60, -7, -17, 81, 62, -128, 94, -17, 45, 93, -30, -99, 103, 115, -112, 72, 84, -38, -28, 56, 23, -103, 50, -13, -102, 14, 42, 117, 19, 24, -62, -34, -105, -94, -116, -42, -91, 57, 60, 55, -79, -51, 47, -105, -28, -6, -7, -111, -32, 43, -21, 123, 124, -53, -89, 79, 61, 96, 70, -38, -74, -98, 24, -86, -50, -77, -81, 79, 77, -56, 81, -99, -115, 4, -5, 24, 52, 6, -100, 97, -128, -43, -63, 116, 49, 94, -48, -90, 29, -79, -16, 120, 116, 121, 42, 45, -109, -100, 54, 86, 91, -56, 70, 39, -46, -51, 83, -105, -88, 96, -92, -79, -36, 117, -76, -68, 19, -9, -68, 35, 3, 107, 67, -86, -58, -42, -9, -90, 84, -67, -18, -26, 1, 65, 80, -124, 77, -12, 75, -88, -8, -100, 58, -39, -14, -33, 43, -15, -110, 69, 77, 80, 97, 37, 121, -125, 67, -67, -4, 127, -70, -108, 97, 60, -44, 127, 110, 93, 58, 19, -32, 35, 68, 6, -47, -115, 107, 1, -89, -91, 94, -28, -15, 86, -128, 48, 29, -3, -74, -91, -72, -81, -67, -68, -26, 106, -96, 99, -73, -43, 61, 61, -93, 109, -119, -77, 95, -44, -68, -28, 23, 60, -119, -50, 77, -16, 114, 126, 43, -72, 68, -84, 2, -30, 45, -110, -25, 37, 63, 120, 77, 99, 81, 6, -24, -74, -68, -70, 122, 51, 20, -63, -46, -43, 31, -12, -42, -48, 62, 12, -104, 115, -104, 27, 50, 24, 78, -78, -61, 1, -117, -12, -70, -1, -66, -116, -14, 65, -37, -71, -101, 105, 59, -124, 54, -84, 79, -62, 39, 46, 3, -70, 36, -12, 126, 126, 105, 22, -74, 2, 30, 62, -122, 39, -41, -47, 107, 81, -48, -107, -49, -32, -95, 48, 95, -123, -91, 11, -106, -72, 10, 4, 85, -71, 82, -114, 20, 38, -66, 25, -92, 67, 106, -8, -18, -63, 74, -31, 46, -89, 54, -93, -64, -75, 67, -104, -38, 113, 47, -32, 18, 126, -65, -30, -37, 111, -44, -62, -124, -30, 3, 54, -127, 123, -122, -64, 40, -80, 101, 120, 1, 29, 63, -11, 52, 41, 7, 25, 59, 83, -36, 9, 15, -116, -45, -24, 35, 9, -1, -111, 98, 52, 72, -87, 21, -45, -52, 38, -82, 41, -37, -101, 123, 14, 4, 55, 19, -49, -3, 111, 48, -28, 13, 57, -12, -93, -107, 123, -96, 45, -36, 38, 105, 35, 46, -10, 107, 125, 19, 48, -125, -81, -95, -9, -52, 13, 10, 81, 118, -18, 104, -80, -76, -98, -59, 57, -96, 104, 117, -122, -29, -111, 62, 63, -89, -15, -102, 35, 7, 89, -106, 60, 43, 84, 61, 108, -76, 3, 21, -125, 62, 124, -87, 22, -20, -127, -36, -127, -43, 9, -26, 66, 48, 5, -89, -36, 94, 36, 86, -101, 60, 115, 18, 43, -71, -13, 91, 44, -32, 47, 2, -123, -19, 11, -42, -128, -57, -119, -125, 58, 93, 89, 78, -52, 111, -128, -102, 122, 5, -42, 91, 17, -24, 41, 114, 94, -92, -109, 56, 86, -29, -46, 13, 121, 13, 110, -67, 89, 76, 32, -7, 101, -24, 64, 26, -24, 73, -8, 98, 92, -110, -22, -9, -9, -96, 99, -54, 60, -33, 113, -55, -78, 60, 24, 65, 101, -83, -3, -94, -119, 69, -81, -123, 9, 10, 61, 53, -126, -21, -10, 105, -116, 107, -91, -48, 8, 60, -6, -62, 109, 89, -125, 78, 74, 28, -1, 4, -11, 57, -37, -64, -6, -106, 32, -10, -95, -13, 0, -10, 56, 24, -93, -31, 52, 69, 15, 45, 15, 93, -115, 22, 30, 88, 59, -113, 15, -98, 54, 77, -23, 105, -58, -20, -83, -12, -91, 59, 32, 97, 36, -104, -23, -96, 43, -26, 66, -81, 37, -63, -15, 60, -41, 101, -53, -119, -7, 104, 47, 125, -107, -126, 46, -84, -26, -103, 62, -15, 52, 44, -60, -39, 121, -48, 127, -51, 108, 70, 56, 17, 62, 57, 73, 88, -71, -2, -92, 121, -14, 116, -25, -39, 49, 39, -11, 118, 121, 66, -2, -27, 98, -9, -72, 124, 94, -34, 47, 44, 15, -30, -85, 57, 89, 15, -120, -76, -125, 72, 81, -74, 53, -43, 114, -126, 20, 79, -62, -112, 64, -83, 13, 51, 10, -82, 123, -97, -125, -33, 63, -12, 42, 43, 40, -119, 115, 102, 18, 60, 48, -70, 0, -70, -69, -125, 80, 48, 101, 127, -54, 69, -33, 86, -68, -7, 26, -118, -80, -72, -77, 2, 18, -93, -60, -24, -60, 104, 94, 110, 47, -85, 25, -115, -23, 126, -41, -106, -52, 121, 95, 86, -16, 86, -68, 5, -96, 126, -93, 62, -53, -106, -76, -16, 26, -23, -33, -74, 63, 49, 57, 1, 115, -4, -99, 19, 57, 105, -118, -41, -54, -43, -117, 117, -23, 103, -46, -128, -99, -13, -5, -35, 5, 90, 18, 57, 120, -42, -38, 123, -12, 95, -72, 46, -49, 117, -56, -104, 109, 30, 123, -63, 103, -16, 2, -52, 2, -128, -68, -22, -12, -109, 116, -29, -45, 12, 51, 87, 72, 123, 97, -101, -42, 71, 10, -90, 114, 33, 10, -89, 110, 82, -102, -111, -44, -117, -58, 92, -88, -76, 114, 89, -116, -59, 117, -6, 126, -67, 64, 90, -68, -78, 93, 121, -80, -11, 117, 85, -6, 102, -73, 63, -54, 33, 73, 70, -99, -82, 39, 50, -25, -97, 9, 1, -27, 58, -54, -122, -70, -128, -29, 107, -23, 21, 63, 92, -82, 115, 64, -82, 61, -64, -39, 60, 3, 54, -13, 15, 124, 78, 3, -104, 106, -11, 41, -26, -124, 111, 15, -64, -18, -120, 110, 33, -26, -30, 90, 15, 72, 1, -125, -56, -6, -50, -46, -20, -123, 74, 4, 70, 77, 76, 33, -74, -56, -87, -3, -102, 99, -26, 114, 117, -6, -63, -39, 79, 20, 97, -53, -95, 70, -111, 112, -63, 119, 105, -44, -4, -14, -77, 70, 42, -70, 37, -128, 103, 117, 44, -30, -51, -32, 28, 119, 108, -118, -127, 74, -78, 64, -42, -2, 89, -50, 40, -83, -29, 33, -117, -34, 3, 70, 9, 21, -5, -123, 49, 15, 65, 51, 55, 23, -128, 98, -27, -103, -19, 52, -32, -20, -14, -48, -63, -37, -70, 111, -64, 115, -6, 118, -101, -50, 71, 107, -91, -64, -125, 18, -39, 102, -71, -14, -6, -121, 108, -22, -75, 31, -121, 45, 77, -116, 23, -57, 39, 92, -109, 115, -13, 52, -93, 43, -84, -105, 51, -101, 5, 95, -22, 50, -14, -98, -95, 88, -77, 47, 47, -126, 19, 10, -56, 98, -11, -127, -121, 28, -53, 1, 59, -5, 56, 19, 28, -90, 108, -12, 127, -91, 125, -23, 83, 30, -113, -78, -42, -121, -91, -30, -37, -127, 66, 25, -124, -9, 17, -19, 74, 110, -25, 41, 63, -124, -37, -39, -38, 123, -114, 103, 69, 75, 91, -106, -128, -5, -62, 5, -56, -13, 32, -117, -83, -103, -60, -66, -101, -81, 74, 48, 6, -8, 2, 67, -85, -48, -68, 122, -35, 65, 49, 38, 48, -3, -32, -114, -23, 110, 109, -67, -94, 59, 122, 107, 91, -34, -51, 76, -99, 17, 42, 4, -23, -104, 76, 83, -28, -116, 56, 67, -3, 105, -81, 20, 31, 123, 106, -40, -108, 50, -112, 94, -37, -44, 121, 4, -79, 4, 27, 35, 31, 55, 115, 102, -58, 45, 127, 65, 110, 89, 19, 124, 57, -50, -107, 109, 71, -48, 9, 87, -69, -119, -16, -111, -104, 30, -2, -76, -106, 12, -41, 63, -89, -80, 84, -30, 125, -57, 121, 64, -73, 19, -6, 22, 8, -82, -1, -10, 53, -2, 1, -109, -34, -73, 54, -100, 25, 108, 73, -48, 69, 119, 0, 20, -54, -58, 94, -36, -5, -19, -118, 5, 103, -51, 38, -69, -81, 120, -117, 18, 23, 22, 11, -120, -36, -37, 73, -96, 104, -110, 18, 95, -20, -115, 43, 31, 94, -57, 8, -101, -67, 21, 123, -107, -97, -74, -77, 45, 95, 83, 5, 119, -54, -101, -78, -81, 63, 30, 97, 126, 0, 118, 20, -59, -110, -65, -47, 35, -60, -72, -64, 123, -90, -121, -84, -40, -70, 50, -103, 49, 121, 34, 73, 3, 42, -53, -87, -122, 48, -12, -79, -68, -1, -43, -62, -68, 60, -64, -120, -33, -73, 89, -11, 60, -46, 7, -31, -116, -47, 68, 0, 126, -3, -102, -1, -9, -63, 121, -102, -15, 51, 124, 79, 35, -7, -39, 10, -110, -3, 79, 62, -27, 78, 97, 56, -111, 116, 66, -115, 42, 43, 71, -90, -15, -62, 3, -36, -99, 112, 54, -17, -72, -77, -85, 74, -84, 12, 97, 72, -11, 74, 103, -35, -56, 34, -30, -17, 110, 16, 90, -121, -7, -65, 122, -113, 98, -75, -67, -27, 73, -47, -39, -54, -110, -33, -44, 16, -22, 117, 92, -4, 120, -62, 101, -42, -81, -45, 111, 81, -7, -46, -64, -67, 101, -54, 126, 11, -39, -116, 114, 13, 35, -67, -49, -128, 41, -17, 45, 119, -101, -55, 69, 68, -42, 66, 86, -8, -101, 83, 25, 6, 83, 87, -92, 53, -35, -17, -94, 8, -42, 97, -25, -105, -76, -15, 123, 38, -66, -44, -124, 76, -34, 3, -41, 23, -8, 108, -87, -86, 2, 101, 19, 7, -95, 45, -37, -13, -12, -114, -66, 85, -54, 109, 60, 20, 8, -67, 21, 59, -31, -112, 27, -93, -102, -36, 84, 82, 123, -21, 41, -13, -1, -128, 107, -118, -86, 43, 79, 98, 63, 47, -24, -65, -120, 0, -8, 39, -96, -1, -78, 1, -91, -22, 54, -117, -75, -38, -8, 62, -14, -100, -71, 40, -123, 127, 117, -82, -89, 122, 102, 86, -20, -11, 102, 106, -77, 15, 39, -18, 109, -107, 114, -121, 51, 103, -82, -14, -25, -33, 23, 29, 19, -52, -17, -47, -117, -123, 51, -100, -64, 42, 37, -42, 90, -1, -66, -99, 37, -60, 100, -100, 18, 28, -74, -69, 92, -1, 50, -82, 97, 4, 100, -111, -105, 28, 7, -80, 87, 126, 100, 110, -30, 117, -42, 30, 105, -73, 14, -46, -90, 89, -96, 86, -123, -82, 48, -93, 40, 77, -3, -7, -109, 103, 89, -7, 23, -81, -34, -7, 104, -106, -91, -40, -96, -81, 73, -58, -3, 115, -32, -94, -93, 106, 126, -67, -70, 72, -5, -64, -106, 88, -33, 105, -47, 23, 119, 36, -53, -37, 72, -1, -38, 97, 79, 91, -82, -94, -76, 29, -19, 93, 73, -86, 110, 29, -54, 65, 5, 112, -128, -8, -50, 117, -65, 100, -83, 37, 116, 50, -117, 74, -86, 92, -91, -85, -40, 59, -50, -76, -18, 39, -79, -36, 56, -24, 122, 66, -102, 53, 98, -21, -81, -54, -55, -76, 121, -109, 6, -81, -7, -88, 41, 103, 22, 51, -61, 77, 118, -70, 7, -127, 97, -52, 85, 23, 80, -83, 113, -63, -33, -80, -3, -25, -48, 115, -44, -93, 4, 10, 36, 57, 123, -79, 92, -86, 20, 65, 111, 56, -83, 21, -95, 63, -109, -49, 90, 93, -11, 44, 110, -36, -31, 50, -121, 15, -68, 101, 27, 124, -127, -81, 68, 14, 81, -83, 71, -109, 122, -62, -97, 4, 121, 84, 90, 73, -3, 77, -73, -123, 48, -122, 52, 114, -65, -23, 13, 98, -8, -111, -38, 58, -13, -90, 69, -121, 90, 82, 114, 39, -12, -51, 85, 86, -14, -28, 94, 65, 81, 72, -95, 66, -64, 33, -89, -77, -21, -78, 121, -91, -104, -43, -119, -13, -78, -78, -34, 59, 98, 115, 3, -4, 82, 7, 37, 66, -53, -110, -103, -112, -24, 14, -40, -25, -108, 56, -100, 22, -108, 52, -113, 126, -6, 122, 4, 0, -73, 111, -90, 18, -76, 73, 38, -58, -50, -40, 46, 110, 61, -59, 97, -22, -50, 35, 42, -61, -40, -29, -60, 50, 127, 88, 47, -51, 22, -108, -22, 53, -123, 101, 89, -95, -12, -86, -87, -53, 116, 3, 120, -50, -104, -19, 27, -126, 30, 21, -42, 52, 59, -127, -109, -9, -91, -77, -82, 124, 79, 48, -53, -22, -114, -127, -4, 86, -111, -59, 53, 48, -57, 78, 110, -40, 119, 105, -77, -70, 23, -95, -70, 32, -18, 8, -48, -63, 22, 88, 1, -18, -113, 55, -58, 24, -94, 6, -90, -18, 73, 75, 49, -120, -14, 114, 73, -3, -2, -109, -53, -51, 72, 41, -120, 88, -52, -43, 0, -108, -11, -28, 94, -115, 93, -7, -18, -75, 108, -8, 83, -28, 117, 55, 46, 40, 111, 64, -30, -68, -40, 37, -127, -110, 67, 38, 15, 95, 9, -74, 122, -72, 45, 22, 82, -110, -76, 9, 106, 69, 93, 7, 85, -81, -26, -112, -125, 50, -106, -88, -27, 58, 98, 15, -44, 8, -101, -2, -55, 56, -51, 44, -115, 111, 9, 34, -121, 23, 59, 38, 95, -49, -13, 98, -127, 27, 125, 79, 34, 9, 108, 75, -30, -106, -87, 25, -63, 5, 9, 63, 91, -17, -128, 83, -40, -114, 113, -72, 100, 79, 118, 68, -33, -38, 15, -101, 72, -46, -120, -62, -14, 25, -62, -105, 69, -48, 41, -25, -5, -60, -120, -3, 72, 0, 39, 54, -101, -28, -13, -13, 21, 16, -26, -77, -80, -14, 15, 37, 48, -63, -80, 33, -35, -53, 89, -127, -117, -26, -96, 48, -22, 80, 110, 46, 93, 6, 0, -105, 35, -119, -85, 4, -53, -128, -45, 1, 19, 45, 26, 94, 51, -35, -50, 6, -24, 99, 118, -71, -102, -68, 89, -6, -119, 122, 65, 46, 23, 24, -126, 49, 35, -34, 71, -117, -30, -22, -27, -18, 22, 28, 44, -15, 25, 57, -121, 109, 78, 27, -126, -115, -63, -48, 47, -78, -112, -46, -44, -82, -110, 81, 55, -40, -14, 5, -96, -86, 87, 2, 82, 83, 50, 89, -4, -25, -110, -8, -99, -106, -16, 32, 16, -102, 101, -70, 96, 40, -105, 90, -98, 7, 6, 67, 74, 28, 19, 99, -32, 32, 54, 8, -81, 46, 103, 24, 88, -112, 55, 110, 8, -12, 122, -82, -92, -68, -96, 109, -64, 49, 69, 75, 117, -75, 92, 68, -47, 33, 20, 19, -89, -18, 110, 43, 67, -91, -26, 9, -103, -92, 77, 22, 126, 0, 37, 31, 116, 6, 29, -90, -65, 103, 33, -60, -67, 38, 19, -43, -35, 91, 48, 70, -114, -22, -35, 6, -122, -65, -15, -111, -26, -27, 1, -118, -82, 108, 89, -84, -41, 122, 48, -30, -18, -110, 12, 34, 27, -24, 87, -78, -112, -78, -128, -53, 74, -127, 101, -12, 60, 3, 56, 127, -39, 96, -16, -74, 110, 44, -96, -51, -11, -39, -113, 98, -37, 97, 36, -119, -80, -88, 31, -4, 11, -19, 59, -84, -121, -70, -79, 97, -25, 22, -8, -79, -60, 39, -108, -79, -72, 46, 124, -9, -18, 121, -93, -128, 95, -98, -24, -17, -79, 62, 95, 64, -55, 85, 70, 116, 41, -8, 35, 18, 82, 15, -13, -106, -92, 96, 84, -17, 102, 75, -33, 6, 74, -108, 56, -46, -77, 60, -47, -31, 112, -23, -64, 27, -15, -126, -94, -72, -86, -48, -73, -49, 99, -23, 66, -108, 109, 8, -28, -105, 73, -7, 109, 85, 31, 66, -128, -4, 42, -61, -18, -61, -122, -4, 69, -80, -119, 93, -89, 119, -128, 113, -76, -98, 99, -115, -55, 105, 72, 25, -87, 40, -98, 79, -117, -87, 32, -77, -45, -37, 73, -105, 74, 113, -6, 38, -113, 66, -25, 45, 19, -77, 51, -29, -15, -79, 42, 50, 43, -25, 94, -92, -116, -28, 78, -96, -17, 42, -81, 68, -124, -43, 91, -25, 115, 5, 33, 40, 59, -33, -69, 18, 57, -39, 117, -45, -18, -90, -108, -67, 11, -116, 112, -99, -77, -67, -55, -127, -109, 48, 76, 15, -85, 65, -29, 79, -102, -74, -12, -42, 18, -73, -66, -122, -40, 61, -59, 63, 46, 121, 27, 104, 23, -3, 87, 112, 78, 87, -66, -26, -61, -42, 24, -52, 40, 90, -5, 18, -34, -47, 25, 9, 7, -79, 116, 102, 110, 95, 0, -68, -1, 56, 61, 11, -127, 60, 107, 117, 89, 10, -49, -115, 89, 62, -32, -14, -10, -110, -59, -51, -113, 75, -120, 48, -17, -97, -58, 106, -81, 22, -27, -46, -121, -75, 88, 29, -103, -3, 73, -38, 22, 96, -79, -47, 84, 72, -77, -73, -41, -75, -50, 81, -106, 79, 70, -45, 97, -121, 62, 70, 9, 71, 8, -116, -29, 67, -90, 69, -89, -16, 84, -12, -38, 64, 95, -34, 98, -45, 109, -52, 70, 28, -1, 25, -46, 120, -86, 86, 4, -21, 29, -42, 20, -42, 22, 11, 49, 76, 24, 113, -71, 35, -117, 7, 50, 64, 9, 105, -77, 108, 87, 93, 59, -124, 45, -82, -49, -38, 79, -88, -5, -41, 108, -15, 42, 29, -126, -97, 4, 42, 45, -106, 114, -50, -112, 122, 22, 31, -9, -56, -103, -98, 116, -127, 17, -14, 70, -10, 22, 123, 78, 114, -43, -10, 7, 57, -108, -5, 28, 118, -6, -12, 52, 25, -115, -112, 78, -109, 104, -24, -15, 29, 55, 6, 120, -2, -63, -74, -91, 115, 124, -127, -29, -119, -32, -23, 66, -11, -125, 104, -60, 106, 17, -69, -45, -67, -39, -8, 99, -10, 40, 72, -122, 126, 103, 10, 93, -30, -49, -105, -67, -41, 71, -43, -9, -124, -89, -66, -55, 11, 45, 79, 68, 48, -128, 40, 39, 3, 62, 40, 77, 51, 73, -90, -89, -23, -48, -37, -64, 56, -83, 119, 29, 57, 86, -111, 65, -21, -117, 59, 53, 22, -72, 117, -65, -22, 67, -86, -26, -93, -50, 103, -87, -65, 69, 80, -85, -67, -40, 106, 95, 10, 55, -98, 83, -35, 124, 110, -60, 61, -16, -92, 101, 29, 103, -106, 116, 114, 98, -23, -99, -19, -54, 60, -112, -56, 42, 87, 88, 123, -93, 0, -87, 15, -45, 81, -21, 51, 113, -91, -93, 107, 13, -1, -86, 62, 23, -8, 4, -58, 94, -65, 90, -37, -23, 109, -71, 124, -109, 99, -76, -45, -14, -76, 82, 42, -91, 62, 89, -80, -118, -105, 75, -77, 115, -54, -102, -101, -60, -18, -18, 33, -19, -19, -22, -12, 104, 97, 31, 46, 91, -128, -6, -41, -108, 80, -96, 57, -117, -36, 31, -109, 41, -123, 106, 5, -58, -88, -14, -102, -44, 60, 52, -22, -8, -116, -29, 38, -106, -22, -118, 83, 7, -23, 86, -69, -25, -76, -84, 41, 82, -20, 6, 124, 5, -113, -59, -56, -103, 30, -84, -60, 47, -109, -83, 0, -128, 58, 4, -41, -126, 18, -87, -78, 91, 57, -23, -81, -56, -83, 29, -19, 106, 75, 33, 75, 117, -49, -98, 41, 4, 8, 48, -61, -21, 92, 73, -51, -53, 23, 123, -25, 45, 59, 49, 40, -37, -56, -3, 122, 73, -123, -108, 127, 115, -46, 3, -104, 126, 72, -38, 69, 18, -99, -70, 59, 110, 2, -127, 3, 6, -102, -41, -43, 90, 47, -102, 3, -84, 27, -87, -121, 80, -43, -74, -26, -93, -70, -23, 39, 14, -23, -94, -78, 5, -32, -1, 73, -105, 90, 88, -47, -6, -83, 68, 36, 6, 72, -74, -106, -103, 27, 40, -3, -127, 92, -53, 107, -20, -127, -78, 83, 14, 62, 41, -117, 28, 61, 74, 105, -56, 88, 2, -65, 98, -33, -47, -66, 111, -100, -98, -119, -68, -103, -62, -17, 63, -103, -89, 1, 113, 49, 24, 27, -11, -18, 61, -111, -80, -10, 6, -85, -15, -74, -17, -26, -123, 104, -88, 49, 116, -110, -50, -93, 30, -27, -41, -81, 101, -88, -4, 32, -36, 50, -106, -3, 51, 5, 89, 31, -121, 44, -67, -84, -6, -25, 18, 55, -76, 98, -77, -81, 61, 67, -66, 85, 90, 105, -12, 126, -29, 45, 1, 18, -118, 103, 120, 50, -123, -105, 7, -70, 38, 46, 32, -123, 127, 65, 65, 13, 4, -27, -96, 32, 79, 4, -94, 78, 83, 36, -101, 5, 119, -86, 111, -96, -118, -3, -94, 38, 88, -47, 26, 56, 9, -98, 40, 86, 3, 96, -117, -25, -121, -1, -65, -55, -105, 78, 89, -2, 111, -29, 115, -103, -31, 1, -99, -116, 64, 121, -7, 107, 17, 96, -63, 18, -117, 55, -83, 52, -8, -10, 15, 25, 50, 17, 79, -87, 18, 60, 70, -119, -59, 33, 14, 55, 15, 99, 48, 28, 39, -105, 68, 22, -4, -63, 62, -45, 108, 112, -55, -95, 17, -14, -79, -117, -121, -3, -66, 124, 89, 18, -80, -102, -103, 105, 105, -82, -38, 34, -104, -73, -90, -123, 51, 75, -34, -114, 116, -81, -119, -5, 81, -9, 38, -111, 54, 71, -79, 66, 33, 30, -102, 71, -119, 62, -106, -105, 85, 60, -78, -83, 82, -115, 46, 87, 105, -79, 99, 24, -69, 41, -19, 107, 71, -109, -85, 29, -5, -26, -87, 13, 31, -37, -96, 37, 7, 2, 43, -11, 2, 112, 28, -51, 61, 56, 0, 10, 13, -70, -85, -88, -21, 58, 70, -111, 71, 106, -112, -50, -90, 15, 91, -93, 70, -14, 11, -20, 45, 15, 29, 47, 127, 47, -41, -85, 58, -49, -104, -22, 77, -93, -76, 122, -101, 58, -2, 73, -116, -124, -8, -69, 108, 35, 115, 73, -91, -18, -13, 1, 8, 71, -94, -113, -92, -102, 30, 64, -89, -40, 65, -60, -77, -101, -38, -94, 85, 77, 83, 14, -98, -16, -5, -111, 117, 71, -102, 66, 102, 48, 21, -32, -36, 98, -104, 22, 21, -33, 8, 44, 46, 98, 58, 48, 38, 119, 92, -23, 66, -21, 28, -12, 71, -19, -66, 36, -40, 15, -71, -35, -110, -89, 31, 74, -52, 41, -28, 31, 107, -115, 88, -46, -70, 79, 90, -58, 32, 76, 67, 87, 112, 69, -35, 98, -116, -45, -15, -2, 66, -119, -80, -53, 10, 87, 116, -73, -53, -91, 84, 11, -115, 57, -29, 71, 56, -52, 120, 65, -34, -45, 0, -21, 0, 97, 41, -89, -18, 10, -86, 119, -11, -103, -37, -97, 113, -58, -84, -56, -113, -21, 72, 56, 63, 8, 14, 57, -9, -39, 6, 50, 95, 44, 26, -103, -86, -28, -84, -127, 32, -74, 22, 67, 95, 54, 116, -80, 120, 114, -3, 86, -34, -91, -102, 113, 64, -97, 111, -5, 17, 101, 48, 117, -6, -2, 109, -105, 12, -75, 9, -123, 72, -17, 105, -110, 57, 68, 70, -61, -38, 40, -123, -97, 36, 87, -31, 68, 120, 21, 71, 26, -59, -55, 14, 118, -21, 119, -68, 68, -39, -11, -96, -62, 89, 45, -55, -80, -126, -104, -112, -9, 52, -127, -112, -118, 19, -18, -75, 93, 107, -50, -47, -72, 40, -66, 62, 126, 47, 45, -121, 121, -37, -3, 69, -81, 63, -14, -65, -124, 83, 108, 52, 116, 115, 67, 16, -81, -41, -11, 9, 80, 111, 64, -61, 3, 20, 90, -43, -90, -33, -11, -68, 107, -25, 56, -3, -4, 100, 27, -59, 23, 13, -115, -28, -14, -55, 109, -39, 22, 54, -17, -25, 45, -15, -95, 104, 109, 126, 33, 125, -101, 101, 42, 70, 80, 24, -99, 127, 110, 45, -37, 20, -65, 65, -67, 107, 35, 75, -56, 36, 122, 25, -75, 22, -16, -95, 7, 111, 40, 41, -8, -54, 16, -82, 1, 127, -96, 69, 17, 60, 63, 101, -83, 34, -21, -118, 100, -94, 95, -21, 106, -54, 72, 55, -24, 47, 79, 116, -41, -122, 5, 7, -109, 46, 15, 118, 22, -15, -55, -9, -42, -25, -3, 8, -126, 68, -57, 125, 84, 49, 0, -5, -98, -117, 107, -11, -86, 120, 73, 74, 0, -49, -104, -37, -28, -105, 26, -107, 60, -103, 96, 126, -45, -80, 105, 19, 113, 114, 99, -22, -109, 111, 7, -39, -80, 10, -72, 86, -17, 6, -1, -107, -99, -65, -15, -51, -112, 120, 119, 121, -93, -88, -20, -112, -103, 15, 116, -122, -46, 20, 25, -107, 99, -121, 33, 38, 48, 114, 56, 44, 67, 29, -30, 110, -41, -97, 103, 29, -45, 50, 112, -70, -115, -117, -47, 39, 40, 3, -33, -8, -103, -87, 68, 9, -5, -2, 26, -49, 23, 71, 89, -49, -102, 84, 71, 26, -96, -80, 39, 35, 70, 56, -49, -21, 50, 3, 81, 61, 98, 15, -71, -70, 12, -31, 68, -76, -107, -115, -72, 28, 7, 97, -3, -17, 124, 27, -39, -87, -44, -88, 63, 119, 38, -10, 94, -75, -51, 113, -126, -54, -7, -71, -30, 105, 24, -37, 51, 7, 102, -98, -114, -125, 41, -81, 65, 117, 92, -101, 123, -19, -41, -108, 81, 105, -123, -70, -7, -3, -109, 114, -47, -100, 46, -48, -122, -14, 54, 98, 67, -79, 95, -3, 17, 90, 56, 70, -18, 79, -75, 23, -87, -95, 24, 37, -105, -87, -85, -120, -67, 4, 81, 16, 25, -3, -3, 123, 110, 47, -10, 47, 24, 8, -10, -49, 61, -122, -103, 69, -11, -58, -8, 97, -77, -35, 69, -66, 121, 118, -63, 97, -41, 51, 120, 22, -38, -126, 69, 88, 1, 68, -76, -102, 74, -30, -6, -48, -92, 59, -118, -14, -31, 27, 104, 119, 94, -81, -78, 1, -81, -50, -117, -39, -25, -76, 54, -40, -14, 57, -120, -86, -12, -108, 61, -59, 127, 92, -34, 83, -102, -122, 26, 111, -85, 6, -61, -116, -32, -56, -127, 96, 43, 63, -102, -18, -45, 110, -85, 25, 86, -109, 4, 46, -70, -100, -96, 5, 38, -63, 90, -126, 66, 89, -10, 78, 72, 124, 40, -112, -97, -110, 0, 126, -110, -7, 36, 31, -58, 80, 75, 53, 39, -9, -34, -2, 79, 84, -28, -23, -90, -76, -44, 25, -93, -38, -27, 55, 78, 87, -45, 113, -52, -123, 44, -66, 46, 80, -38, -108, -21, 52, -7, 25, 108, -92, -60, -71, 94, 44, 113, -89, -47, 30, 42, -100, -79, -119, -38, -14, -121, -100, -59, -79, 71, -127, -116, 121, 13, 12, 87, -6, 82, 63, 56, 49, 84, -84, -45, 15, -65, 73, -35, -125, 103, 76, -53, 57, 82, -109, -2, 5, 45, -16, 109, 52, 98, -76, 18, -32, -80, 24, 48, -74, -53, -65, 75, -2, 31, 21, -61, -90, 48, 6, 126, 51, 80, 22, 111, -89, -116, -35, 60, -20, -47, 33, 0, -127, -73, 63, 2, 60, 57, -2, 104, 107, 53, -26, 81, 20, 110, -108, -107, 64, 35, -84, 14, 101, -59, -113, -47, 57, -35, -7, -61, 47, -62, -15, 61, 78, 23, -95, 0, 27, -78, -5, -46, 36, -32, -12, -116, 3, 54, 46, 93, -6, -6, 13, -73, 50, -102, -37, -76, -96, 0, -13, -125, 44, 76, 91, -7, -93, 70, 72, -60, 95, 112, 86, 2, 86, -72, 8, -7, -91, 88, 34, -16, -105, -119, 78, 28, -25, -34, -20, 63, 63, -125, 84, 87, 124, -58, 118, 114, 64, 62, 34, -94, 118, 22, -80, -108, -103, -85, 39, -61, 124, -36, -116, -112, 32, 47, 96, -116, 76, 19, -23, -65, -112, 78, -14, 36, -118, 91, -12, -1, 71, 6, 6, 37, -20, 29, -108, -101, 84, -94, -40, 16, 16, -113, 62, -32, -12, -42, 25, -72, 62, 124, 85, 101, 62, -111, 67, 62, -70, -113, -106, -9, 86, -15, 1, -56, -33, 74, 95, 55, 25, -83, -92, -20, 66, 69, -60, -59, -48, 20, 26, 43, 49, 62, 42, -69, 78, 111, 81, 127, -4, -97, -77, -124, -65, -60, -125, -28, -127, -70, -53, 60, -97, -11, 71, 34, -45, -128, -1, 123, 20, -73, 71, -4, 35, -10, -25, 49, 98, -19, -85, -123, 42, -90, 57, 56, 114, 64, 106, 34, 110, 44, 29, -109, 62, 97, -68, 72, 106, 53, -50, -14, 116, 109, -85, -30, -106, 51, 127, 35, 62, -81, 108, -61, -99, -84, 118, -114, -35, -93, 14, 123, -94, -15, 4, 56, 17, -127, 103, -123, -111, 13, 60, -41, -79, -65, 95, 89, -73, 116, -18, -125, 70, -91, 102, 47, 86, 59, 21, 106, -84, -37, -25, -64, -115, -92, -21, 37, -14, -123, 19, -86, 111, -75, 27, 113, 19, -7, -7, -68, 48, -97, 78, -103, 25, 23, -84, -52, 5, 12, -94, -76, 14, 40, 65, 76, 16, 123, 118, -54, -31, -110, -49, -82, 107, 18, -46, 4, 107, -4, -123, 13, 101, 91, 102, 42, 100, 20, 108, -21, -13, -4, -114, -16, 57, 123, 42, 114, 31, -82, -119, -73, 78, 15, -17, -84, -91, 50, -6, 89, 76, -53, -42, 101, 74, -89, -29, 52, -128, -32, 39, 21, -46, 58, 79, 71, -99, -126, 55, 113, -113, 37, 52, -81, -18, -124, 50, -24, -24, -36, 101, 59, -7, 2, 28, -83, -81, -127, 57, -102, -107, -44, 17, -43, 111, 113, -102, -108, -62, -53, -59, -37, -128, 41, 105, -15, 111, 73, -13, 85, -6, 62, -107, 0, -119, -35, -39, 18, -21, 105, 113, -110, 111, 4, -92, -53, 9, 48, 120, 44, 72, 75, 123, -42, 9, 86, 122, 42, -80, 55, 75, -40, -125, 3, 31, -109, -37, -47, -91, -17, 21, 117, 71, 67, -113, -84, -27, 11, -21, 32, -51, -29, -101, 82, 30, -84, 13, 123, -97, 46, 0, 53, 46, 9, -42, 34, -128, -100, 7, -19, 95, -27, -79, -21, 71, 10, 3, -70, -92, 43, 109, 76, -38, -69, -28, 68, -16, 55, -126, -35, 116, 120, 59, -19, 108, 72, 67, -56, -91, -43, 81, 101, -30, 69, -49, 88, -87, 82, -55, -111, -124, -71, 45, -38, 31, 62, -95, 25, -99, 62, 19, -99, 81, -30, 115, 118, 52, 102, -89, -39, -30, 17, -83, -94, -11, -33, 69, -16, -128, -3, -126, -65, 33, 115, -25, -52, -41, 112, -122, 48, -28, -8, 108, -37, 44, 71, 58, 99, 112, 55, -17, 104, -68, 37, 13, -3, -16, 113, -128, -64, -1, -112, 80, 51, 50, 10, -62, 11, -113, -94, -67, 33, -121, -93, -6, -80, -12, -90, 76, -81, -13, 13, 19, -52, -96, 71, 96, -29, -63, 43, 116, -33, 12, -73, 63, 29, -119, 57, 46, 126, 117, -45, 58, -89, 52, 86, 105, -40, -36, 67, 50, -82, -14, 75, 102, -93, -30, -53, -120, 83, -59, 99, 89, -105, 102, -3, -65, 27, 66, -1, -103, -115, -37, -100, 97, 108, -82, -5, -10, 38, -64, 77, -124, 110, -54, -27, -16, -68, -115, -95, 19, -65, -27, 73, -22, -109, 46, 76, -35, 101, 125, 104, -32, 21, 79, -59, 71, 42, -79, 115, -46, 4, 6, 95, -125, 102, 121, -55, 30, -36, 71, -123, -125, -126, 47, 112, 31, -80, -124, -13, 126, 6, 117, 39, -6, 2, 98, 68, -20, -64, 32, -17, -62, 31, 110, -103, 98, 92, -69, 78, -7, -94, -7, 41, -4, -23, 83, -84, 124, 99, -115, 16, 16, -79, -65, 12, 69, 71, -60, -78, 105, -66, 43, -114, 53, -73, 99, -20, 22, 125, -107, 47, -111, 126, 25, 55, 121, 120, 120, -52, 87, -119, -22, -66, 112, 68, 96, -109, -118, -44, 125, -72, 69, -57, -91, 34, -60, -117, 36, 127, 68, -84, 43, 18, -27, 35, -116, -12, -94, 9, -78, 83, 127, -43, 109, 7, 61, -98, 8, 25, -39, -4, -91, -1, 45, -42, -87, 24, -58, 107, -103, 79, -40, 115, 51, 53, 92, 18, -66, -112, -14, 109, 100, 60, -35, -91, 41, -63, -28, -53, -100, -106, 70, 107, -78, 88, -97, -57, -96, 127, -25, -127, -50, -119, -101, 69, 101, 28, 94, -30, -47, -125, -38, 12, 9, 83, -108, 17, 107, -109, -46, 15, -19, -13, 105, 108, -97, -88, 34, -117, -96, -90, -103, 123, -59, 84, -74, -87, -17, -8, 11, 36, 107, -24, 38, 24, 73, -57, 81, -28, 75, 59, -87, -119, -58, 110, 125, -29, 110, -66, 108, -90, -31, 41, 118, -44, -67, -127, 67, -11, 83, -48, -127, -116, 10, -33, -85, 85, -46, 26, -54, -37, 112, -26, -117, 79, 25, 1, -27, 96, -100, 49, 126, 111, -37, 14, 58, -124, 78, -33, 7, 34, -110, 71, 30, 91, 104, -118, -12, 112, 117, -102, -5, 105, -45, -31, 26, 13, -115, -18, 46, 45, -69, 69, -66, 66, 62, 88, 67, -107, 64, -126, 29, 76, 17, 107, 23, -120, 82, -122, -3, -62, -56, -75, -24, -119, -119, 54, -12, -109, 82, 25, -101, -106, -86, -83, 33, 62, -39, -122, -68, 53, 19, -118, 118, 69, 94, -78, -27, -54, 65, -127, 55, 52, -36, 9, -38, 72, 119, 35, 47, -94, 6, 38, 78, -45, -51, 7, -49, -99, -99, 71, -19, -10, -81, 5, 34, 37, -26, 23, -55, -14, -21, -66, -113, -50, -19, 111, 92, -15, 122, 82, 0, 106, 124, 107, 84, -8, 61, -77, 62, 110, 38, 112, 30, -73, 114, 58, -18, -35, -38, -117, -97, 111, 33, 50, 53, -40, 9, 14, 9, 37, 82, -20, 9, 76, 86, -59, 72, -58, -109, -57, -19, -27, 33, -7, 47, -54, -45, 29, -95, -38, -58, -51, -43, -58, 94, 74, -7, 75, -39, -43, -37, -67, 45, 14, -26, 44, -38, -115, 80, 84, -109, 10, -32, -19, 56, 43, -49, -35, -38, 58, -11, 87, 74, -87, -111, 117, 77, -8, 105, -5, 73, 108, -67, -75, 117, -44, 36, 43, -92, -72, -84, 73, -118, 120, -104, 90, -23, -89, 78, 91, 30, -14, 74, -93, 73, -5, -5, 48, -29, -31, -122, -49, -52, 91, -126, -114, 111, 44, 120, 56, -116, -123, 83, -86, -40, -42, 33, 124, -44, 40, -126, 46, -54, 5, 86, -49, -105, -4, -64, -23, -13, -19, -72, 35, -35, -93, 57, -58, 40, 112, 72, -100, -120, -2, -63, -15, 124, 6, -7, 20, -44, -1, -19, -31, -55, 73, -4, 53, 91, -8, 17, -28, -121, -96, 36, -7, 39, -69, -87, 48, 55, 21, 104, 63, -94, -126, 32, -114, 18, 126, -112, 32, 91, -15, 36, -92, -80, -97, -125, -12, -125, -31, 25, -48, 117, -29, -109, -67, -46, 113, -36, -61, -120, -53, 113, 72, 81, 8, -49, -121, 106, 26, -19, -94, 29, 122, -6, 103, 44, -18, 20, 57, 13, -99, 67, -113, -107, -94, 80, 22, -112, -23, 23, 38, 34, 47, -36, 23, -96, -109, -1, -68, 116, -110, -9, -24, -25, 41, -81, -109, -29, 81, -13, 118, -36, -35, -122, -97, -14, 87, -106, -46, -55, -69, 76, 35, 34, -98, 30, 45, 64, 30, 108, 83, 88, -36, -78, -26, 118, 15, -60, -109, 80, -115, 87, 94, -113, 100, -71, 121, 55, -90, -115, 49, 2, 7, 33, -7, -9, -25, -6, -16, -23, 113, -100, 4, 55, 103, -92, -119, 6, 50, -75, 127, 103, 51, 73, -101, -57, -9, 91, 102, 60, 77, 57, 103, -113, 18, 38, -73, 125, 40, -14, -106, -116, -115, 116, -60, -128, -101, -97, 85, -116, -22, -69, 62, -44, 73, 109, 127, -83, 102, -128, 121, 38, -118, 98, 26, 40, -46, -58, 102, -10, -51, 1, -128, -115, -77, -4, -9, 88, -127, 36, 46, 49, -31, 87, -17, 41, 9, -103, 97, 91, -59, 91, 65, 68, -72, -41, -47, 117, -58, 7, 52, -3, 126, -69, -98, -121, 17, -119, 120, 99, 43, -124, 94, 74, -88, -94, 112, -1, 127, 15, 109, 43, -78, 45, -13, -80, -16, -76, 70, -9, -121, -64, -35, 125, -51, 17, 59, 111, -42, -55, 112, -84, 74, -101, -20, 108, 35, 59, 4, 41, 44, 117, 68, 32, 126, -3, -92, 13, -77, 65, 106, 122, -114, -11, -16, 84, -80, 85, -83, 17, 68, 31, -31, -104, 29, 4, -88, 30, -38, 64, -16, -106, 105, 27, -109, -42, 7, -80, 89, -74, 111, 93, 18, 68, -30, 104, 53, -32, 11, -5, 6, -17, -121, -19, -35, -43, -104, 18, 121, -102, -65, 92, 36, -126, -105, -78, 27, -18, 34, 102, 26, 60, -43, -72, -47, -99, 63, -86, 25, 38, 115, 40, -23, -45, -43, -19, -4, -88, -106, 31, -80, -61, -41, -38, -66, 74, -19, 65, 75, -20, -64, 11, 56, -14, 42, 2, -39, -63, 27, 86, 28, -100, -43, 70, -1, -118, 40, -53, -2, 40, -58, -13, 16, 106, 100, 116, 64, -18, 113, 124, -65, -38, 2, -107, 31, 41, -47, 110, -76, 50, 64, -114, 105, -58, 74, 73, -70, 103, 30, 25, 39, 11, -13, -113, -75, -71, -40, 66, -106, -41, -126, -122, 44, -47, 16, -70, -2, -10, 13, 19, 106, 97, -63, -67, 40, -61, -98, 56, -67, 73, 108, 107, 98, -3, 100, 6, 11, -66, 78, 5, -80, 46, -18, -2, -29, 115, 109, -90, -40, -26, 55, 29, 110, 60, -115, 59, -116, -68, 102, 115, 115, 73, -36, 81, 84, 28, -108, -5, 33, 75, -7, 86, 112, -70, 1, 34, 31, -28, 108, 65, 21, -43, -20, 93, 118, 61, -20, 99, -99, -113, -116, -122, -13, -64, 83, 99, 14, -104, -57, -58, -17, 22, 70, 36, -127, -55, 78, -32, -72, 126, -54, 30, 80, 30, 69, -122, 86, 76, 107, -12, -110, -102, 105, -19, -124, 72, -36, -34, -12, -3, -71, 38, 52, -126, 110, -20, -79, 126, 95, -86, 3, -12, -45, 62, 95, 60, 28, 65, 75, -112, 33, 117, -20, -103, 86, -76, 29, 39, -113, 54, -74, 4, -112, -100, 81, 77, 90, 40, -96, -22, -19, -60, 124, 119, -93, -65, 92, 43, 77, -106, 83, -68, 119, 58, -30, -40, 44, -120, -64, 55, 80, -26, 12, 71, 80, 85, -34, -116, -45, -122, 70, -76, -57, 78, -111, 99, 119, -1, -57, -41, 32, -90, 123, -73, -97, -99, 118, 17, 87, -42, 97, -23, 10, -110, 84, 60, 54, 72, 60, 119, -26, 27, -27, 51, 39, -99, 8, 28, 80, -98, 116, 67, 0, 11, -53, 11, -41, -95, 69, 71, 118, -74, 76, 101, -30, -95, 108, -6, -93, 117, -128, -107, 52, 51, -23, -102, 50, 70, -51, -120, -37, 117, 64, -122, 124, 115, -72, 23, 120, -60, 23, 111, -55, 28, 32, 78, 74, -20, 44, -48, 10, 70, 86, 48, -125, 15, -34, -58, 5, -104, -14, -103, 86, 119, 26, -106, -61, -2, 108, -48, -57, 109, -128, 39, 75, -32, 82, -104, 17, -55, 8, -1, -77, -51, 60, -38, 110, 38, -117, 117, 83, -36, -88, 13, -70, 27, -14, -14, -47, -107, 126, 65, 47, -119, 120, -93, -44, 96, 2, -49, 67, 93, 74, -50, -61, 40, 51, -21, 71, -48, -41, -97, -84, -108, 71, 81, 92, 50, -33, -102, 14, 27, 63, 29, -88, 76, -33, -93, 112, -67, -3, -6, 56, 104, 25, 57, 81, -125, 35, -57, -89, -118, 10, 42, 82, -127, 30, -120, 29, -25, 95, -4, 18, -72, -95, -71, -89, -22, -72, 115, 23, -125, 61, -46, -88, -39, 119, -119, 5, 39, -91, 110, -37, 13, 69, 1, -127, 71, -106, -101, -17, 62, 46, -39, 30, -83, 92, -51, 92, 117, -63, 25, 58, -16, -39, 54, 88, -52, 75, 49, 42, -121, 46, -17, -53, -59, 41, -20, -47, 100, 40, -95, -33, 79, -106, 34, -37, 100, -16, 122, 73, 110, 2, 42, 56, 11, -15, 119, -4, -14, -37, -13, 38, 11, 25, -15, 116, 95, -90, -30, 125, -94, -90, -41, -89, -52, -38, -93, 18, 6, 99, 44, -69, -86, 61, 104, 48, 91, 120, -6, -56, -71, -39, -20, -84, -17, 124, -14, -99, -84, 92, -42, 12, -38, 116, -42, 34, -21, 47, 78, -18, -41, -113, 66, -22, -15, 119, 14, 95, 38, 4, -2, 59, 97, 13, 110, -32, -101, 92, 97, -48, -71, -81, -40, -32, -89, -27, 77, 64, 104, -18, -3, -58, -2, 115, -30, 86, -69, -50, -68, -22, -60, 90, 88, 14, 116, -43, 122, -67, 103, -30, 55, 47, 33, -90, 65, -51, -108, -1, -124, -34, 2, -54, -81, -125, 34, 125, 15, 74, -66, -12, -103, 114, 98, -26, 92, 42, 89, -66, 114, 125, 84, 124, -120, 93, 106, 84, -115, 117, 33, 102, 9, 74, 60, 5, -47, -57, 84, 123, -21, -107, -90, -58, -77, -60, -70, -62, 82, -21, 105, 107, 104, -74, -35, -53, 123, -105, -68, 5, 4, -23, 86, -121, -10, -12, 37, -59, -71, -100, -105, -48, 16, -124, -108, 50, -125, 68, 50, 71, -48, -72, -118, -96, -98, 117, 127, 99, -117, -124, -60, -15, 43, -43, -14, 77, 9, 50, 113, 75, 114, 11, -53, -7, -20, -14, 111, 116, 4, -102, -116, 67, -57, -103, 111, 51, 37, -102, -48, -92, -123, -7, 87, -40, -54, -71, -97, 108, -3, 98, -79, -14, 79, 70, 71, 113, 67, -121, -44, 105, 98, -112, -73, 12, -50, 26, -40, 16, 127, 51, -16, -97, 52, -68, 34, 104, 24, 70, -115, 113, -61, -51, -87, 75, 127, 29, -111, -110, -22, 60, -90, 54, -110, 1, 21, 77, -22, -99, 54, 40, 108, 53, -39, -20, -18, 77, -114, 81, -73, 72, 44, 100, 83, 126, 12, 22, -21, 78, -43, 41, 59, -124, 39, 117, 8, -103, 104, 88, -100, -76, 40, -9, 65, -73, -94, -21, -121, -19, -19, 112, -10, -3, 22, 86, 25, 104, -83, 73, 124, -58, -79, 83, -81, -83, 110, 34, -96, -90, 15, 94, -120, -20, 23, -96, 33, -100, 37, 14, 68, 83, 59, 64, -40, -90, 27, 82, -96, 35, 37, 102, -107, -26, 121, 94, -121, -42, -23, -19, 79, -92, -50, -33, -104, 59, -59, 9, 60, 101, 87, -32, 28, -90, 77, -39, 59, 38, 50, 87, -88, -39, -98, 43, -66, -24, -32, 93, -43, -117, 19, -100, 67, -75, 53, 72, 115, -27, -22, 84, -92, -118, 108, 91, 117, -54, 21, -70, -64, 105, 79, -108, -34, -64, -118, 88, 43, -82, 96, 70, 75, 13, -76, -24, -88, 70, -63, -41, 60, -74, -97, -72, -58, 37, 20, -86, 89, 54, 79, 114, 5, -73, -44, 115, 83, 96, 86, 2, 102, -62, 75, -44, -128, 7, 29, -41, 21, -2, 63, 35, -90, 9, 96, -12, -62, 82, 47, 53, 32, -30, -46, -128, 83, 90, 35, -3, 40, -126, -50, -18, -32, -1, -69, -84, -25, 114, 24, -76, -34, -36, -127, -43, 115, 91, 64, 122, 59, 36, 125, 48, -69, -109, -43, 115, -40, -106, -27, -12, -78, -37, 52, 119, -31, 64, 27, 8, 96, -90, -33, 61, -92, 119, -105, -13, -25, -100, 29, -75, -26, -6, 50, -128, 19, 48, 83, 37, 30, -68, -9, 93, 72, 56, 82, -32, -74, 35, 37, 13, 3, 18, -77, -102, -107, 79, 7, 25, 86, -19, -59, 27, -34, 26, 16, 1, -108, -95, -86, -103, 51, -43, 66, 68, 58, -107, 36, 10, -47, -56, -50, 59, -79, 37, -107, 63, 84, 125, -95, -2, -19, -59, 52, 83, -69, 71, 102, 86, 32, 121, 25, -109, 93, -24, 65, -64, 6, -90, 15, 80, 66, 111, -120, 41, 72, 16, -7, 121, 51, -76, 31, 93, -109, -8, -121, 60, -84, -2, 15, -49, 68, 29, -15, 40, 74, 44, -93, 79, -115, 87, -112, -122, 89, 52, -2, -94, 111, 123, -110, 99, 44, -12, -93, 31, 13, 36, 23, -80, -37, -33, 116, 8, 107, -17, -126, 116, -119, -114, 59, -32, -109, -38, 95, -76, 47, -20, 49, 108, 91, 118, 121, -9, 91, 32, 0, 41, -14, 67, -65, 12, 109, -6, 45, 80, 57, -35, -83, -108, 53, -27, -22, -19, 56, 116, -2, -66, -11, -113, 74, -51, -16, 104, -56, 56, 79, -71, 42, -58, 69, -38, -56, -112, -47, 35, 50, 35, -45, -18, -42, 106, 46, -102, 1, 0, -27, -75, 22, -87, 125, -56, -120, -33, -123, -128, 6, 60, -81, -45, 4, 21, -108, 46, -37, 72, 53, 104, -35, -60, 10, 52, 45, -52, -25, 36, -119, 108, 55, -122, -64, -33, 63, -29, 78, 54, 6, -44, -92, -72, 101, 121, -61, -41, -25, 78, -2, -10, 27, 22, -93, -69, 39, -112, 32, -114, -66, 95, -37, 42, 95, 4, -124, -59, -68, 21, 125, -124, -6, -114, 72, -53, 50, 72, 116, -109, 114, -62, 10, 92, 112, 10, 52, -116, 51, -15, 124, 98, 66, -97, 126, -97, -93, -45, 84, -99, 13, 58, 87, -78, 19, 93, -87, -71, -14, 33, -112, -44, -115, -63, -110, 113, 5, -118, -7, 116, 9, 82, 23, -118, 26, -57, 62, 5, -9, -19, -86, -89, -5, 86, -68, 83, -108, 79, -65, -81, -59, -33, -109, -88, 14, -39, 71, -107, -115, -104, 39, 13, 44, -71, 35, 111, 120, 99, 22, 85, -33, 57, 86, -121, -30, 50, -29, -11, -122, 23, 113, -41, 31, 46, -119, -84, 49, 90, -83, -5, 6, 47, -97, -76, 44, 53, -48, 107, -95, -4, -88, 102, -16, 19, 80, 126, -29, 109, 75, 110, 90, 17, -40, -104, 105, -56, -7, 27, -61, -25, -8, 126, -32, -39, 122, -119, 5, 28, -19, 97, 28, 35, -37, 94, 110, -41, 46, -124, 10, 27, 80, 12, 20, 98, 82, 10, -122, -123, 93, 65, 105, -67, 6, 31, 36, -15, -64, -64, 45, 52, -3, -72, -109, 82, 30, -85, -64, 33, 101, 87, 112, -83, -94, -120, 123, 104, 100, 116, -73, -70, -93, -6, -25, 75, 106, 98, 15, -48, -75, 60, -81, -74, 50, -90, 96, 22, 112, -35, -36, -48, -26, 93, -9, 10, -45, -41, 51, 4, 38, -80, -85, -75, 106, -52, -99, -6, 64, 76, 72, -35, 126, 56, 117, -103, 67, -90, 2, 16, -93, -38, 74, -39, -62, 1, -1, 17, -37, -117, -122, 87, 83, 98, -23, -45, 60, 39, -32, 58, 117, -112, -65, -15, -97, -83, 91, 109, 123, 12, 113, -12, -5, -64, -90, -12, 49, 25, -17, 67, 1, 92, -123, 105, -97, -119, 101, -67, 30, 34, -45, 0, -92, 89, -58, -127, 40, 89, -51, 64, 65, 31, 97, -118, 71, 84, -86, 66, 90, -53, 23, 99, -27, -4, 119, 78, 88, 116, -89, 121, 99, 4, 64, 88, -54, 83, 102, -8, -59, -62, -6, 65, -58, -70, 115, -94, -39, 16, 115, 83, -106, -18, 105, -14, 97, -8, -35, 125, 22, -66, 14, 70, 21, 59, -109, 109, -118, -28, -55, 119, 13, 48, -58, -89, -118, -56, 59, -46, -82, -124, -65, 44, 9, 96, -90, 74, -12, -36, -72, -70, -16, 83, -103, 94, -58, 63, -4, 5, 124, 35, 96, 38, 41, 125, 46, -88, 16, 44, 65, -47, -82, 78, 85, 64, 92, -78, -115, 114, 38, 41, -119, -10, -36, 64, -21, 87, -51, -70, -21, -47, 108, 70, -66, -31, -104, 63, -127, 99, -103, -3, -117, -126, -6, -18, -94, 115, -12, 116, 122, -57, -31, -8, -76, -23, 31, 57, 84, 89, -35, 87, -28, -83, -60, 94, 45, 64, 77, -58, 44, 55, -57, 100, 40, 72, -109, -25, 14, -11, 70, -126, 73, -21, -73, 86, 93, 118, -29, 8, -124, 36, 28, -62, -81, -79, -64, -49, 127, -42, 114, -98, -58, 19, 61, 33, -45, -100, 113, -56, 61, 0, -89, 124, 115, 49, 31, 57, -97, 47, 103, 37, -58, -82, 102, -86, -48, 119, -73, -71, -65, -59, 98, 73, 7, -69, -51, -38, -107, -102, -14, -87, -6, -63, -25, -5, -96, -84, -68, -123, 102, -99, 68, 3, 74, -77, -46, 50, 70, 47, -62, -76, -22, 45, -88, 6, -66, 26, 101, -15, 114, -36, -54, -6, 95, -113, 27, -46, -45, 46, 64, -28, -109, 29, -98, -70, -16, 75, -110, -34, -65, -17, -112, -16, 6, 32, 85, 50, -16, -84, -84, 58, 124, -43, -111, -11, 0, -37, -88, -27, 73, 99, 121, -21, 15, -88, -88, 42, -9, -117, 56, -43, -109, 79, -76, 67, -126, -76, 116, 53, -60, -128, -47, 40, 6, 82, 127, 22, -11, -94, -1, -13, 58, 120, -107, 39, 91, 112, 126, -82, -102, -79, -59, -77, 91, 36, 63, -88, 108, 113, 47, 118, 98, -75, -19, -40, 58, -119, -59, -75, 30, 59, 99, 127, 53, -80, -55, 8, -23, -96, -64, 42, 9, -22, 112, 57, -44, 115, -113, 88, -105, -48, 18, -9, -58, 112, 6, -32, 115, -121, -11, 69, -20, 98, 55, 2, 99, -118, 29, -35, 35, 79, -2, -84, 126, 117, -11, -127, -88, -104, -30, -47, -123, -33, -117, 78, -11, 46, -79, 86, 56, 95, -54, 105, -79, -73, 113, 125, 82, 91, 49, 118, 116, -127, 25, 123, 30, 122, -75, 96, -101, 86, -58, -127, 6, -43, 64, 52, -109, 35, -21, 22, 101, 28, -31, 90, 123, -13, 119, -34, -84, -91, 55, -47, -33, 70, 18, -124, -21, 49, 43, -19, -125, 21, -105, -119, -103, 123, -93, 64, -126, -47, 99, -46, -7, -16, -91, 49, -43, -25, -34, -78, -95, 50, -102, -51, -67, -93, -82, 8, -70, -96, 44, 27, -13, 37, 109, -32, -115, 81, 66, 103, 1, -84, -113, -83, -21, -76, -89, -14, -123, 117, -16, 86, 66, -24, 111, 118, 34, -68, -65, -121, 69, 118, -77, -53, 79, 122, -24, 4, 120, 99, -68, 62, -5, 7, 54, -61, -67, 29, -49, -77, -61, -43, 87, -80, 82, 121, 3, 43, -114, -78, -33, 63, 21, -35, 60, -78, 59, 69, 119, 118, 119, 32, -102, -106, -6, 95, -87, 29, -112, -5, 4, -12, 37, 52, 88, -115, -108, -87, 1, -63, 106, 121, -13, -121, -52, -4, -56, 70, 58, -8, -81, -13, 26, 24, -56, 113, -43, 40, 118, -99, 106, -128, -59, 36, 61, 40, 104, -27, -128, -1, 97, 85, 47, -24, 14, -46, -67, 103, -32, 46, 22, 93, 85, 77, 18, 89, -106, -87, 22, -54, -78, -110, 14, -107, -120, 56, 106, 76, -79, 126, -89, 80, 77, 53, -114, 27, 110, 45, -127, 26, 79, -93, -70, 45, 103, -9, -121, 42, -88, 45, -28, -127, 92, 74, 75, -17, -38, -114, 28, 4, 84, -103, -92, -50, -56, -65, -92, 1, 102, -32, 91, -64, -120, 115, 109, 39, -75, -120, -101, -125, -64, -83, 72, -68, 30, 94, -97, 54, -17, 44, -119, 37, -44, 66, 13, 28, 77, -118, -20, -38, 104, -34, -43, 36, 37, -8, 125, -125, 60, -64, -58, -46, -50, 116, -51, 13, -83, 123, -96, 41, -7, 120, -113, -63, 88, -126, -30, 19, -51, 17, -107, 5, 15, 85, 32, -49, -102, -108, 99, -67, -116, 50, -105, 30, 93, 52, 17, -74, 58, -28, -85, -75, 71, -57, -59, -106, -116, 111, 3, 106, -74, -27, 41, 102, -43, 7, 59, 79, -111, -50, 92, 27, -104, -69, -92, 94, 114, -110, -43, 9, 98, 124, 21, 83, 109, 32, -14, 94, -97, -85, -2, 56, -53, -26, 108, 126, -104, -95, 28, 33, -80, -34, 98, 38, 71, 75, -71, 30, 59, 126, 43, -111, 120, 119, -47, 38, 76, -95, -64, 39, -104, -71, 12, -116, -4, 74, -53, -74, 91, -32, 30, -82, -88, -30, -93, -19, 41, -53, 20, -102, 109, -115, -28, -16, -77, -66, 0, 20, 94, -98, 49, -5, -62, -36, 120, -7, -41, 126, -116, 87, -100, -38, 2, 67, 10, 36, 46, 86, -18, -104, -90, -29, -17, -87, -118, -114, -69, 48, 75, -101, -33, -115, -37, -87, 57, 70, 86, -77, -3, -108, 11, 86, -21, 54, 3, -91, -63, 125, 49, -109, 1, 62, -112, -57, 18, 19, 121, -99, 19, 112, 81, -10, -22, 91, 64, -119, 102, 109, -71, -4, 7, 126, -82, 59, -17, -85, -122, 41, 113, 118, 4, 72, 11, -4, 96, 122, -80, 33, -43, -120, 35, -37, 49, 27, 12, -80, 46, 3, 5, -82, 126, 55, 124, 98, 120, -94, -77, 64, -28, -99, -76, -125, -118, 101, 12, -49, -84, -77, -25, -118, 98, -73, 48, 71, -23, -98, -19, -41, 43, -98, 92, 93, 25, -102, -110, 0, -88, 108, 38, -46, 37, -36, -38, 8, 22, 78, -27, -16, -30, 11, -55, -97, 18, 96, 43, -112, 20, -121, -125, -53, -91, -124, -35, 115, -68, 81, 27, -123, 7, -15, -105, 104, -116, 89, -54, -51, -23, 118, 81, -56, 50, 23, 126, 41, 26, 51, 1, 59, -36, 81, 59, -40, 20, 117, -117, 112, 66, -10, 80, 113, 49, 58, -113, -41, -92, 43, 118, -46, 79, 0, 114, 20, -41, -108, 68, -112, -8, 7, 7, -62, -80, 94, -81, 111, -55, -91, 30, 12, -92, -69, -109, 79, 37, -122, 2, 94, 105, -78, -34, 74, 17, -99, 76, -60, 63, 36, -84, -96, -126, -70, -77, -30, -14, -40, 117, -74, 35, 63, 87, -46, 122, -56, -106, 55, 60, -4, -49, -11, 59, 124, 95, -112, -32, -34, 78, -97, 122, -56, -32, 8, 35, -87, 12, 36, 54, -2, 61, 30, -32, -58, 2, 120, -128, -29, 38, -66, -127, 7, -79, -22, 30, 67, 28, -104, -103, 6, 110, 116, -111, -8, -20, -117, -29, 84, -85, -66, 43, 107, -121, 112, 125, -75, 57, -12, -10, 0, -38, -117, 27, 117, -45, -48, -116, -1, -119, 122, -56, 50, -110, -108, -127, 60, -120, 51, -46, -120, -82, -88, 93, -104, 43, 118, -67, 48, 102, 42, 109, 16, 1, 75, 88, 26, 11, 0, 4, 28, 116, -122, 104, 9, 80, 59, 24, 100, 126, 23, -31, 16, -6, 53, -66, -91, -122, -112, 37, -97, 27, -74, 58, 48, 66, 64, -19, -11, 31, -12, -44, -64, -121, 38, 126, 30, -100, -110, 78, -107, -96, -60, -86, -39, -74, 57, 97, -122, -94, -119, 66, -61, 30, -93, -70, -117, -57, -113, 30, -29, -126, 123, -84, -90, -39, 58, -33, 30, -83, 14, -106, 30, 125, 14, 127, -125, -114, -110, 88, 19, -74, -102, -95, -35, -101, -40, -107, 53, 114, 29, 10, 22, 106, -67, 121, -102, -68, -12, 10, 41, -72, 73, -89, -9, 36, 96, 119, -35, 117, -25, 105, -66, -23, 26, 20, -124, 70, -92, 1, -13, -67, 124, 108, -18, -103, -79, 35, -11, -36, 26, -101, 120, -19, 123, -70, 3, 49, -3, 66, -73, -104, 92, 79, -47, 70, 111, 40, 32, 124, -6, 9, -60, -123, 36, -54, -80, 99, 21, 36, -103, -60, -123, -117, -60, 113, -67, -92, -13, 22, 84, 11, -111, 107, -7, -125, 32, 84, -35, -40, 32, 100, -59, 57, 19, -25, 23, -111, 88, 50, 1, 95, -90, 123, 8, 101, -59, 36, -13, -105, 16, 25, -43, 54, -88, -92, -61, 60, -23, 38, -52, -43, 61, 25, -86, 98, -86, 31, -58, 15, 27, -61, -115, 11, 121, 36, 104, 88, -9, 74, -35, 106, -119, 1, 98, 14, 32, 112, 93, 24, -65, -10, -49, 71, -72, 122, -86, 71, -125, -75, 97, 124, 31, 124, -52, -68, 67, -93, -5, -36, 51, 41, 122, 3, -95, -112, -84, -101, -80, -18, -127, -7, -32, 127, 74, -75, -103, -101, 124, -74, -70, 93, 80, 115, 60, -41, 10, -85, -20, 37, -23, -95, 89, 79, 32, 19, 23, 20, 55, -107, 107, -128, -9, 75, -128, -118, 26, -39, -60, 101, 27, 124, 83, 29, 111, -124, 10, 75, 100, -94, -11, 104, 16, 57, -3, 49, -119, -96, -69, 93, 65, 55, 86, 71, -47, -90, -37, -120, 90, 107, -53, 0, 17, 81, 111, 57, -120, 0, 91, -16, -20, 64, -90, -105, -61, 93, 120, -56, 64, 47, -70, -34, 53, 8, -46, 105, -99, 19, -36, 80, 12, -90, -39, -49, -53, 20, 10, -1, 81, 64, 58, 20, 42, 39, 30, -127, -20, -37, -117, -3, 66, 5, -126, -126, 96, -127, 84, -125, -24, -11, 81, 107, -59, 83, -67, -40, -2, -89, 126, 71, -73, 45, 28, 109, 14, 64, 72, 53, 31, -56, -76, 12, 84, 77, 30, -95, 11, 78, 102, 32, 74, 127, 37, 97, -8, -27, -26, 64, 96, 110, -1, -62, -29, 110, 28, 98, -41, 27, -43, 55, -53, -81, 72, -125, 26, -13, -103, 2, -110, -120, 10, 1, -70, -31, -35, 36, -12, 124, -50, -38, 1, -82, 120, 74, 50, 5, -71, 56, -96, -103, -75, -51, -74, 19, -14, 110, 68, -56, -43, -98, -125, 91, 12, 105, -66, -87, 45, -99, -21, -31, -53, 108, -45, -124, 107, 16, -110, 60, -89, -118, -93, 64, 98, 14, 34, -74, -29, 66, 7, -112, 49, 125, 112, -11, 48, 82, -31, -108, -121, 21, -101, -17, -55, 105, -72, 32, -12, 104, 83, 19, -13, -52, 105, -87, 68, -34, -5, -1, 4, 64, -106, -43, -40, -95, -68, -6, 14, 61, 48, -88, -66, -124, -17, -38, 111, -40, -89, 105, 17, 101, -128, -81, 13, -46, -49, 49, -23, 18, 107, -82, -75, 69, 122, 79, -101, 52, -125, -70, 80, -100, -18, 79, 0, 108, -110, -115, -47, -34, -31, -80, -66, 89, 83, 42, 36, -4, 116, 33, -80, 111, 23, -35, -21, 13, 51, 55, -5, 60, 109, 12, -116, 111, 121, -16, 73, 100, -121, 42, -127, 115, 21, 3, -89, -94, -99, -112, 4, 28, 37, -56, -25, 30, 93, -117, -108, 25, 88, 83, 68, 108, 49, -126, 26, -16, 38, 80, -19, -119, -77, -60, -119, 20, -12, 4, -112, -117, 30, 107, 68, -73, 86, 113, -75, 5, -109, -45, -56, -97, -27, 41, 8, -123, 47, -33, -17, 58, 1, -105, 66, -89, -124, 27, 56, 7, 70, 104, -98, 104, -103, 64, 111, -117, -2, 97, -19, 63, 77, -37, -125, 65, -83, 89, 97, 52, 55, 78, 120, 74, 124, 12, 50, -107, 95, -114, -38, -99, -76, 48, 34, -71, 126, -13, -75, -57, -50, -112, -111, 37, 97, -44, -80, 108, 1, -67, -83, 66, 76, 59, 54, -24, -103, -57, 40, -94, -50, 93, 64, -75, -73, -79, -32, -72, -105, -45, 32, 49, 77, 93, -31, -122, 81, -123, -15, 16, -110, -93, 47, -59, 61, -69, -51, -84, 28, 33, 102, 110, -128, -73, 24, -53, 59, 1, 34, 44, 77, 35, -22, 34, -124, 126, 10, -36, -61, 101, -52, 11, 114, 5, -113, 24, -35, 33, 53, 123, 81, 43, -124, -105, -54, -14, 57, 58, -4, 122, 110, 71, -38, -26, -48, -13, -12, 6, 46, 17, 85, -80, 4, -55, 17, 115, 52, 41, 122, 115, 47, -104, 46, -114, -97, 102, -55, 28, -37, -19, 45, -87, -119, 76, -100, 93, 35, 90, 90, 4, -85, -6, -79, -51, 49, -39, -73, 6, -113, 64, 124, 63, 41, -45, 99, -45, -88, 56, -124, 62, 18, -88, 109, 36, -69, 91, 124, -77, 103, 17, -30, -48, -17, 40, 63, 9, -53, 101, -106, -119, -10, -104, 106, -82, 124, -93, -30, 3, -94, -93, -34, -75, 126, 73, -59, 56, 36, 54, -9, 65, -125, 15, -32, 116, 2, 123, 125, -86, 29, -104, -69, 46, -39, -96, -28, -115, -27, 1, -125, -42, 67, 38, -121, 38, -110, 18, -116, 126, 105, 62, -62, -126, 94, 62, 110, -45, -113, 81, -59, -118, 83, 100, -37, 36, -12, -112, -68, 36, -60, 114, 3, 15, -113, -108, 64, -40, 39, -73, 43, -126, -108, 98, 25, 18, 32, -45, 78, 126, 19, -109, 112, 107, 16, -91, -21, -78, 54, -98, -89, 111, 61, -96, -34, 14, -68, -3, -58, 100, -34, -10, -25, 81, 67, 28, 91, -120, 21, 107, -25, 63, -74, -61, 26, -98, -95, 121, 58, 73, -40, 110, 77, -24, 102, 89, 123, -29, 109, 95, 24, -21, -38, 59, -44, -12, 110, -64, -86, 5, 28, 56, -90, -76, -23, 68, -36, 59, -87, 40, 94, 95, 84, 88, -39, 63, -59, -32, 8, -110, -6, 22, -108, 47, -112, 8, 91, 17, 27, -68, 115, 25, -94, 31, 51, -86, 17, -14, -84, 36, 37, -7, -103, 119, 123, -26, 77, 2, 86, -98, -51, 76, -42, 121, 125, 29, -12, -10, -58, 88, 0, 86, 39, -99, -90, 41, -107, -50, -82, -24, 105, -90, 46, -115, 94, 79, 28, 72, 89, -29, -118, 13, 74, -88, -39, -67, -16, -53, 54, -66, 101, -35, 53, -43, -13, -17, -57, 37, 102, -51, -64, -87, -59, -49, 100, 54, 80, -43, 55, -52, -27, -25, -16, 73, -65, 26, -66, 19, -12, -20, -71, 24, -106, 66, -94, 51, 50, 70, 122, 121, -32, 73, -88, -59, -108, -79, 61, 23, 55, 75, 77, 59, -5, 69, 56, -17, -21, -74, 120, -99, -81, -34, 30, 46, -59, -79, -23, 118, -53, -36, -115, 122, -63, -71, -104, -91, 10, 72, -120, -19, -94, -99, -44, -64, 27, -49, -49, -1, 106, 84, 30, 5, 52, -14, 7, 2, 7, -19, 65, 94, 35, -28, -118, -98, -25, -39, -58, -30, -84, 126, 83, 59, -12, -43, -109, -4, 38, 92, 34, 24, 30, -104, 121, -89, -36, -5, 119, -96, -121, -121, 71, -30, 25, -13, 57, -54, 99, 12, -39, 62, 61, -94, 14, -125, 103, -123, -83, 59, 0, -110, 29, -98, -76, 42, -60, 37, 124, -97, 113, 38, 39, 127, 78, 17, 53, 19, 28, 106, -76, 72, -53, 8, -123, -107, -2, -15, 49, -68, 58, -31, 77, -45, 7, 48, 86, 38, 69, -23, -18, -46, -72, -103, 20, -94, -124, -114, 55, 0, 85, -49, -54, -66, 34, -114, -52, 28, -63, 103, -112, -35, -23, -14, 13, 123, -115, 0, 80, 85, 29, -1, 51, 11, 121, 84, 127, 36, -59, -51, 15, 61, -63, -48, 106, 55, -11, 14, 8, -109, 110, -15, -50, 73, 120, -92, -115, 29, -39, -111, -32, -13, -19, 51, 114, 47, 13, 109, 85, 125, -4, -61, 13, -109, 73, -25, 109, 70, -90, 55, -26, -124, -27, -24, -17, -112, 89, -97, 36, 32, -62, 4, 49, -1, -55, -88, 24, -48, 122, -128, -6, 95, 100, -87, 62, -87, -70, 12, 88, -103, 111, -75, -27, -88, 20, -12, 76, 115, -18, -54, -22, -28, 98, 90, -91, 40, -39, -29, -94, 61, -15, -55, -7, 101, -81, 53, -1, 110, -38, -125, 109, -7, 94, 102, -88, 16, -31, 118, -104, 69, -115, -2, -77, -39, 8, 5, 22, -1, 73, 107, 32, 91, 84, 0, -3, 109, -85, -69, 54, -120, -68, 110, 59, -43, -61, 75, 120, -84, -85, 3, -55, 100, 3, -84, 35, 114, 22, 71, 109, -74, -101, -26, 56, -113, 115, -121, -63, 70, -127, 28, 67, 94, -13, -30, -36, -109, 29, 32, -80, 124, 96, 48, -77, -13, 1, -63, 127, 114, 37, -1, 38, -87, -92, -28, -30, 104, 16, 0, -13, -107, 33, -9, -26, 13, 4, -10, 44, -94, 49, -117, -35, -29, 126, -36, 106, 32, -32, 10, 5, 68, -2, 3, 13, 110, -99, 18, 116, -126, -86, 44, 104, 28, 85, -86, -99, -127, 121, -105, -116, 15, -58, -66, -51, -109, -88, -90, -20, -33, -68, 32, -16, -28, 89, -90, -101, 80, -21, 94, -41, 86, -6, -4, 73, 18, -22, 35, 56, 118, -16, -128, -71, 37, 84, 79, 106, 125, -51, 101, -92, 6, -84, 92, -26, 18, -7, -9, -40, -91, 46, -60, 4, -127, -122, 110, -32, 28, -28, -120, -104, -80, 60, -120, -50, 9, 13, -25, 40, -91, 25, 29, 82, 92, 119, 14, 112, 109, 84, 50, 30, 59, 86, -112, -119, -90, 120, -2, -106, 122, -4, -85, -47, 38, -68, -20, 114, -121, 112, -38, 122, -95, -117, 107, 111, 127, -36, -112, 34, 22, -61, 76, 1, 28, 87, 110, -56, -10, -57, -66, -75, 105, -122, -84, -28, -107, 94, -124, -5, 0, 26, 68, 127, -92, 3, -37, 40, 46, 31, 52, 29, 56, -16, -99, -29, -44, 17, -40, -14, -69, 46, -80, -29, 25, 23, 114, 105, 70, 81, 71, 103, -83, 20, -65, -13, 50, 26, -61, -79, 90, 112, -44, -23, 107, -42, -21, 43, -104, -21, 30, -10, 72, 116, 17, -99, -76, -48, 0, -50, 90, 42, 83, 21, 127, 58, 65, 37, 46, -81, 121, 17, 40, 47, 21, -103, 27, 111, -118, -16, -64, -92, 40, 41, -69, -43, -70, -42, 9, 30, 54, 124, 85, -29, -5, 120, 5, 24, -73, 45, -109, -7, -108, 113, -96, -52, -1, -106, 82, 102, -34, 124, 118, 118, -50, 86, 115, -127, -19, 75, -70, 107, 78, -26, 77, -20, 39, 123, -122, -62, 42, -15, 58, -22, 90, -7, 71, 95, -13, 86, -59, -116, 69, -31, -9, -28, -45, 76, -81, -21, -90, -124, 4, 32, -120, 2, -9, -112, 82, 88, 32, -52, -106, -66, -117, -85, 91, 74, -21, 35, -109, 14, 86, -26, 119, -3, 92, 121, -26, -106, -25, 14, -54, -61, 28, -26, -102, -18, 45, -18, 66, 35, -93, -29, 16, 37, -97, 110, 109, -20, -84, -118, -104, 3, -116, 76, 64, 88, -55, -2, 12, -109, 127, -14, -78, -90, 127, 93, -61, 74, -99, 35, -107, -53, 14, -114, 118, 45, -24, -27, 13, -88, 104, 26, -114, 96, -9, -44, -62, -18, 46, -13, 57, -80, -22, -99, -8, -80, 47, 80, -122, 19, 19, -121, -54, 120, 118, -115, 89, 82, 100, 4, -112, -58, -126, 108, -9, -112, -81, 39, 27, 78, 38, 83, -101, 124, -19, -90, 112, 67, -45, -21, -91, -63, -22, -96, -47, -71, 20, -125, 69, -112, 27, 60, 124, 28, 25, 7, -127, -18, 114, -75, 54, -26, 73, 127, 7, -75, -7, -44, 75, 95, -76, 44, -120, 120, 56, -72, 44, 27, -98, -92, 127, -111, 109, -30, 24, 91, -98, 111, 33, 61, 107, -45, -45, -46, 45, -93, 11, -47, -1, -91, 107, -18, -117, -92, -108, 89, -125, -114, -1, -50, 56, 19, -51, -26, -73, 16, 2, 95, 107, -36, -26, 57, 45, -122, 20, 58, -94, -96, 27, 113, 65, 72, 72, 59, 91, 5, -105, 43, 118, 54, 97, 8, 30, -88, -106, -113, 46, -97, 87, -97, -97, 119, -28, -81, 7, 72, -103, 63, -112, -27, 49, 81, 37, -43, 8, 73, -78, -22, -111, 63, -105, -37, 77, -115, -34, -41, 72, -125, -76, -120, -26, -73, -77, 115, -16, -97, -33, 39, 87, -11, -112, -2, -119, -64, 126, 65, -92, 101, 58, 77, 127, 34, 51, -114, -5, 24, 43, -36, -26, -71, 32, -63, -73, 7, 44, -87, -63, 103, 20, -19, -24, -41, 7, 119, 1, -54, -51, 47, 106, -119, -73, -19, 7, -120, -54, 115, -62, 114, -98, 2, 35, -17, -113, 57, -68, -15, 100, -26, 87, -10, -64, 85, -74, -41, 3, 44, 24, -63, -18, 24, -51, -116, -4, -78, 27, 108, -74, -117, -38, 77, -110, 82, -37, 112, -17, -33, 71, -8, 96, 101, -67, 57, 16, 58, -38, 111, 97, 81, 28, -27, -42, 105, -24, 7, -127, 49, 29, -109, 11, -16, 121, 15, 17, 111, 123, -29, -114, 94, 111, -49, -69, 56, 50, 112, 118, 78, -43, 10, 35, 101, 72, 118, 108, -31, 63, -48, -69, -69, 62, -69, 6, 108, 114, -128, 100, -18, -97, 19, -89, -7, 19, 84, 11, -25, -15, 79, -29, 79, -116, -47, 55, 66, -82, -58, 93, -81, 35, -69, 68, -96, -6, -68, 108, 22, -41, 89, 53, -32, 92, 83, -42, -85, 87, -28, 90, -22, -114, -14, -72, -35, 44, 15, -25, -20, -1, 101, -67, -79, -90, -1, 51, -75, 5, -28, -62, 25, -13, -27, 67, -84, -23, -62, -22, -114, 28, 11, -66, 69, -50, 65, 97, 109, -118, 57, -91, -12, 74, 115, 103, -58, 74, 78, 60, 82, -45, 91, 95, 124, 4, -59, -23, -58, 68, 98, -85, -113, 86, -119, 99, 10, -93, 21, 25, -77, 111, -93, -70, 79, -39, -11, 92, 79, -22, 121, 12, 116, -24, 39, -14, 114, -66, -69, 78, 83, 51, 15, -27, -68, 23, -12, -116, -3, 90, -1, 56, 1, 92, 82, -16, 71, -64, -125, -12, 116, 73, -104, 105, -60, -128, 84, -80, 90, 29, 98, -120, -84, 90, -77, 117, 53, -99, 17, 18, -124, -82, 39, -107, -122, 69, 101, -122, -46, -10, -75, 122, -103, 49, 99, 0, 49, 18, -108, -47, -28, -70, 62, -44, 121, 127, 29, -48, -114, -98, -7, 88, -5, 101, 97, -23, -47, 114, 87, -64, 91, 66, -88, -69, -47, 14, 25, -73, 121, 66, -40, -50, 95, -83, -122, 40, -46, 66, 95, -60, -85, 64, 38, -28, -49, -120, 57, -92, 117, -43, 82, -73, -59, 52, 41, 34, -23, -120, 94, 31, -105, 90, 40, -34, -30, 104, -57, 27, 88, 21, 4, 118, -106, -5, -31, -92, 10, -73, 7, 99, 84, -78, -97, 72, -54, 61, 48, 12, 41, 55, 126, -21, -127, 27, 12, 82, -30, 57, -37, -104, -112, 92, 29, -100, -81, -10, 103, -22, -83, 102, 90, -70, -85, -112, 86, 97, 113, 84, 119, -116, -10, -39, -120, 8, -28, -14, -107, 54, -38, 23, 69, -2, 9, -115, 87, -9, 2, 29, -98, 54, 98, 112, 97, -42, -119, 48, -41, 126, -48, 80, 122, 78, -89, 10, -54, 45, 9, 16, 90, 27, -127, -33, 17, -62, 29, -50, 68, 13, 31, 55, -47, -4, -74, -28, -2, 119, -50, -110, -13, 110, 58, 11, 90, -23, 89, -31, -19, -127, -106, -103, -66, 31, -46, -100, -22, 117, -71, 8, -28, 126, 113, -78, 92, -23, 86, 105, 31, 44, 93, -18, -31, -104, -39, -74, 27, 126, 49, -84, -97, -27, -82, 26, 12, 57, 95, 2, 70, -67, -38, 114, -117, -114, -118, 87, 105, 63, -21, -124, -29, -38, -115, 97, -69, 39, -114, 101, 9, -60, -82, -50, 29, 125, 18, -70, 9, -100, 25, 28, 47, 25, -70, -18, 1, -70, -41, -37, 105, -39, -10, -69, -89, 96, 104, 10, -67, -90, -79, 50, -98, -94, -28, -80, 30, 117, -24, 86, 111, -121, -78, 18, 96, 40, -62, -14, 91, -35, -46, 109, -37, -74, 116, -17, 68, 115, -67, -118, -76, -80, 119, -128, -97, 104, -25, -32, 79, -99, -121, 46, -123, -53, 117, 84, -30, -82, 95, 116, 89, 94, 93, -109, -112, -115, -19, 114, -94, 104, 0, 79, 37, 64, -26, -106, 25, 62, 58, 104, 20, -11, -55, -12, 116, -24, -88, -14, 123, -124, 125, -11, -89, -57, -124, 70, -63, -125, 47, 76, -62, 127, 109, -92, 11, -81, -77, 25, 90, -58, -29, 60, -126, 41, -74, 96, 121, -64, 110, 127, 30, 25, -11, 78, 95, 32, 118, -26, -88, -15, -28, -66, 122, -66, 10, 100, -64, 45, 93, 5, -71, -95, -114, 122, -24, 61, -82, 72, -39, -26, 71, -41, 102, 31, 11, -102, 97, -4, 125, -93, 116, -46, -33, -103, 105, -96, -121, 25, 49, 90, 58, -1, -74, 57, 30, 18, 32, -120, -103, -122, 114, 27, -104, 23, 44, -88, -92, -73, 127, -17, 107, 11, 32, 90, 89, 47, -50, -92, 74, 66, 69, 76, 124, -108, -74, 93, -24, 46, 63, -55, -43, -83, 114, -98, -80, 13, -41, -51, -13, -127, 112, -57, -99, 107, 102, -2, 28, 42, 119, -54, 93, -109, 11, -58, 84, -38, -41, 2, -102, 76, 115, -93, 38, -13, -77, -7, -23, 38, 91, 91, -107, -96, -14, -41, -48, 8, 73, 91, -9, 21, -91, -96, 82, 99, 26, 100, 24, 25, -50, -89, -84, -19, 19, -38, 63, -20, -19, 121, -128, 24, -104, -45, 95, -68, -99, -48, -106, 14, -28, 77, -106, -105, 99, -66, -32, 32, -50, -16, 27, 54, 99, 123, 73, -41, -124, 24, 90, -26, -58, 86, 73, -88, 58, -34, 4, -7, -102, 69, 20, 80, -17, 96, 75, 42, -4, -36, 47, -87, 8, 17, 118, 44, 46, -19, -111, 39, -84, 63, 15, 83, -119, 89, 70, -77, -39, -58, -47, 70, -26, -47, -121, -45, -46, -52, -90, -34, 95, -110, 81, -75, -82, 89, -126, 93, 28, -2, -101, -55, -90, 65, -119, -95, -20, 99, -50, -93, 72, -4, -68, 4, -17, 116, -40, -60, 36, 88, -103, 118, -20, -27, -3, 62, -113, 27, -83, -3, -113, -8, -108, -83, -58, 21, 38, 52, 122, 12, -101, 121, 47, 112, 52, -117, -33, -58, -15, 102, 79, 12, 96, -25, 110, -80, 126, 34, -46, -34, -6, 33, 91, 42, 63, -121, -18, -116, -72, -80, -126, 34, 3, -111, 79, -50, -81, 32, -128, -62, 43, 72, -7, -128, -32, -99, 2, 98, -65, -89, 71, 114, 11, 60, 65, -40, -51, 47, 56, -81, 122, -37, -38, -37, 34, 123, 53, 39, -23, 16, -119, -63, -13, -17, -37, -75, -4, -51, 85, -19, -115, 82, 59, -116, 83, -13, 39, -76, -63, 82, -123, -74, 64, 110, -16, 118, 31, -21, 107, 124, 6, -46, 58, 14, -66, 48, -30, -26, 93, -59, 114, 70, 96, 114, -46, -28, -17, 31, 57, -118, -124, 19, -7, -51, 27, 67, -105, -53, -46, -92, -21, 127, 120, -18, -37, -35, 98, -34, -34, -96, -36, 51, 108, 60, -110, -11, -34, 51, 20, -71, -106, 30, 24, -121, 62, 52, 5, 9, -26, 44, -71, 24, 78, 28, -122, 61, -1, -55, -66, 15, 112, 115, -78, -6, 79, -24, 29, -62, -80, 106, -20, 88, 54, -126, -109, 35, -123, -60, 126, -112, 56, 33, -41, 3, -106, 0, -120, 29, 107, 31, 54, -26, 17, 48, 87, 73, 27, -47, -16, -3, -59, 85, 32, 45, -117, -86, 68, 69, 61, 66, 32, 125, -114, 84, 80, 74, 38, -18, -64, -94, 15, 28, -62, 69, 65, -36, 34, -123, 66, 43, 80, -123, 56, 73, -92, -98, -91, 24, 62, -51, -48, 111, 39, 88, -82, -6, -120, -39, -116, -76, -122, 49, 12, 19, -62, 14, -5, -123, 103, -38, 67, 12, 63, 41, -1, 104, -71, 3, 102, -55, -88, 70, -89, -55, 16, -115, -104, -52, -96, 14, -115, -11, -7, -17, 115, 80, -38, 112, 17, -22, -62, 99, 53, 52, 115, -76, 42, -83, -90, -69, -90, -97, -12, 86, -52, -21, -24, -80, -109, 10, 19, 109, 33, -11, 121, 123, -22, 105, 81, -20, 11, 112, -12, 49, 44, -43, 8, 23, 127, 64, -29, 75, 111, -48, 44, 126, 111, -31, -56, -119, -73, 50, -34, -50, 125, 119, -39, -5, -89, 32, 113, -90, 15, -54, -25, 99, 19, 47, -92, 102, -121, 82, -115, 4, 39, -65, 110, -116, 9, -110, -124, -94, 100, 74, -37, 118, 16, 11, 91, 55, 48, -109, -76, -95, 56, -41, -67, 127, -87, -105, 65, -93, -55, -25, -63, 11, 58, 4, 12, -8, -6, 89, 86, 23, 82, 116, -107, 104, -75, 63, 67, -93, 17, 124, -96, -89, 88, -4, -32, 56, -13, 61, 8, 94, 52, 102, -81, -24, 51, 30, -76, -37, -109, 81, -76, -86, 32, 27, 73, -97, -7, 42, -41, -11, 26, -66, -115, 119, -93, 15, -54, 74, 35, -50, 37, 116, -125, -57, 12, 72, 87, 22, 86, -96, 8, 113, -34, -5, -101, 99, -23, -106, -99, -57, 32, -85, -26, 79, 83, 17, -116, 56, -30, -86, -91, 14, -23, 44, -69, 63, -34, -37, -58, 68, 127, -54, 86, 117, 12, -6, 103, 115, -126, -21, -67, -37, 36, -121, 125, 20, 45, 63, -106, 112, -32, 101, 48, -103, 117, -111, 96, 125, -53, 76, 15, -62, -97, 101, 60, 126, -65, 49, -26, -13, -49, 112, -69, -20, -76, -111, 0, 109, -15, -108, 15, -77, 67, 64, 33, 70, 125, -62, 60, -83, -126, -60, 45, -9, -124, -30, -10, 105, -92, 68, 123, -113, -42, 49, -61, 11, -43, 106, -52, 65, -96, 87, -46, 43, -97, 47, 84, -100, -115, -94, 10, -76, -105, -4, -55, -110, 96, -69, -20, 127, 90, -42, 22, 125, -102, -4, -48, -35, 1, 116, -41, 101, 77, 123, 126, -64, 40, 103, -93, -50, -57, 16, 1, -123, 60, -51, 126, -97, 4, 85, -42, -109, -21, 57, -24, -59, 62, 71, -78, 18, 19, 68, 127, 40, 12, 68, 30, 39, -114, 27, -74, 3, 36, 88, -79, 98, 111, 37, 103, 97, -127, 49, 120, 56, 99, -122, -34, 72, 54, -57, 95, 92, 116, 36, -24, 58, -68, 120, 81, -34, -86, 2, -25, 104, 49, -46, 40, -57, 47, -72, -89, -110, 80, -46, 92, 98, 107, -94, 37, 58, -112, -19, -119, -83, -99, -57, -5, 115, -1, 59, 34, -75, 105, -69, 120, -128, -19, 27, 20, 45, 66, -105, -116, -98, 113, -20, -61, -115, 123, -64, 123, -4, -3, 127, -70, 49, 75, -109, 26, -95, 34, 127, -11, -104, 74, 4, 44, -91, 83, -86, -99, 33, 36, 66, -12, 109, 31, 98, 97, 50, 33, -120, 110, 73, -51, 72, -17, -79, 48, 71, -37, -94, -65, 114, 102, 70, -74, -35, -90, 108, 125, -24, -97, 105, -45, 86, -12, -62, -57, 90, -120, 37, 48, -126, -47, 92, 119, 73, -62, 53, 52, -120, -73, 93, 16, -78, -70, 98, 48, -68, 92, -45, -23, 54, -3, -46, -10, 25, -42, -85, 120, -125, 24, -14, -108, -111, 7, -99, 48, 50, 23, -44, 106, 19, 61, -120, -49, -35, -82, 61, -3, 19, -25, -95, 28, -45, 62, 97, 4, 61, -104, 124, -125, 12, 82, -122, -75, -1, -60, 40, -55, -15, 20, -88, -126, 51, -115, 52, -68, 94, -114, 112, 4, 51, -4, -14, 37, 4, 124, -41, 72, -110, 85, -91, 21, 56, -33, 76, -40, -4, 124, 11, -3, -51, 28, -95, -114, 108, -123, -71, 101, 16, 87, -74, -53, -21, 52, -99, -119, 61, 9, 30, 85, 21, -94, -51, -2, -90, 12, 66, -52, 57, 38, -44, -60, -25, 68, -24, -64, 95, -119, -60, 55, 6, -125, -125, -105, -70, 103, -36, -85, -9, 73, 95, 82, -52, 86, -49, 97, -103, 38, -120, -61, -62, 15, 77, -66, 39, 119, -17, -108, 106, -71, 108, 57, 118, -71, 53, -26, 112, 6, -123, -1, 60, 121, -125, -59, -126, 95, -89, 86, 13, 46, -92, 21, -54, -59, 124, -37, -37, -43, -34, 14, -110, -56, 3, -10, -51, 104, -104, 40, -12, 1, -5, -26, -122, -11, -99, -4, -33, 75, 95, 28, -75, 36, -67, 109, -111, 40, -40, -30, -9, 12, -94, -45, -117, -61, 89, 46, 86, -118, 126, -8, 8, 121, -121, 89, -117, 53, 16, -93, -120, 29, 41, -69, 87, -76, -63, -5, -128, 105, -43, 47, -103, 36, -63, 106, -106, -107, 42, 68, -35, 15, 24, 7, -90, 6, 12, -111, 17, -102, 28, 33, -50, -36, -97, 61, -127, -76, -121, 93, -77, -110, -55, 117, -80, 69, 109, 76, 5, 30, -102, -103, -64, -87, -95, 119, -87, -3, 45, 8, 66, 29, -29, -110, -57, 120, 69, -60, -5, 115, 116, 86, 5, -92, 86, 105, 119, -58, 17, 35, 113, -14, -28, -19, 24, 58, -21, 13, 34, -100, -100, -56, -101, -83, 91, -96, -114, -10, -104, -35, 64, -67, -121, -33, 25, -50, -117, -23, 49, 10, 76, -78, -37, -10, -96, -110, -51, -10, -67, -55, -127, -73, -84, 66, 74, -75, -86, 94, 16, 69, -86, 5, -47, -11, -43, -48, 82, -51, 110, -117, 90, 113, -70, 73, 69, 88, 99, 93, 119, 110, 3, -80, 88, 117, -93, 105, 78, -45, 62, -80, 30, 117, 26, 99, -42, -103, -82, -83, 60, -23, 59, -29, 36, -64, -31, -44, 92, -34, 87, -48, -56, 102, -113, -6, 89, -28, -15, -90, -121, 51, -28, 84, -21, 61, -104, 57, 47, 45, 55, -22, -42, 24, 99, 40, 51, -45, 119, -26, 3, -26, -18, 42, 75, 98, 59, 94, -113, 79, 74, 4, 116, -82, -50, -15, 59, 56, -26, 114, -38, 14, 72, 44, -109, -85, 27, -12, 93, -127, 87, 6, 75, 37, -94, -26, -2, -103, 118, -106, -83, 14, -100, 12, -52, -55, -46, -62, -110, -27, -94, -14, 5, 83, -88, -33, 22, 106, -15, 54, -91, 47, -77, -120, 27, 3, 46, 86, -86, -125, 59, -117, -58, 65, -46, -31, 23, -4, -61, -41, 116, 54, -124, -113, 83, 70, -102, -20, 77, 116, -75, 63, -90, 25, 78, 13, -115, -82, -55, 5, -89, -113, -105, 51, 122, -67, 18, 67, -128, -18, 87, -11, 101, -102, -83, -117, -68, 55, 5, -81, 113, 25, -12, 84, 83, -15, -19, 116, -62, -11, 53, -78, 121, -48, 101, -127, 20, -86, 11, -112, -83, 102, -30, 41, 107, 18, -67, -86, 103, 124, 30, -78, 65, -72, -80, 63, -99, 2, 78, -98, 73, -61, -3, 89, 123, 40, 125, -114, 55, 45, 20, -106, 62, -12, 52, -104, 104, -95, -39, -73, 45, 121, -69, 99, -103, 81, 14, 103, 48, 4, -23, -80, -1, 39, 84, 110, -116, -76, -103, -74, -29, 103, -96, -41, -38, 114, 48, -71, 77, -21, -58, 114, -38, 99, 31, 77, 7, -113, 119, -92, 91, -38, 96, 68, -75, 78, -70, 114, 92, -78, 17, 113, 12, -89, -105, 8, -101, 33, -79, -78, -80, 18, -48, 49, -94, 56, -124, 44, 115, -46, -126, -27, 71, -14, -4, 18, -93, 17, 88, 4, 66, -88, 84, 0, -10, -28, -82, -61, -24, 97, 120, -40, 46, 112, 65, 89, 73, 43, -74, 26, -94, -48, -62, 105, -13, 71, -81, 123, -85, -47, 111, 119, 22, 55, -46, 125, 13, 21, -63, 68, -65, 25, 57, -78, -119, -14, -92, 16, -17, 0, -29, -5, -79, 46, -33, 40, -9, -90, 122, -75, 100, 61, -12, -86, 78, -103, 114, 122, -52, -65, 102, 99, 63, -6, -80, -91, 83, -5, 91, -32, -75, -53, 122, -95, 7, 5, -20, 112, 50, -83, 22, -85, 12, -29, 44, -103, -101, -84, -50, 122, -127, -32, -18, 72, 3, -126, 106, -93, 49, 55, -21, -18, 107, -114, -123, -128, -123, -76, 28, 95, -18, -79, -105, 109, 98, 18, -4, 71, 124, 3, 121, 69, -104, -109, -33, -21, -121, -75, -124, 15, 66, -123, 109, 69, -104, -74, -74, 105, -116, 50, -128, 93, -5, 124, -87, 19, 23, -66, 11, -16, 87, 3, -105, 115, 9, -15, -61, 73, -91, -16, 107, -113, 58, -77, 55, -114, 60, 45, -45, 10, -11, -65, 120, 95, -40, -128, -65, 62, 69, -76, -120, -17, -109, 124, 47, 118, -60, 86, 51, -76, -23, -103, 102, -16, 101, -115, -112, 61, 28, -95, 0, 45, -92, 2, -87, -29, -28, -53, -33, -57, 108, -92, -48, -63, -67, 86, 9, 37, 104, 23, 58, 124, -23, 126, 43, 74, -128, -92, -123, 23, 96, -121, 61, 25, 104, -12, 92, -68, 44, 85, -40, 67, 100, -124, -2, -17, 13, -50, 53, -123, -108, -50, -50, -66, -64, -101, 106, 34, -14, -42, -51, -46, 28, -35, -110, 124, 93, 98, -87, 10, 104, 33, 113, 120, 70, 49, -103, -59, 73, -121, 107, 49, -83, 14, -72, -33, -114, 30, 79, 40, -76, -99, -16, -104, 10, -39, 105, -85, 68, -96, -127, -17, -117, -22, 94, 126, 30, 102, 51, -63, -12, 82, -22, 117, -37, -99, -2, -114, -50, -49, -77, 125, 9, 110, 115, -44, -111, 103, 108, -74, 34, -54, 100, -61, 109, -4, -35, -75, 89, 17, 124, -16, 105, -27, 5, 104, 110, 43, 40, -77, 22, -16, 23, 108, 43, 49, 65, 7, 69, 49, -8, 58, 46, -126, 114, -39, -8, -60, 122, 67, -3, -125, 23, -34, -17, 53, 62, -83, 63, 8, -4, 102, 41, -12, -46, -82, -49, -39, 97, 37, -78, -95, 34, 112, -60, 68, -38, -68, 125, 48, 76, -111, 104, -85, -16, -36, -122, -102, 96, 51, -102, 56, 121, -100, -10, 91, -35, 126, -20, 4, -100, -87, 35, -116, 102, 75, -102, -122, 40, 76, 3, -114, -55, 101, 42, 21, 116, 14, -115, -103, -66, -100, -46, -33, 1, -6, -72, -61, -37, 16, -116, 113, -94, -46, 20, 95, -22, 48, -95, -111, -118, 87, 59, 41, -71, -122, 9, 44, -41, 118, 20, -115, 20, 110, -13, 31, -121, 33, 91, 13, -7, 56, 17, -101, -38, 8, 11, -92, 125, 93, 77, 55, -118, -48, 21, 57, -48, -18, -7, 53, -59, -102, 58, 103, -106, -101, 94, 118, 90, -5, -62, -37, -8, 85, -54, -95, -80, -55, 34, 102, -114, 108, 115, -95, 47, 30, 29, 96, 61, 59, -110, 29, -81, 62, -93, -127, -116, -62, 35, -81, 31, 27, -32, -69, -56, 62, -66, 36, -105, -68, 84, 59, 34, -107, -87, 46, -122, 84, 83, -80, 5, -36, 3, -98, -89, -117, -57, -49, 30, 18, -114, -122, -42, 55, -9, -108, 115, -92, 28, -79, -27, 42, 118, -63, 11, 93, 34, -31, -36, 69, 71, 110, -47, 42, 24, -44, 108, -15, 51, -119, 113, -70, 15, -119, 106, 65, -112, 25, 24, -70, -43, -34, -95, -28, -36, -44, -92, -47, 21, 106, -48, 64, -128, -92, -29, 55, -121, -108, -99, -90, 61, -120, 0, 89, -83, 9, -72, 10, 127, -56, 24, -119, -78, -94, 90, 31, 80, -103, -51, 82, 79, 9, 81, 64, -45, -74, -119, -58, -24, 88, -107, -66, 78, 73, 63, 28, -97, -78, 36, -16, 50, -64, -21, 66, -33, -77, 106, -95, 62, 43, 40, -102, 22, -120, -18, 36, 113, -51, -12, 71, -74, 41, 104, -40, 11, 5, 40, 104, -77, -9, 67, 1, -111, 96, 9, 57, 65, 116, 95, 62, 3, 121, 67, -76, -88, -22, -83, 94, -60, -39, 127, -14, 119, 72, -10, -37, 114, 104, 27, 44, -77, -119, -38, -99, 13, -23, 3, -14, -83, 54, 119, -114, -54, 104, 127, -54, 52, 126, 99, -52, 106, -17, -24, 111, -15, 62, -71, -15, 54, -71, -9, -62, -25, -31, -47, -56, -54, 62, -120, -67, 7, -65, 53, 102, 61, -1, 106, -32, -84, -97, 10, -107, -109, -100, -109, 109, 72, 4, 111, -110, 13, 10, -98, 68, -37, 45, 110, 99, 86, -93, -88, 63, -16, -59, -120, -84, -59, -104, 103, 96, -17, 40, 59, 50, -118, 107, 35, 2, 25, 7, -30, -128, 14, 75, -114, -94, 115, 51, -51, 94, 108, -24, 97, -128, -89, 16, -73, 109, -82, 127, 68, 74, -22, -118, 5, 32, 18, -85, -62, 4, 97, 46, -74, 84, -7, -35, 81, 87, -33, -89, 68, 73, -19, -111, 6, 30, 0, -62, 48, -58, -42, -67, -128, -30, -95, -125, 126, -38, -44, -108, -122, 84, 50, 56, 88, -86, -21, -60, -90, 12, 38, -120, 2, 44, 48, 101, -56, -63, 111, -4, 41, 124, 4, -50, 63, -58, -94, 24, 58, -64, -54, 34, -31, -48, -31, -14, -51, 115, 92, -73, 30, 61, 16, 119, -5, 57, 125, 59, 63, 44, 81, -79, 106, -58, -75, -64, 99, 88, -9, -5, 106, -99, -36, 0, 20, 63, 52, 14, -25, -91, -65, 63, 14, 20, -21, -94, -9, -114, 58, -29, -90, -14, -70, 100, -96, 3, 34, 15, -54, -121, -12, 33, 49, 13, -12, -24, -43, 62, 121, 40, -119, -75, 119, -30, -78, -120, -76, -111, 44, -57, 6, 65, -16, -14, 22, 65, -42, -75, 121, 43, 100, -93, 24, -94, 68, 58, -42, 110, 13, 7, 70, -10, 124, 6, 20, 41, 2, 73, -57, 113, 105, 41, -84, 119, 46, -25, 37, 108, -38, 22, 46, 98, 40, 43, -100, -116, 64, 36, -60, -10, -106, 42, 44, 48, 126, -12, 39, -125, -108, -28, -18, 17, -4, 58, -113, -48, -60, -40, -38, 86, 37, -32, -48, 120, -88, -127, 104, -70, 109, -69, -89, -71, 52, -127, -94, 68, 26, 31, -43, 51, -76, -108, -117, -29, 57, 90, -63, -31, -108, -57, 65, 57, -71, 17, 108, 15, 94, 77, 19, -3, -113, -23, -15, -19, 99, 112, 14, 76, -91, 54, 123, 50, -62, 78, 43, -29, -125, 120, -108, -95, 79, 30, -68, -87, -62, 21, -124, 19, 52, 26, -120, 90, -37, -44, 127, -80, -111, -114, -75, -22, 83, 111, -118, -112, 93, 48, -43, -50, -100, 5, -48, -59, 17, -29, 64, -56, 58, 11, 69, -1, 49, 1, 85, -98, -66, 65, 39, -3, 59, -14, -74, -6, -110, 83, -89, -23, 92, 48, -27, -97, 27, 2, -86, -112, 52, 81, 0, -43, -71, 126, 53, 100, -11, -6, 42, -100, -60, -13, -51, 33, 88, -35, -78, 63, 24, -94, 65, 43, -79, 51, 39, 49, 109, -40, -26, -14, 24, -2, -108, 50, 4, -47, 105, -37, -47, -125, 99, -119, 17, 63, -99, -117, 54, 66, 111, -125, 52, -88, -5, -19, -39, 75, 46, -125, -22, -125, 41, 82, -93, -99, -105, -57, -106, -95, 51, -124, 49, 77, 115, 28, 53, 43, -108, -58, 8, -43, 78, 28, -19, -17, -103, 50, -46, 72, -35, -103, 18, -21, 24, 61, 13, 25, 113, 108, 116, 76, -83, -57, -92, -35, 72, 47, 79, -114, -118, 71, -108, -54, 50, -105, -118, -35, -94, 37, -99, 73, 29, -18, -63, 56, 58, -99, -83, -118, 98, -50, 35, -100, -11, -105, 1, -54, 81, 21, 55, 97, -111, 12, -17, 124, 104, -3, 32, 116, 26, 97, 98, -71, -17, 123, 24, -124, 113, -126, 39, -91, -35, 51, 38, -6, 94, 125, 106, 79, 15, -26, 3, -63, 115, -54, 21, -94, 38, -89, -55, -97, 85, -102, 7, 121, -81, 66, -3, 111, 114, 88, 78, -117, -22, -10, 29, -49, 89, 8, 108, 79, -113, -116, -83, 41, -50, -7, 91, 126, -48, -118, 16, 104, -81, -115, -13, 94, 22, 110, -118, -50, -75, -12, -99, 58, 8, 34, -15, -122, 70, -46, 15, -5, 109, 107, 100, -30, -101, 118, 95, 91, -121, 69, -33, 96, -107, 9, -69, 71, -45, -115, -5, -67, -41, 97, -69, -83, 119, -84, 23, -16, -15, 101, 57, -61, 112, -54, -74, 30, 84, -52, 9, 117, -88, -75, -74, 1, 2, 70, 87, -18, -128, -50, 11, 81, 124, -27, 95, 15, 83, -43, -32, 80, 32, -28, -31, -98, -110, -4, -102, 42, 125, 99, 124, 81, -113, 5, -117, 74, 60, 46, -59, 106, -32, 7, -30, -40, 94, 39, -42, 106, -14, 96, 99, -92, -10, -90, -76, -16, -2, -74, -24, -75, -26, 106, 12, -22, 119, 86, 97, -115, -118, 124, 115, -104, -112, -65, -7, 51, 20, 17, 116, 99, -43, 118, -64, -66, -55, -93, -42, -70, -88, -111, 3, -13, 62, -55, 12, -69, 85, -128, 90, 110, -20, -67, -86, 11, -119, -11, -82, 102, 11, 75, 24, -33, -54, 48, 38, -124, 51, 36, 63, 48, 36, 109, -125, 19, 45, -58, 79, 111, 55, -64, 46, 110, -128, -17, -61, 63, 114, -38, 34, -11, 9, 54, 90, -7, 96, 84, -45, -24, 79, 79, 118, -97, 70, -29, 1, 1, 93, -122, -63, 63, -107, -118, 89, -37, 0, -85, -4, -112, -15, -18, 86, -100, 123, 19, 11, 125, 122, 118, 65, 122, 102, -61, 119, -62, 70, -75, -59, 11, -84, -70, 49, -127, -24, 43, -14, 10, -81, 82, -8, 126, 6, -75, 45, -108, 41, -115, -66, 103, 15, -21, 69, 89, -74, 121, -1, -73, 80, -83, 95, -109, -106, 80, 70, -67, 33, -127, 116, -49, 106, 45, -23, -32, -118, -42, -77, 16, 105, 87, -22, -33, 112, 104, -69, -116, -34, -68, -79, -39, -124, -72, 30, 60, -32, 119, -92, 89, 77, -87, 5, -89, 73, -64, -93, 2, -81, 96, 127, 14, 12, 90, -41, 48, -45, -9, 124, 70, -72, 111, -66, -114, -86, -9, 61, -87, 105, -121, -38, 22, 6, 13, 67, 67, 45, -2, 127, 118, -66, 6, -105, -11, -3, -85, -15, 56, 101, -50, 54, -31, 98, -29, 55, -25, 100, 113, -4, 40, 110, -104, 78, -31, -100, -90, 12, 117, 101, 53, 55, -38, 111, 74, 96, -103, 37, -77, -100, -29, -46, -88, 48, 122, -84, -12, -19, -107, -47, -117, 45, -25, 78, 121, -48, -68, -111, -112, -115, -64, 86, -112, -46, -54, -53, -64, -124, 29, 6, 81, -98, 60, -6, 102, 13, 30, -104, -118, 14, 20, 0, 104, -86, -7, -77, -16, 68, 42, -67, -23, 33, 122, 91, 16, 42, 57, 41, 77, 55, 25, 90, 66, 119, -56, -67, 72, -92, -54, -83, -47, -13, 123, 39, 34, 39, 123, 40, 74, -99, -48, 11, 89, 15, 21, -8, -85, -16, -87, 20, 56, -15, -38, 18, 55, 24, 14, 96, 57, 84, 5, -111, 57, 13, 20, 105, 76, -102, -31, 98, 99, -62, 35, -17, 108, 65, -22, -28, 92, -17, -5, 122, -96, 109, -23, 79, -13, 56, -68, 114, -65, -50, -117, 58, 120, 127, -72, -127, 51, -54, 106, 118, -32, 47, -68, 2, 49, -52, 56, -114, -79, 54, -90, 124, -40, -40, -70, -37, -39, 79, -96, -85, 125, -40, -82, -120, -40, 107, 84, 44, 84, -5, -34, -12, -71, 11, -81, -64, 90, -19, -65, -126, 110, -6, 22, -8, 109, -112, -8, -98, -101, 90, 123, -48, 87, 120, 122, 80, 22, -24, -29, -101, 91, -26, -43, 29, 61, 110, 78, -20, 12, -35, -17, 109, -30, -73, -81, -103, -73, 71, -72, -73, 123, -40, -29, 77, 40, -7, 98, -5, -99, 101, 2, 95, -21, 28, 65, 94, 100, -94, 59, 84, 99, -40, 73, 47, -6, -48, 38, -28, -124, 19, 109, 79, 103, 46, -56, 99, 9, 26, 58, -87, -51, 64, 59, 49, 100, 85, 105, -43, -54, -68, -49, 82, -14, 57, -83, -70, -99 );
    signal scenario_output : scenario_type :=( -39, 26, -23, -19, 28, 82, -22, -25, -13, -48, 28, 41, 8, 9, 3, -64, 59, 19, -7, 41, 38, -64, -9, -62, 9, -44, 89, 14, -14, 1, 27, -61, 11, -29, -60, 63, 64, 80, 35, -11, -90, -69, -20, 48, -19, 53, 51, 46, -47, -48, -82, 31, -23, 28, -31, 18, -74, 30, 22, 46, -32, 79, 34, -57, -44, 82, -12, 1, 93, 6, -93, -8, 1, -23, -1, -11, 6, -3, -1, 13, 0, -55, 26, 32, 17, 32, 30, -27, 30, 2, 21, -13, -14, -39, 66, -53, 24, -15, 8, 14, 85, -40, 24, -14, -39, -42, 71, 28, 29, -23, -128, -68, 83, 31, -54, 8, -19, -80, -17, 71, 78, 52, 36, -18, -23, 0, -35, -106, 36, -11, 31, -28, 13, 14, 112, -26, 10, 24, -37, -76, 8, -24, -38, 66, 11, -62, -6, 12, -17, -47, -38, -59, 30, 127, 59, -59, -31, -12, -40, -31, 24, 46, 80, 1, 23, -2, -23, -42, 23, -14, -23, -43, 5, 65, 29, -11, -9, -71, 38, 13, -2, 21, 49, -30, 97, 5, -37, -5, -47, -20, 102, -26, -56, 73, -34, 3, -30, 0, 34, 80, -17, 38, 32, -25, -47, -34, 28, -47, -28, -60, -49, 8, 97, 91, 45, -14, -7, -43, -87, 14, 51, -68, 43, 26, -93, -73, 36, 69, 102, -8, -76, -9, -4, -31, 0, -3, -7, 14, -4, 76, 59, -65, -60, 30, 3, 9, 12, 39, -46, -34, -19, -22, -49, 86, 15, 57, -8, 42, 45, 19, -96, 36, -18, -27, 0, -40, 13, 59, 1, 3, 32, -44, 28, 17, -35, -24, 70, -37, -15, 25, -69, -36, 48, 45, -14, -44, -11, 4, 66, -12, 6, -45, -12, -78, 56, 44, 44, -14, 58, -26, -61, -64, 38, 20, 1, -26, 13, -19, 7, 10, -12, 41, 10, 21, -12, -35, -100, -6, 73, 112, 25, -78, -25, -19, -24, 19, 103, 45, -28, -39, -8, -27, 0, 127, -22, -41, -54, -65, -68, 29, -23, 51, 45, 38, 62, 61, -96, -34, -72, -23, 88, 96, -43, -15, -27, 18, 39, 27, -93, -25, 75, 12, -83, 25, 21, -12, -2, -12, 5, 14, -14, 22, 42, 10, -23, -26, -2, -3, -63, 32, 23, 51, 0, 71, -61, 14, 24, -14, -80, -5, -39, -3, 59, 51, 42, -21, -57, -25, -21, 8, 35, 39, -51, -2, 3, 34, 55, -12, -9, 19, -91, 0, 82, -40, 21, 12, -11, -22, 80, -54, 8, -71, -10, -62, 97, 36, -23, -35, 8, 43, 17, -73, -23, 85, 74, -9, 2, -102, -42, 32, 71, 14, 61, -17, -1, -15, -81, 20, -10, -36, 36, 19, -2, 43, -83, -59, 7, -78, 21, 27, -9, 20, 109, 59, 28, -92, -26, -23, -58, -4, 11, 8, 32, 40, 3, -30, -82, 96, 22, -36, 68, 57, -128, 12, 39, -63, -45, -4, 19, 51, 90, -14, -9, 31, 8, -87, 22, 32, 6, 58, -35, -30, -70, -52, 59, 27, -60, -45, -24, -3, 54, -13, -4, 1, 81, 58, -7, -106, 19, 10, 56, 43, 6, -65, 13, 2, -13, -73, 31, 65, -2, -51, -46, -23, -21, 54, 64, 102, -9, -8, -106, -38, -25, 24, 94, 64, -71, 18, 66, -48, -55, -42, -9, 86, 90, -32, -74, -38, 12, 73, 2, -12, -27, 8, 0, 38, -5, -12, -47, 27, 25, -65, -24, 119, -15, -60, 32, -30, -5, -6, 23, 31, 54, -73, 18, -13, 52, 47, -18, -45, -82, -57, 42, 24, -28, 42, 56, 56, -28, 9, 30, -62, -47, -4, -59, -35, 25, 30, 19, 32, -47, 60, -37, 55, -48, 57, 19, 116, -73, -6, -74, 1, 7, 0, -73, 25, -11, -52, 51, 20, 71, 11, 0, -1, 48, -51, 95, 1, -48, -10, -83, -53, 92, -26, 29, 23, -52, -55, 98, 0, -34, -69, 9, 20, 116, 66, -32, -79, -29, -56, -29, 27, 126, -8, -3, 39, -8, -69, 26, 19, 39, 11, -74, -70, -4, 15, -13, 51, 108, -8, -83, 30, -34, 20, 29, 21, -37, 18, -40, -12, -66, 56, 57, -43, -7, 2, 19, 74, -51, 9, 62, -71, -24, 2, -53, 41, 78, -35, -7, 91, 42, -61, -91, 32, 22, 17, 3, 9, -59, -19, 62, 48, 60, 48, -32, -51, 32, -46, -38, 59, -61, -37, 26, -21, 58, 22, -77, 43, 4, -116, 34, 48, 28, -13, 28, -22, -29, -58, -18, -40, 68, 30, 52, 37, -28, -4, -8, -31, 60, 30, 6, 29, -35, -59, -24, 46, 22, -111, -13, 75, -19, 20, 51, -55, -106, 17, 10, 65, 64, 19, -97, -27, 36, 40, 24, -37, -37, -27, -31, -20, 66, -12, 45, 76, -17, -46, 24, -38, 11, 29, -56, -14, 34, -29, -8, -8, -26, -12, 6, -1, 17, 3, 43, 3, 10, 63, 51, -9, -25, -19, -28, 62, -3, -22, -10, -29, -26, 20, 61, 17, -92, 6, 40, -23, -61, 14, 26, 81, 25, 30, -2, -69, -40, -45, -18, -13, 29, -11, -47, 70, 82, 42, 4, -1, -72, 41, 30, 34, 87, -41, -61, -7, 34, 19, 27, -95, -49, -3, -36, 13, 102, 42, -59, -24, -7, -8, 63, -36, -5, -46, 19, 23, 17, -109, 63, 14, 7, -49, 41, -42, 71, -35, 21, 27, 14, -87, 48, 18, -74, -15, 10, -19, 90, 39, -9, -71, -6, -46, 24, 68, 36, 10, 8, 27, 11, 31, -128, -53, 72, 0, 11, -2, 0, -63, -2, 6, 52, 19, 17, -14, -12, -1, -86, -77, 6, -22, 31, 32, 51, -92, 72, 12, -22, -43, 26, -34, 73, 30, 18, -5, 26, 4, -3, -43, 31, -34, -41, 20, 4, 17, 38, 72, -41, 5, -20, -11, -72, -18, 10, 45, 3, -80, -31, 66, 75, -12, -43, -17, 34, 26, -37, -88, -27, 15, 62, 44, -8, -12, 39, -10, -44, 37, -46, 2, 9, 0, -69, 80, -3, 19, 9, -5, 6, 37, -36, -60, 8, 22, 4, -54, 112, -59, -13, 42, 38, -94, 28, -17, 72, -28, -29, -70, 57, -6, 23, -19, -31, -59, 63, -20, 4, 41, -6, -66, 73, 20, 0, 51, -11, -29, -24, -34, 0, 127, -5, -3, -71, -44, 39, 17, -17, -1, -19, -79, 36, -24, 62, 38, 12, 9, -10, -60, 45, 34, -23, 40, -27, -61, 85, 14, -81, -36, 41, -30, -44, 22, 6, -34, -31, 28, 60, 93, 0, -47, -42, 71, 26, 12, -43, -20, 30, 25, -103, -29, 25, 47, 55, 10, 58, -25, -108, 31, 4, -55, -7, 13, 11, 80, -57, -10, -21, -43, 53, 68, -49, -90, 24, -12, -70, 34, 91, -11, 61, 13, -2, -18, -4, -77, -2, -29, 117, 28, -31, -64, -27, -55, 17, 59, 102, 56, 61, -68, -104, 5, 36, -65, -44, 70, 20, 45, 29, -3, 17, -14, 3, -17, -18, -92, -6, -59, -1, -15, -38, 9, 127, 43, 27, 5, 29, -31, -52, -93, 104, -8, 32, 31, 44, -61, 2, -11, -28, -128, 29, 70, 0, -3, 21, 17, 71, 19, -98, -54, -53, 9, 92, 3, -51, 69, 46, -71, -8, -10, -1, 71, 59, -66, -32, -18, 80, -2, -43, -3, 56, -57, -53, 31, 1, -36, 20, 32, -31, -37, -31, 30, 79, 74, -13, -34, -36, 59, -12, -38, -96, 45, 8, 47, -40, 36, 4, 41, -31, 12, -82, 1, 38, 70, 22, 59, -21, -36, -7, 30, -30, -69, -48, 63, -22, 34, 28, -104, -51, 63, -10, 27, 43, -81, -1, -10, -34, 81, 22, -126, 36, 9, -14, 96, 29, -61, -23, -57, -23, 44, 42, -1, -14, -66, 43, 4, -28, -25, 86, 1, -81, 0, 5, -1, 79, 28, -128, -4, 5, -64, 26, 77, -63, 0, 12, 13, -28, 24, -106, 30, 86, 70, -63, -8, 6, -48, 6, 72, 95, -47, 6, -5, -15, -23, -8, -92, -23, 42, 49, 81, 55, -2, -60, -56, 41, -18, -46, -74, -44, 25, 82, 22, 47, -43, -66, 21, 11, 47, 35, -87, -35, 32, 59, 0, -52, -89, 1, 14, -19, 31, 18, -78, -29, 104, 34, 37, 54, -54, -52, -63, -74, -28, 64, -5, 39, 96, -43, -20, 2, 47, 9, -7, -41, 46, -2, 47, -51, -34, -10, -53, -32, 85, -60, 4, 78, 75, -15, -25, -94, 40, -1, 31, 60, 0, -93, 25, 0, -25, 6, 41, -11, -17, 17, -8, 6, -18, -22, -8, 83, -53, -49, 28, 20, -30, -49, -49, -31, 57, 99, -6, 14, -28, 24, -60, 17, 1, 93, -8, -75, -44, -17, 8, 83, 41, -36, 42, 10, -122, -37, 38, 43, -26, 4, 40, -6, -111, -20, 106, -34, -14, 108, -21, -53, 23, -29, -39, -5, -42, 63, 55, 30, -7, -1, -44, -31, -45, 63, -41, -39, 0, 22, -34, 1, -45, -6, 32, -47, 0, 105, 39, 34, 62, -58, -64, -56, -24, -45, -23, 19, 93, 44, -51, 34, 39, -62, -30, 56, 28, -52, 42, -23, 8, 15, 54, -60, 7, 26, -14, 14, 17, -74, -91, -10, -27, 11, 39, 42, -10, 51, -6, -48, -24, 54, 1, 69, -28, -72, 12, -6, -3, 29, 3, 0, 68, -57, -86, -20, -23, 36, 20, -25, -51, 3, 28, 93, 59, 35, -25, -110, -34, 32, 9, -30, 38, -30, 11, 6, -13, -41, 69, 26, 61, -24, -71, -34, 44, -72, 21, 23, -35, -69, 75, 31, 72, 10, -30, -54, -30, -53, -24, 79, 21, -76, 31, 48, -31, -40, -22, -4, 53, 42, 52, 65, 45, -40, -60, 13, -52, -26, -4, -31, -10, 94, 28, -1, -47, -29, -9, -31, -52, -17, 71, 62, -20, 7, -31, -44, 0, 70, -30, -38, -6, 13, 102, 21, -19, 7, -38, -29, 49, -7, -58, 40, 8, 1, 28, 105, 18, -62, -31, -11, -45, -97, 56, 48, 12, 30, 37, -62, 14, -3, 21, 36, -11, -65, 31, -42, 21, 44, 57, 39, -14, -56, -94, 27, -43, 70, 12, 71, -23, 26, -128, 8, 88, 35, -27, 56, -34, -71, -3, 13, 64, 29, -24, -2, -53, -42, 21, 24, -20, 68, 46, -29, -58, 11, -35, -22, 54, 14, -9, -14, 14, 9, -15, 58, 45, -22, 26, 9, -18, 7, 10, -61, 38, 43, 13, -28, -65, -31, -74, -11, 69, 60, -47, 21, 89, -25, -80, 41, 8, -34, -38, 47, -64, 8, 59, 52, -41, 21, -53, -26, 39, 6, -55, 73, -37, 5, 43, 96, -10, 32, -9, -70, -39, -5, 32, -56, 22, -12, -12, -29, 111, 79, -73, -28, 44, -36, -51, 72, -34, -18, 48, -20, -88, 41, 32, -27, -37, 8, -48, -29, 42, 74, 47, 41, -22, -17, -83, 54, 21, -11, -47, 56, 31, -5, -49, -43, 51, 96, -21, 15, -69, 1, -46, 4, -75, 76, -7, 34, 5, -61, -28, -34, 4, 96, 73, -51, -25, -65, -27, 92, 108, -38, -34, -29, 23, -29, -6, 0, 31, 60, 35, -65, -81, -13, -30, 23, -8, 44, 48, 58, 19, -28, -24, 47, 65, -22, -45, -49, 57, 14, -29, -68, -53, -2, 72, 104, -14, -22, -59, 0, -54, 12, 36, 56, -82, -7, -3, 28, 43, -2, -55, 22, -2, -78, -37, 5, 26, 100, -11, 1, -48, -6, 45, 71, -61, -25, 15, -35, -45, 15, 81, 0, -39, 14, 61, 42, -36, -40, 99, -28, -44, 30, -34, -6, 54, -35, -31, -26, -86, 18, 42, 10, 38, 65, 65, -49, -61, -12, -47, 2, 63, -31, -98, 9, 42, 22, 20, 27, 26, -41, 27, 8, 71, -30, -10, 6, 2, -77, 49, -20, -35, -11, 25, -17, 20, 10, 27, 14, 9, 24, -55, -5, -32, -29, -39, 66, -21, 24, -18, -37, -41, 77, -34, -8, 46, 17, 4, -12, -43, 41, 10, -100, -46, 38, 9, 14, 79, 25, -48, -76, -22, -55, 25, 94, 34, -20, -8, -25, -92, -15, 26, 86, 10, 47, -12, -46, -57, 56, 3, 107, -24, 22, -96, 29, -53, -9, -60, 119, 37, -41, -26, 43, -48, -53, 38, 2, 20, 35, 38, 46, -20, -94, 25, -11, 13, -1, 28, -30, 62, -87, -31, 61, 40, -76, -39, -9, 37, 8, -35, 64, 32, -108, 6, 12, 1, 4, 52, 53, 7, -11, -7, -55, -24, 65, -15, 6, 39, -9, -110, -55, 73, 11, -34, -3, -39, -37, 1, 25, 51, -27, -19, 64, -13, -39, -28, 47, -2, -8, -39, -6, 36, 91, -54, -9, 39, 28, 40, -49, -74, -10, 29, 17, 66, 2, 40, -58, -115, -47, 85, 41, -19, -25, 21, -7, -48, -49, 62, -51, 0, 64, 104, -58, -30, -72, 8, -42, 13, 51, 82, 18, -42, -45, -53, -35, 28, 106, 31, -6, -17, 3, -18, -77, 31, -11, -51, -42, 14, 9, 30, 53, 4, 36, 34, 18, -30, 9, 38, 11, -87, -53, -44, -112, 10, 127, 2, -23, 40, -47, -86, 37, 82, 75, 2, -40, -56, -38, 2, 75, 77, -23, -60, -36, 8, 7, 65, 36, 35, -19, -57, -90, -22, -9, 66, 37, 47, -6, -35, -38, 43, -13, 35, 35, -20, -83, -24, -8, 47, 0, -51, -26, 7, 20, 20, 58, 51, 2, -114, -85, 2, 43, 18, -30, 0, -29, -5, 48, 43, -44, -5, -54, -29, 18, 97, -68, 19, -4, -2, -29, 90, -17, 64, -49, -32, -41, 79, -55, 20, 14, 44, -15, -72, -6, 10, 22, -22, 12, 17, 103, -77, -48, 0, 82, 13, 46, 5, -103, -82, 76, -5, -19, 12, -55, -24, 91, 81, -29, 2, -44, -66, 40, 37, -36, -36, -28, 42, 52, -2, -58, 39, -11, 38, 3, 9, -39, 21, -60, 34, 60, 12, 29, 28, -51, 74, 40, -68, -18, -7, -51, 17, -22, -14, 31, 69, -42, 55, -14, -87, -9, 99, -37, -49, 12, 15, 13, 62, 24, -83, -44, 114, -42, 26, 42, -53, -17, 49, -34, -8, -39, -53, 37, 21, -27, -9, 70, 52, -27, 46, -28, -66, 76, 60, -43, -14, 44, -15, -90, -25, 82, 20, -6, 9, -77, -2, 41, 28, 15, 20, -44, 21, 72, -19, 12, -18, -26, -43, 83, -46, 8, -83, 23, -73, 24, 48, 46, -15, -14, -25, -6, 71, -36, -21, 1, 43, -25, -47, -45, -23, 62, 63, -37, 14, -37, -23, -14, 39, -19, 59, 65, 11, -51, 8, 14, -3, -26, 24, -58, -18, -11, 80, 3, -22, -73, -12, -21, 103, 42, -28, 47, -11, -105, -36, -4, -32, 27, 93, 18, -83, 37, 60, -35, 41, 8, 14, -40, 36, -39, 40, -27, -26, -53, 71, 23, -7, 17, -2, -2, 18, 18, 10, -71, -39, -10, -27, -30, -32, -71, 59, 39, 44, -19, -8, -21, 42, -21, -25, -34, 44, 79, -62, 0, -7, 40, 32, 3, -99, -78, -37, 42, 105, 73, -1, -107, -1, 80, -19, -3, 37, 42, -37, 15, -7, -11, -77, -80, 5, -5, 35, 61, 63, 26, 47, -99, -88, 35, -1, 1, -1, -20, 8, 19, 43, -19, 1, -30, -45, -19, 93, 49, 11, -15, -35, -93, -23, 56, 26, 9, 37, -41, 43, -45, 0, -36, -13, 44, 123, -71, -72, -42, 6, -26, 22, 38, -17, -28, 56, -17, -46, 22, 127, 22, -69, -76, 23, 38, -20, 10, 106, -4, -119, -10, 15, 0, 12, 21, -10, -20, -9, 35, 58, 14, -1, -103, -27, -51, 68, -6, 12, 21, 63, 9, -11, -27, 20, -15, -77, 41, -55, -20, 13, 47, 29, 40, -36, 2, -38, -18, 40, 9, -5, -46, 24, 25, 0, -99, 12, -12, -28, 1, -13, 34, 26, 21, -3, 51, 39, 78, -66, -22, -13, 19, -2, 46, -108, -62, 27, 76, -61, -65, 9, 26, 43, 75, 7, 17, -42, -69, -64, 73, -85, 42, -2, 24, 3, 39, -42, 11, -34, -41, 27, 39, 15, -57, -46, 57, 29, -57, 1, 2, 11, 18, -58, -27, 121, -14, 8, 86, -5, -86, -21, -79, 44, 58, -47, -28, 95, 9, 9, -41, -22, 19, -3, -48, -55, -22, 127, 54, -44, 31, 24, 14, 14, -7, 45, -19, -123, -17, 20, 12, -6, -59, -58, 15, -25, -36, 77, 7, 38, 14, 24, -56, 97, -34, -3, 9, 38, 9, -55, -15, 7, -80, -12, 82, -32, -19, 83, -90, -24, 115, 36, -116, -3, 55, -18, 35, 32, 20, -64, 23, -6, -19, -39, -29, -26, 85, 13, -22, -11, 6, -7, 23, -44, -29, -36, -4, -17, 44, 100, -13, -51, -31, 56, 21, 9, -89, -15, 76, 44, -63, 48, 43, -107, -7, 68, -12, -69, 8, 4, -9, -42, 45, 20, -7, 22, 74, -22, 45, -35, -51, -23, 65, -57, -37, 3, 63, -26, -29, 46, 29, -92, -5, -2, 17, 18, 27, 11, 8, -38, -13, -63, -19, 62, 34, 45, -18, -21, -58, -3, -23, 44, 34, 55, -128, -43, 95, 6, -89, 11, 11, -2, -12, -26, -32, 46, -11, -56, 86, 45, 14, -24, -23, -5, 88, -37, 38, -6, -46, 38, 34, -44, -37, 10, 18, 78, 4, 4, -111, 7, 8, 0, 30, 19, 13, -12, -42, 35, 34, -76, 0, -34, -54, 57, 105, 15, -58, -25, -52, 9, 66, -5, 19, 30, -115, -32, 77, 86, -1, 19, -76, -32, -6, 31, -43, 23, -7, 2, 109, -18, -17, 4, -1, -10, -24, -21, -27, -51, 45, 68, -71, 4, 53, -37, -17, 65, 21, -48, -45, 0, 44, 59, 9, -54, 1, -2, 12, -24, -3, -45, 27, 60, 94, -28, -28, 1, 63, -38, -40, -26, 15, 1, -17, -54, -23, 27, 41, 6, -8, 19, 25, -45, -64, -26, 29, 56, 5, 8, -63, -95, -12, 15, -3, -41, 78, 24, -27, 26, 95, 18, 52, -17, -128, -61, 9, 71, 73, 4, -44, -65, -69, 39, 68, 14, -4, -60, -45, 12, 49, 28, 15, -5, 52, 26, -48, -40, -49, -34, -38, 109, 15, -36, -34, 94, -41, -39, 15, -22, -106, -6, 45, 45, 1, -7, 66, 17, 0, -65, -77, 18, 60, -47, -2, 110, -9, 59, -1, -9, -54, 2, -28, 53, -17, 15, -22, -24, -34, 18, -5, -56, -66, 58, 52, -56, -13, 94, 94, 0, -15, -77, 1, 38, 44, -85, -32, -23, -7, 51, 9, -36, -10, -37, 25, 98, 35, -32, -23, -59, -66, 66, 87, -34, 21, 53, 25, 56, 6, -128, 9, -30, 31, 69, 9, -102, 64, 8, -12, 49, 66, -39, -25, -28, -89, -21, -3, 29, 56, 124, -42, -22, -77, 11, -11, 95, -35, 1, -60, -18, -2, 85, -19, 9, 2, -63, -18, -18, 13, -8, 56, -79, 11, -72, 60, -14, 4, -69, -9, 13, 78, -9, -48, 2, 51, 30, -57, -17, 34, 29, -5, 1, 35, 9, -128, 4, -48, 25, -7, 77, -28, 10, -39, 71, -100, 22, 63, 15, 1, 112, -21, -117, -59, 72, 30, -30, -70, 26, 27, -41, 43, -3, -9, -8, 46, 19, 37, -81, -37, -1, 52, 13, -12, 51, 1, -110, -47, 1, -13, -44, 22, 4, 44, 56, -13, -34, -10, -53, -17, 7, 17, 21, 8, 64, 90, -54, 6, -3, 13, -39, 23, -39, 51, -13, 46, -23, 10, -88, 3, 24, 62, 19, 2, -82, -10, 39, -26, -17, -11, 23, -2, 38, -22, 1, -28, -18, 6, -25, 40, -2, 48, -35, -53, -17, 104, -39, -1, 55, 32, -114, 9, 38, -82, -6, 27, -27, 49, 14, -47, 48, 51, 35, -10, -128, -6, -6, -19, 43, 95, -66, 3, 15, -66, -23, 64, -40, -98, 54, 5, -34, -13, 90, 9, -30, -24, 17, 1, 15, 8, 53, -31, -7, -27, 75, 15, 81, -29, -30, -18, -31, -72, -35, -10, 11, 40, 42, 28, -60, 11, -4, -25, 41, 75, -15, 2, 2, 29, -2, -4, 8, 15, 1, 22, 0, -14, 38, -53, -8, -60, -8, -39, 58, 0, 80, -89, 5, -28, -3, -24, -4, -70, 36, -49, 26, 45, -20, -8, 82, 18, -40, -30, -9, 109, 39, -106, -28, 87, -53, -9, 68, 21, -90, -28, 5, 18, -37, 13, -8, -11, 0, 78, -2, 29, -65, 76, -27, 5, 21, 64, 2, 2, -73, -25, 18, -71, 46, 18, -42, -6, 64, 28, 9, -4, -86, -13, 23, -23, -51, 109, 34, -51, 3, 100, -15, -58, -38, 0, -55, -40, 7, 115, 44, -79, -2, 69, 49, -62, 30, -60, 7, -36, 76, 4, 27, -114, -45, -47, 65, 90, 28, -47, 15, 10, -30, 46, 63, -108, -25, 104, -36, -10, 32, -17, -28, 6, 15, -7, 5, 12, 9, -19, -7, 3, -13, 6, 0, 107, 0, 18, -85, -47, 12, 31, -23, 34, -3, 0, -13, -7, 37, 25, -31, -65, -6, -11, 3, -57, 12, -39, 45, -48, 54, 15, 19, 3, 7, -17, -53, 44, -36, 10, -32, 78, -19, -11, 43, 24, -60, -89, 15, -52, 49, 30, 58, -4, 113, -18, -117, -15, 20, -82, 35, 51, -73, 81, 11, -24, -5, 3, -31, 61, -48, 38, -2, 14, -46, -40, -12, 105, 18, -56, 1, 30, -31, -27, 90, -28, -43, 59, 37, -64, 18, -44, 3, 36, -31, -51, 53, -1, -11, -43, -17, -29, 91, 34, -9, 75, 7, -107, 2, -55, -26, 121, 38, 7, 36, -77, -27, 19, -52, -89, 53, -35, 39, 32, 38, -26, 89, 22, -58, -35, -73, -30, 65, 61, -52, 54, 9, -3, -25, -9, -29, -12, 0, 64, 34, 28, 17, 13, -13, -117, -35, -1, -59, 3, 99, 28, -19, -42, -36, -13, -52, 29, 9, 36, -18, 35, 20, 87, 64, 34, -81, -128, 22, -14, 62, -42, 80, -65, 51, -21, 29, -76, 25, 57, 42, -76, -19, 55, -39, -96, 2, 93, 52, -12, -47, -27, 11, 24, 0, 100, 2, -52, 14, 28, -58, 7, 7, 36, -39, -79, -69, 25, 10, 48, 25, -45, -61, -76, 11, 93, 56, -36, 30, 10, -11, -23, 10, 5, -11, 6, 92, 49, -53, -61, -54, -30, 52, 32, 15, -70, -14, 46, 104, -36, -44, 0, 48, -7, 18, -36, -53, 12, 75, -26, 9, -10, 34, 14, -70, -17, -8, -46, 10, 26, -102, 15, 37, 41, 74, 72, -12, -98, -11, -1, -52, -46, 20, 59, 51, -59, -92, -3, 45, 78, -46, -12, -48, -11, 64, 72, -46, -27, -44, -77, 49, 30, 73, 56, -39, -77, 62, 27, -49, 22, -88, 1, 47, 92, -29, -63, -19, 69, -18, -90, 61, 3, -28, -25, 27, 0, 91, 44, -3, -1, 40, -44, -104, -31, 15, 52, 18, 22, -52, -11, -20, 55, 34, -14, -61, 2, -31, 20, 34, 35, -44, 29, 25, 49, -21, -9, 28, -6, -74, -46, 40, -14, 13, 3, -55, -37, 37, 3, -32, 0, 83, 22, -2, -58, -14, 43, 81, -6, -26, -66, 47, 32, 0, 31, -3, -17, -29, -18, -52, 68, 18, -34, 43, 18, -19, 3, 100, 7, -18, -90, -24, -19, -52, 27, 52, 62, 47, -9, -89, 35, 6, -11, 6, 38, -2, -39, -8, 18, -14, -72, 1, 37, -2, -3, 45, 102, 47, -38, -73, 8, 22, 11, 38, -23, -36, 7, -25, 18, -4, -13, 13, 26, -65, -39, -3, -6, -17, 22, 4, 15, -8, -5, -103, -1, 18, 53, 30, -27, -22, 4, -44, -17, 112, -39, -76, 8, -51, 13, 74, 53, -103, -12, 40, 20, -12, 102, -2, -73, -37, -15, -27, 26, 26, 31, 44, 7, -15, -9, -17, -121, 35, 36, 6, 10, 61, -44, -1, -18, -47, 17, 14, 51, 0, -35, -25, 8, -11, 77, 93, -96, 38, -26, -25, 26, 15, -83, 28, -1, -90, 14, 94, 100, 29, -86, -19, 21, -27, -99, 85, 19, 9, -74, 74, -26, 32, 48, 6, -53, 62, 23, 4, 0, -17, 24, 46, -54, -68, -62, 27, -8, -29, 39, 111, -22, -63, -3, 44, -38, -64, -10, 15, 25, 76, -26, -38, 1, 40, -19, 41, -73, 9, -21, 42, -17, -11, -20, 81, 94, -26, -9, -74, -17, -77, 6, 18, 47, 27, 25, -41, -96, 26, 54, 51, -66, -35, 17, 14, 68, 71, 20, -72, -36, -63, -60, 48, 103, -57, -77, -10, 22, 55, -23, 17, -35, -9, 72, 58, -27, -22, -6, -2, 89, -3, -51, -42, 41, 0, -25, -70, -36, 11, 98, 5, 21, -17, -53, -79, 62, -37, 26, 65, 0, 1, 68, -13, -77, -23, 39, 72, 40, 0, -70, -94, -7, -14, 45, 47, 37, -10, -1, -39, 47, -36, 26, -4, 71, -42, 35, -47, 12, 6, 38, -6, 13, 37, -75, -47, -22, 4, 31, 19, -76, -32, 72, -34, 25, 49, -5, -97, 6, -31, -3, 8, 83, -20, -23, 34, 96, -31, -22, -69, 35, -44, 1, 53, 41, -128, 1, 69, 15, -20, 4, -27, 3, -18, 49, 35, -1, -85, 2, 7, -26, 25, 40, -21, -2, 24, 0, -2, 56, -1, 62, -1, -28, -116, 0, -3, 75, 35, -4, 17, -47, -30, 30, -43, -64, 119, 52, -55, -58, -48, 14, 19, 64, 0, 47, -48, -8, 6, 102, -77, 0, -10, -79, -19, 8, 1, 64, 95, -47, -29, -52, -11, 26, 28, 10, -69, 1, -39, -3, 28, 81, 29, 59, -25, -28, -42, -82, 1, 47, 29, -9, 42, -29, -1, -27, 7, -36, 35, -13, 7, -64, 43, -36, 14, 3, -47, -47, 79, 48, 25, 31, -31, -5, 20, -55, -24, -17, 18, -44, -62, -29, 25, -13, 32, -8, -27, 4, -62, 12, 53, 36, 55, 56, -71, -59, -9, -58, -22, 59, 97, -38, -27, 7, -7, -115, 0, 19, 65, 6, -14, -36, 72, -52, -21, -53, 13, 6, 66, 57, 54, -63, -83, -35, 34, -32, 27, 25, 2, 58, 83, -53, -76, -43, -20, 21, 53, 5, -25, -19, -40, 12, 111, 64, 0, -54, -82, -90, -8, 80, 72, 3, -18, -88, -22, 89, 46, 19, 17, -1, 4, 41, -46, -36, -40, 18, 36, 66, 0, -64, 0, -7, -89, -41, 27, 35, 1, 7, 10, 66, -26, -42, 24, 48, -70, -51, 60, 68, -11, -65, -36, 10, -1, 11, 19, 40, 62, -42, -7, -24, -97, -26, 102, 2, 46, 35, -77, -25, 18, -80, 13, 62, -7, -5, 82, -39, -52, 21, -7, -38, 68, 32, -71, 25, 37, 0, -65, -14, 3, 26, -6, -35, 14, 0, -71, 13, 63, -66, 22, 82, 9, -51, -58, -56, -27, 72, 18, 32, 75, 13, -52, 2, -55, -70, 48, -17, 13, 63, 112, -36, 8, -53, -17, 28, 23, -23, -6, 9, -32, -81, -54, 37, 27, 44, 82, 20, 8, -85, -92, 12, -17, 12, 61, -41, -74, 74, 12, 17, -31, -48, 23, 74, -14, 17, 40, 42, -37, -73, -60, -11, 36, 96, 1, -37, -79, -20, 0, 38, -30, 38, -11, 44, 21, 52, -37, -36, -56, 28, 5, 26, -78, -22, 2, -1, 6, 26, -36, 31, 100, 4, -18, -10, -72, -4, 62, -30, 81, -9, -36, -47, 5, 44, 21, -79, 41, 75, -48, 35, -26, -60, -121, 13, -26, 82, 79, -18, -2, -17, -31, 5, 54, -6, 88, -21, -60, -17, 52, -93, 10, -23, 4, -6, 25, -23, 36, -69, -5, 53, -73, 43, 1, 6, 4, 32, -61, -9, -14, -9, 60, 12, 53, -28, 2, -8, 51, -54, 12, -23, 10, -10, 69, 21, 47, 6, -22, -31, 34, -49, -87, -19, 48, 85, 39, -52, -75, -86, 14, 54, 4, 0, 48, -48, -26, -23, 10, 61, 19, -46, 30, 26, -39, 47, 59, -11, 28, 18, -7, -15, -17, 12, 14, -37, 24, -55, -46, 18, 55, 14, 0, 45, -49, -70, 0, -11, -14, 49, -9, 2, 11, -26, 76, -1, -86, -17, -71, -19, 24, 31, -2, 41, -13, 55, -28, 36, 57, -11, -71, -105, -52, 79, 47, -45, 26, -2, 10, 39, -28, -57, 42, 13, 32, -60, -41, 68, 21, -41, -92, -17, 53, 127, 5, 21, -109, -20, -22, 35, 5, 43, -102, -5, 11, -30, 37, 40, 1, 55, 46, -3, -28, -37, -47, -35, 0, 96, -9, -8, -25, -10, 18, 62, 22, -15, -17, -88, 12, -11, 32, 12, 69, 5, 44, -25, -71, -28, 0, 3, -21, 22, 23, 48, 31, -9, -54, -82, -42, 57, 10, 17, 64, 82, -48, -54, -87, 51, 49, -9, -35, 9, -69, 8, 36, 17, -57, 48, 57, 56, 14, -32, -47, 11, 56, 10, 32, 28, -54, -44, -8, -77, -59, 1, -4, 24, 38, 90, 72, -100, -24, 1, 41, -8, 12, 15, 23, -62, 30, 5, 2, -29, -66, 1, 4, -38, -21, 57, -2, 3, 21, 24, -35, -14, 2, 44, 39, -45, 26, -13, -52, 1, 57, 3, -90, 0, -13, -69, 29, 97, -10, -63, 12, -15, 3, 23, 119, -27, -37, -96, -40, 6, 10, 2, 49, 42, 42, 2, -102, -24, 4, 40, -34, 35, 10, 14, -44, 18, -1, 60, 24, 28, 1, -52, -1, -43, 44, -10, -14, -83, -11, 46, 81, -73, 6, 36, -65, -15, -18, 20, 44, 38, -78, 36, 47, -35, -27, 52, 12, -39, 4, 17, 20, -38, 22, 48, 40, -35, -54, 41, 5, -23, -35, -32, 0, 73, -31, -3, 44, 3, 61, -14, -97, 0, 32, -83, -27, 75, -13, 20, 11, 9, -59, 83, -56, 24, -39, -17, 24, 86, -128, 36, 44, -53, -19, 4, -30, 91, 27, -64, -12, -61, -17, 53, 34, -7, 66, 0, 5, -9, 32, 17, 20, -58, -42, -43, -19, 10, 0, -45, 51, 105, 0, -37, -32, -20, -8, 102, 37, -51, -32, -57, 0, 30, 34, -47, -65, -57, 89, 70, -1, 49, 12, -30, 41, 18, -73, -58, -57, -73, 65, 31, 27, 25, -25, 10, 11, -47, 66, 39, -65, 10, -24, -59, 32, -4, 59, 13, 8, -46, 0, -4, 1, -73, -7, 15, 22, -3, 46, 21, -40, -51, 25, 55, 39, -35, -79, -3, 35, 65, 39, -56, -75, 36, -38, -26, 104, -22, -28, 0, -62, 37, 75, -107, 61, 7, -76, 68, 29, -95, 39, 39, -97, 24, -29, 6, 53, 48, -40, 21, 23, -4, 13, -60, 17, -11, 40, -89, 37, -37, 20, 10, 21, -19, 24, -58, 0, -12, -26, 14, -4, 29, 29, -58, -9, 29, 15, 12, -25, -7, 74, -38, 5, 18, -46, -51, 75, -8, -32, 29, -51, -42, 23, -21, 47, 62, -55, -15, -1, -42, 19, 99, 4, 27, -25, 10, -31, 0, -125, 20, 37, 1, -18, 102, 25, -96, -11, 6, 28, -11, -53, 11, 27, -59, -29, 11, -43, 20, 0, -5, 86, 74, -46, -58, 82, 23, -8, 5, 1, -43, 20, 37, -45, 14, 26, 0, -48, -38, 21, 103, 1, -10, 28, -110, -35, 127, 75, 8, -59, -42, -1, 44, 60, -29, -36, 47, -6, -94, 57, 31, -55, 24, 38, -77, -30, 37, -8, -10, 40, 0, -29, 9, 55, -76, -36, 80, 40, -4, 24, -36, -57, -20, 29, 69, 26, -83, 61, 27, -85, -57, 32, -39, 12, -34, 57, 28, 54, -30, 78, -35, 41, -4, -73, -78, 120, -21, -15, 46, 35, -15, 6, -27, 13, -72, -52, -29, 36, 47, 0, -12, 0, -3, -17, -9, -19, 18, -38, 2, 63, 27, 41, -59, -23, -48, -27, 5, 57, -22, 66, 18, -19, -63, -14, 43, 66, -52, 29, 34, -72, -20, 13, 25, 30, 0, -59, -47, 40, 26, 6, 27, 82, -82, 17, -3, 39, 37, 12, -77, -27, -59, 2, 105, -39, -17, 36, 48, 56, 17, -128, -6, 31, -68, -2, 23, 14, 4, 79, -6, -40, -115, 26, -21, 46, 1, -3, 25, 63, 66, 22, -73, -21, -3, -9, -10, -54, -37, 110, 57, -25, -51, -57, 46, 9, 80, -10, -36, -113, 18, 74, 21, -45, 63, 49, -74, -3, -7, 21, -54, 40, 27, -19, -68, -41, -12, 39, 11, 28, 41, -55, 3, 57, -74, 23, 41, -60, -89, -38, 14, 72, 94, -38, 1, -21, 39, -46, -27, -42, 27, 70, -10, -39, 9, 18, -61, 21, 66, 89, 15, -119, -13, -7, -56, -12, 49, 42, 98, -53, -8, -9, -79, -66, 76, -25, 3, -3, 32, -25, 42, 61, 57, -24, -27, -88, -86, 54, 47, 68, 32, -19, -24, 19, 42, 22, -87, -106, 3, 15, 28, 93, 18, -128, -37, 8, 37, 0, -47, -55, 43, 60, 23, 2, 0, 26, -127, 8, 0, 3, 55, 38, 9, 2, -52, -51, 42, 2, 3, -49, -13, -37, 27, 25, -35, 12, 42, -9, 34, -18, -86, 0, 35, 31, 30, 9, -11, 5, 25, -24, -30, 14, 26, 14, 80, 39, -55, -3, -14, -44, -8, 32, 5, -28, -32, 92, 3, -96, -25, 64, 43, 3, 31, -4, 3, -87, -8, 29, 26, -77, 68, -31, -23, -6, 0, 14, 41, -44, 34, 2, -65, -12, -18, 23, 21, -20, 38, 26, -93, 7, 79, -9, 15, 31, -82, -18, 9, -21, -30, 64, -62, 54, -32, -6, -26, -23, 7, 77, -80, -9, 96, 30, -29, 27, -2, 29, -9, 0, -37, -37, -15, 46, -24, 20, 7, -26, -41, 52, -47, 29, 2, 14, 20, 66, 32, 0, -75, -35, 42, -30, -22, 43, -24, -29, -76, -10, 34, 41, -24, 64, 43, -54, -34, -31, -61, 11, 53, -5, 47, 42, -21, -59, -17, -6, 96, -3, -24, 18, 42, -70, 21, 26, 1, -45, -36, 22, -12, -8, 32, 22, -46, 46, -15, 11, 9, 10, 3, -32, 6, 0, 31, -54, 31, -19, -53, -47, -31, -26, 90, 44, -58, 44, 20, -74, 14, 46, -2, 9, -46, -11, -1, -45, 61, 52, -49, -24, 70, 23, 1, -51, -28, -63, 24, -2, 26, 65, 87, -55, -19, 26, 23, -45, 64, 1, -5, -25, -38, -32, 18, -9, 56, 20, 19, 28, -38, -65, -22, -3, 22, 114, -30, -21, -21, 36, 30, -1, -73, 56, -9, -8, -5, -59, 28, 13, -110, 43, 32, -86, 27, 15, -65, -75, 60, 59, 20, -83, 18, 48, 95, 39, 3, -58, -71, -71, 39, 70, -7, 9, 8, -25, -20, 25, 90, -36, -38, 25, 1, -76, 61, -18, -17, -46, 52, -10, -57, -36, 107, 27, 4, 29, -38, -14, -34, -51, -94, 36, 27, 57, -46, 29, 3, 26, 83, 48, -128, 29, 4, -75, -21, 21, -23, 54, 73, -9, 41, 24, -80, -68, 32, 45, 20, 21, -51, -73, -13, 39, 8, 3, 100, 7, -48, -98, -43, -5, 53, 7, 11, -39, 27, 39, -13, -40, 59, -63, 1, 75, -4, -17, -11, -13, 24, 103, -5, -45, -66, 0, 17, -4, 3, 72, -5, -42, -40, -14, 17, -2, 28, 32, 0, -3, 13, -128, 10, 39, 105, 65, -12, -82, 19, 12, -29, -27, -27, -42, 58, 10, 2, -106, 9, 45, 72, 59, -8, -107, 23, 35, 11, 39, -49, -41, 47, 28, 15, 18, -81, -128, -29, 100, -23, 2, 77, 19, -128, 20, 21, 25, 22, 96, -57, -78, -77, -36, -18, 48, 75, 22, -46, -26, 75, -2, 10, 2, 19, -56, 32, 41, 0, -12, -30, -44, 8, 69, 63, 24, -104, -69, 17, 53, 1, -85, -57, 5, 14, 107, 5, -63, 22, 15, -39, -47, -40, -36, 48, 39, 54, -55, -14, -94, -18, 79, 91, 44, 8, -63, -47, 44, 39, -15, -36, -36, 7, -56, 52, 0, -10, 42, 87, 38, 18, -103, -64, 94, 14, -49, -58, 59, 32, 8, -57, -25, -34, 48, 81, 25, -35, -27, 21, 35, 43, -19, -61, 28, -29, -2, -4, -2, -35, 39, -90, 18, 102, 37, -53, -47, 13, 75, 27, -31, -74, -4, 42, -20, -46, 12, 62, 35, 54, -47, -36, -7, 29, -28, 45, -1, 18, 3, 9, -95, -42, 9, 66, -37, 26, -26, -36, -82, 65, 15, -56, -39, 56, 52, 58, 54, -21, -56, -58, -65, -94, 32, 111, 29, 38, 38, -20, -128, 9, -45, 0, 104, 38, -26, -1, -22, -55, 3, -78, 24, 74, 28, 78, 0, -22, 23, -41, -46, 29, -29, -53, 32, -63, 48, 37, 54, -7, 0, -89, -23, 47, 107, 57, -52, 1, -38, -23, -12, -3, -7, 76, -65, -29, 79, 15, 80, -18, -89, -14, 10, -24, 0, 15, -26, -42, -19, 34, 24, 24, 13, 27, 20, -32, 9, -3, 7, -38, -44, -19, -44, -90, 5, 104, 1, 47, 10, -30, -21, 56, -90, 28, 63, 9, -31, -30, 20, -40, 28, 2, -55, -52, 76, 58, 77, -10, -20, -45, -43, 0, 23, -46, -40, 21, -22, 13, 100, 34, -66, 19, -28, -43, 65, 47, -15, 22, -27, -8, -38, -12, -44, 2, -40, 77, 18, 14, 54, 10, -10, 82, -9, -60, -83, 8, 27, 35, 31, -7, -109, -13, -32, -5, 94, 79, 14, 36, -98, -34, 9, -56, -19, 99, 69, -25, 28, -43, -69, -28, 19, -34, 47, -28, -75, 63, 69, -7, -37, 14, 38, -48, 6, 51, 39, -34, 29, -15, -41, 5, -26, -30, -36, 45, 32, 8, -80, -9, -45, -21, 11, 59, 104, 19, -71, -2, -21, 26, 20, 2, 1, 45, -63, -11, 68, 42, 5, -100, -18, -1, 26, 53, 48, -64, -8, -35, -11, 54, 17, -72, 2, 10, -31, -78, 6, 53, 52, -7, 45, 20, 20, -27, 6, -34, -35, -47, -27, 2, 121, 55, 20, -58, -47, 61, 9, -71, 44, -20, -35, 31, 43, -20, 0, 0, 13, -3, 0, -11, 7, 12, -93, -38, 37, -44, -45, -26, 8, -42, 46, -2, 53, 29, 57, 13, -34, -98, -60, 28, -22, 34, 60, 29, 3, 0, -2, 0, 10, -70, -63, -37, 12, 47, 70, -71, -53, 85, -36, -76, 43, 83, -25, -58, -103, 5, 74, 48, 12, -47, -36, -64, 0, 22, 114, 57, 14, -70, -105, -60, 10, 5, 42, 15, -46, 48, 63, -91, 25, 94, -25, 4, 0, 2, -32, 40, -20, -1, 27, 56, -128, -4, 29, -94, -18, 85, 7, -49, 5, 18, 32, 38, 5, -19, -23, -18, -22, 21, 25, 2, -65, -37, 32, -41, -32, 71, -4, 5, -2, -1, 42, 12, -10, 58, 52, 15, -37, -89, -94, 18, 22, 37, -1, 3, -74, 27, 43, 24, 4, 35, -12, 42, -45, -10, -26, -43, -46, -5, -47, 53, 121, -15, -11, -22, -8, -48, -9, -19, 54, -4, -11, 0, 54, 61, -3, -79, -30, -31, -56, 70, 32, 22, 59, -41, -114, 58, -32, 1, 2, 9, -57, 95, -37, -46, 15, 27, -38, -19, 27, 29, 55, 6, 49, -29, -116, -23, 64, 6, 40, -19, 18, -48, 20, -71, 1, -42, 127, -9, 22, -25, -22, -46, 53, 13, 63, -12, -95, -29, 73, 15, 15, -13, -13, 47, 26, -91, -94, 17, -3, 76, -13, 14, -92, -1, 46, 94, -23, -43, -35, -44, -18, 105, 32, 5, -8, -55, -77, 104, 47, -12, 15, -30, 27, -6, 55, -25, -27, -60, 88, 1, -65, 17, 51, -31, -22, 62, 28, 30, -69, -43, 17, 9, 23, 42, -18, -74, -30, -24, 65, -7, -35, -58, 57, 58, 47, 46, 11, 2, -34, -68, -69, 48, -20, -60, -25, 73, 68, 32, -57, -91, -9, 81, 53, 1, 46, -18, -87, -13, 11, -35, 10, -23, -58, 44, 42, 19, 55, 2, -34, 53, -27, -100, -66, 56, -22, 18, 20, 26, -75, -19, -85, 62, 34, -14, 21, 127, -28, -59, -83, -9, -26, 23, -21, 35, 106, 25, -56, 32, -34, -36, 77, 0, -70, -28, 8, 59, 19, -3, 28, 0, -57, 7, -19, -41, 9, 13, -55, 39, 89, 45, 7, -45, -103, 38, 40, 15, -4, 34, 0, 24, -69, 37, 17, 12, 30, 14, -26, 75, -43, -109, -55, 7, 53, 116, -27, -76, 0, 46, 21, -3, -73, -91, 2, 20, 37, 52, 96, -81, -36, -22, 34, -41, 7, 17, 73, 1, -43, -62, -61, 28, 4, 11, -36, 86, 10, -43, 17, -2, -41, 17, 11, -59, -31, 31, 12, 55, 19, 14, -31, 40, 59, -22, -107, -58, 2, 12, 77, 13, -41, -57, 10, 7, -62, -22, 82, -7, 45, 63, 13, -51, -94, -64, 78, 27, 22, 20, -55, -82, 32, 19, 24, 68, 2, -106, -14, -31, 19, -2, -23, 32, 52, -53, 81, 68, -111, -45, 6, 15, 15, -31, -28, 56, 61, 35, -49, -17, -3, -25, -117, 48, -44, 34, 76, 68, -5, 80, -46, -76, -65, 11, 8, 6, 6, 12, 39, -7, -39, -31, 37, 54, 55, -65, -72, -52, 10, 62, 4, -6, 58, -43, 0, 13, 45, -46, 30, -21, 37, -9, -6, -10, -27, -71, 23, 40, -94, -18, 58, 66, 63, -26, -29, -45, -35, 49, 35, -30, -64, 12, -18, -19, -35, 89, -19, -1, 10, 34, 5, 31, -22, -87, 25, 25, -10, 7, -11, -83, 106, 40, -96, 22, 53, -66, -18, 88, -18, -40, 57, 18, -42, 34, 57, -27, -56, -36, -43, 35, 22, 59, 27, 56, -12, 23, -30, -62, -107, 0, 42, 2, 8, 48, -4, -61, 39, 26, -21, -6, -10, -115, -54, 110, 36, -6, -17, -56, -36, 59, 92, 19, 8, -3, 6, 20, 11, -108, -17, -29, -28, 81, 73, -37, 3, -48, -74, 61, -18, 4, 36, 82, -66, -14, -104, -18, 46, 53, 10, 65, -14, -94, -58, -32, -28, 58, 123, 75, -42, -78, -8, -1, -12, 2, 95, -43, -6, 88, -20, -62, 56, 56, -94, -20, 22, 17, -51, 52, -4, -10, -29, -70, -22, 74, 42, 3, 57, -46, -29, -7, 30, -19, 15, -100, 29, 22, 8, -49, 43, -27, 85, -20, 7, -35, 37, -44, -21, 40, 37, -46, -40, -32, -27, -41, 60, 37, 48, 34, -7, -95, 104, 25, -85, 39, 4, -76, -32, 4, -18, 69, 57, -3, -25, 2, 85, 10, -52, -11, 94, -43, -18, 17, -55, -8, 59, -18, -59, 42, 7, 44, 22, 9, 0, 9, -85, -18, -38, -14, 24, 59, -108, 56, -36, -15, 85, 23, -90, 47, 25, -19, -43, -8, 61, -10, -17, 6, -85, -87, 77, 5, 42, 40, 45, -71, 35, 23, 18, -40, -31, -61, -27, -18, 2, 46, 55, 57, 88, -22, -75, -70, 14, 15, 72, 0, -21, -19, 38, -18, -51, 44, -23, -11, 34, 7, -60, -9, -30, 60, 21, 20, 35, 2, -36, -7, 7, 53, -63, -52, -5, 62, -3, -83, 4, 11, 7, -10, 31, -34, 5, -70, 63, 1, 29, -10, -48, -90, -14, 44, 89, 39, -46, 37, 5, 0, 34, 25, -119, -30, 56, 45, 18, 49, 12, -115, -44, 79, -7, -4, 69, -11, -37, -57, -11, -46, 35, 25, 5, -31, 22, 11, 23, -44, -74, 21, 40, 3, 20, -39, 38, -34, 26, 5, 85, -71, 2, 32, -18, -107, 13, 32, -64, -2, 44, 64, -47, -7, -15, 71, 26, 34, -89, 29, -58, -14, 44, 30, -30, 43, -98, -66, 44, -28, 22, 38, -14, -3, 34, -2, -38, 5, 29, -10, 29, 74, 20, -27, -19, -64, 55, 10, -26, -80, 35, -6, 36, 34, 10, -12, 0, -29, 40, 15, -79, 0, 4, -62, 45, 59, -21, -55, 5, 30, -18, -11, 28, 98, -29, -6, -13, 6, -28, 5, -70, -3, 27, 14, -32, -25, -8, 30, 79, 97, -4, 15, -40, -13, -40, -68, -18, -20, 2, 48, 98, 37, -11, -8, -6, -117, -41, 69, 54, 28, -37, -52, 20, 25, 19, 19, -103, 24, 0, 11, -49, 19, -91, 27, 57, 7, 46, 82, -102, -32, 42, -40, 36, 64, 9, 34, -10, -44, -19, -70, -54, 39, 65, 4, -30, -65, 17, 39, -10, -46, 6, 3, 69, 23, -64, 20, -1, -40, 54, 73, -20, -35, 41, 0, 9, 65, 15, -95, -82, -81, 5, -10, 22, 120, 38, -100, 46, -18, -72, 39, 44, -39, -69, -7, 100, 65, -47, -24, 19, 25, -35, -4, -56, 21, 18, 9, -47, 70, -38, 20, 14, -3, 8, 25, -1, 5, -63, -5, 88, 21, -15, 79, -45, -11, -30, 37, -78, 4, 37, 53, -39, 9, -73, -21, 41, 30, 83, 23, -73, 44, 28, -48, -18, -85, -10, 63, 44, -71, 39, -52, -1, 19, 79, -80, -10, 26, 4, -96, 36, 59, -45, -30, 39, -21, 42, -3, -12, 30, 11, 29, 23, -43, -9, 42, -32, 2, -13, -74, 10, 66, 7, -43, -13, -27, 8, -43, 42, 47, 32, -47, -40, -1, 37, 56, 29, -29, -45, -19, -30, 18, 75, -11, 70, -17, -17, -76, -55, 1, 59, 61, 12, 12, -81, 17, -30, 29, 13, 1, -21, -21, -47, 43, 105, -49, -19, -92, -42, 98, 60, -10, 21, 36, -45, 1, -46, -37, -35, 91, -35, 3, -28, 9, -22, 15, -61, 54, -10, 20, 2, -37, 12, 38, 91, -9, 13, -76, -10, 4, 65, -44, 43, -1, -66, -47, 14, 57, 20, -13, 71, 26, -93, 5, 36, -27, 0, 24, 51, 44, -42, -75, 25, 31, 96, 30, -82, -48, -2, 2, -48, 43, 25, -8, -73, 113, -22, -4, 34, -22, -90, 76, -46, -35, 64, 95, -63, 0, -30, -39, -66, 81, 31, -51, -38, 27, -62, 43, 51, 19, 15, 94, -11, -37, -64, -85, -29, 36, 46, -17, 43, 9, 3, -13, 73, 14, 17, 17, -78, -27, 26, -6, 28, 0, -72, -82, -49, 24, 47, 56, 86, -26, -104, 43, 75, -22, -41, -80, 0, -29, 46, 22, 100, -53, 26, -39, 1, -12, 106, -6, -17, -39, -29, 34, 3, -25, -55, 14, -47, -28, 55, 81, -6, -70, 1, 28, 45, -8, 99, -51, -30, -74, -31, -1, 127, 12, -5, -19, -6, -57, -34, 5, -56, -28, 96, 0, -11, -13, 19, -14, 81, -55, -6, 48, 43, -48, -51, 15, -36, 27, -11, 75, -36, 53, 42, 24, -60, 53, -48, -63, 0, 46, -41, -5, -26, -39, -71, 24, 119, 29, -39, 74, -10, -59, -31, 82, -6, -56, -26, 92, 12, 41, 76, -72, -78, 59, -5, -128, 8, 90, -26, -5, -37, -8, 5, -6, -42, 124, 21, -91, -4, 64, -12, -62, 34, -40, 19, 23, 49, 5, 23, -103, 19, 72, 46, -41, -26, 26, 15, -7, 13, -25, -57, 39, 45, 32, 62, -64, -86, -5, -17, -85, 60, 13, -54, 20, 47, -20, 61, 24, -47, -10, -12, 18, 0, -68, -27, 85, 17, 8, -13, -6, 42, 45, -70, 0, 20, 35, 26, -56, -51, 62, -44, 5, -22, -38, 23, 99, 7, -2, 15, -43, 35, 4, -30, -44, -17, -75, -12, 20, 59, 72, 7, 52, -44, -15, -46, -54, -83, 72, 69, 18, 6, -57, -34, 60, 24, 27, -6, 9, -43, -38, -64, 75, -8, 66, 40, -71, 1, -3, 38, 39, -44, -106, 23, 9, 70, 52, -23, -116, -28, 120, 26, 15, 0, -23, -17, -4, -36, 4, 13, 31, 3, -14, 57, 6, -58, -17, -40, -26, 56, 52, -8, -35, -12, -59, -24, 74, 34, -31, 26, 82, -64, -7, 5, -17, -7, 38, 3, 42, -46, -11, -47, 5, -92, 41, 48, 74, -108, 5, 13, 73, 21, 42, -90, -26, -13, 5, 37, 25, -71, 10, 10, -3, 57, -69, -29, 40, 0, 11, -41, -11, 13, -20, -45, 77, -36, 30, 48, 17, -31, 44, -51, -65, 7, -41, 10, 122, -28, -4, 0, -68, -13, 75, -38, 21, 3, -93, 12, 114, -5, 2, 2, -49, -51, -1, -19, -36, 75, -5, 15, -71, 51, -41, 42, -35, 1, -20, 109, 6, 26, 54, -12, -59, 37, -13, -96, -4, 55, -41, 6, 14, -97, -23, 35, -44, 25, 87, 19, 34, -44, -23, 4, -24, -61, -15, -39, 124, 64, 13, 3, -17, -19, -34, -21, 42, 35, 4, 6, -20, 39, -32, -80, -52, -6, 4, -21, 6, 31, 76, -47, -6, -32, -13, -44, 22, -20, 12, 66, 78, -1, -115, -43, 63, 54, -24, -42, -72, -25, 88, 21, 29, 53, -12, -58, 9, 41, 31, -55, -64, 75, 22, -30, 1, -42, -21, 44, 52, -46, -47, -58, 97, 22, 61, 4, -29, 0, 11, -103, 46, 48, -18, 2, -4, -15, -22, -69, 21, 71, -6, -19, 6, -46, 22, 28, -32, 10, 127, 29, -51, -9, 47, -64, -14, 83, 22, 0, 75, 0, -89, -24, 40, -10, 10, -51, -27, 37, 7, -24, -40, 0, -32, -26, -11, 82, -4, 12, -5, 2, 35, 12, -27, -12, -47, 39, 25, 59, -43, 12, 4, -25, -114, 34, 19, -41, -13, 21, 10, 76, 15, -35, 5, -12, 20, 86, -65, -36, -9, -19, 65, -3, -29, 35, -2, -63, 1, 0, 53, 45, -56, 26, -66, 9, 21, 0, -105, 92, 20, -7, -52, -2, -29, 46, 54, 69, -113, -38, 31, 44, 36, 43, -75, -99, -7, -51, -13, 63, 89, 49, 21, -42, -56, -78, -27, 8, -23, 15, 104, 47, 60, -30, -39, -10, 61, -70, -46, 23, 64, -19, 53, -60, -14, 7, -49, -76, -3, -15, -4, 34, 27, 108, 6, -41, -25, 36, -27, -6, 1, 34, -42, -42, 27, 28, 15, -18, -37, -73, 8, -15, 18, 22, 88, -30, -19, -57, -79, 23, 79, -17, 63, -42, -42, 39, 39, -82, -24, -51, 7, 48, 25, 51, 56, -12, -89, 12, -4, -32, -58, 83, 28, -57, 29, 80, -32, -52, 34, 0, 49, 0, 3, 30, 4, -88, -46, 30, 11, 94, -19, -18, 9, -24, -102, 24, 3, -47, -8, 78, 18, 3, 58, -28, -44, -53, 26, 26, 99, -70, 42, -57, 0, -2, 104, -78, -4, -7, 2, 25, 46, 0, -31, 6, -49, -75, -14, -17, 17, 11, 12, 15, 124, -34, -56, -52, 8, 24, 93, -12, -4, -44, -48, -45, 127, -11, -10, -49, 17, -21, 105, 10, -2, -27, -79, -57, 93, 29, -69, 30, 2, -54, -38, 93, 18, -22, 11, 9, -100, 40, 32, 7, -2, 75, -15, 41, -54, -51, -7, 80, 35, -25, -91, -28, 15, 73, 24, -14, -42, 23, -39, 41, -71, -20, 46, 79, -56, -25, -49, 39, 10, 20, -1, -5, -9, 89, -35, -17, -18, -63, -53, 26, 21, 62, -17, -44, 63, 0, -7, 47, 61, -53, -41, -103, -29, 1, 40, -7, 111, -29, -8, 47, 55, -85, -29, -61, -44, 12, 38, 97, 46, 5, -65, 1, -20, 31, -20, 34, 4, -39, -40, 53, 18, -6, -22, -79, 0, 69, -27, 48, 7, -121, -76, 127, 0, -41, -48, -13, 32, 45, -63, 19, 51, -4, 27, -18, 11, -26, 46, 19, -14, -68, 75, -7, 17, 36, -42, -38, 6, 9, 2, 20, 91, -27, -32, 25, -6, -96, 24, -31, -56, 3, 94, -8, 37, -57, -5, -5, -1, -41, 103, -31, -32, -38, 34, -23, 24, -76, 17, 57, 73, -59, 51, 3, -77, -57, -48, 8, 10, 40, 51, -4, -25, 52, 0, 55, 9, -11, -38, 0, 31, 31, -35, 43, -64, -70, 4, 53, 30, -47, -43, 2, 0, 62, 64, -78, -20, 35, 31, -4, 83, -51, -55, 20, -55, -86, 44, 95, 10, -83, -60, 65, -2, -26, 20, 75, -25, 7, -56, -10, 0, 8, -83, 36, 61, 0, -12, 39, 1, -49, -60, 0, 48, 107, 9, 20, -45, -93, 6, 30, -51, 31, 45, -18, -47, 27, 21, 86, -66, 36, -74, 26, 13, 14, -120, 80, -1, 41, -15, 9, -1, 95, -66, -13, 5, 28, -51, 3, 35, -26, -7, -10, -94, 10, 85, -51, -32, 56, 24, 23, 78, -58, -39, -11, 32, -39, 75, -9, -43, -71, -25, 20, 38, -41, -20, 27, 68, 1, 36, -51, 7, -99, 75, -31, 14, 2, 83, -19, 20, 14, -41, -74, 38, 49, -24, 9, -11, -99, 17, -4, 37, 35, 52, -88, -40, 7, 29, 65, -2, 22, 28, 25, -117, -5, 8, -53, -8, 73, -13, 27, 44, 38, -41, 3, -126, 11, 74, 59, -34, -29, 0, -39, 75, -32, -5, 7, 106, -72, -34, -51, -51, 15, 13, 8, 102, 31, 12, 45, -80, -82, 62, 14, -41, -26, 18, 78, -12, -35, 42, -38, 20, 26, -20, -107, -7, -32, 92, 38, -32, -27, 55, -2, -14, -9, -52, 30, 40, 37, -8, 35, 8, 38, 19, -42, -64, 19, 41, 2, 35, -25, -12, 35, -39, -46, -95, -43, 35, 17, 5, 34, -25, -28, 63, 59, 58, 38, -46, -53, -35, 27, -22, 14, -32, 44, -60, 68, -57, 4, -90, 3, -48, 113, -36, 28, -5, 59, -31, -14, -45, 51, 24, 27, -38, -93, 22, -2, -12, 51, 54, -63, 13, 30, 1, 34, 35, -62, -82, -47, 20, 18, 66, 68, -22, 5, 31, -106, -32, 58, -6, 48, 93, -69, -35, -82, -43, 34, 105, -47, 48, 20, -53, -14, 27, -98, -2, 96, 13, -3, 29, 41, -48, -77, -93, 7, -6, 58, 87, 68, -97, -39, 40, -5, -76, 35, 2, -79, 7, 34, -85, -10, 116, 1, 19, 77, -9, -46, -14, -19, 17, 43, -54, -43, -24, 58, 9, 23, -34, 31, -36, 42, 13, 5, -85, -66, 13, 82, 9, -70, -6, -27, 35, 71, 66, -24, -77, 6, 2, -31, 25, 21, -14, 47, 17, -86, 26, -27, -17, -41, 105, -48, 5, -46, 29, -38, 2, -29, 49, -29, -20, 0, 62, 66, -7, 5, 78, 8, -75, -5, -51, -74, 74, 0, -3, 26, 25, -97, 38, 49, 74, -44, -28, -75, -7, -28, 42, 31, 59, 71, 14, -54, 24, 29, -51, -53, -79, 3, 2, 46, 38, 35, -47, 9, -63, 60, -23, -8, -79, 74, 14, 15, -35, -36, -37, 60, -21, 12, 89, -26, -93, 4, 5, 3, -25, -11, 61, 86, 24, 7, -4, -13, -41, -44, -66, 86, 27, -31, 75, -1, -40, 9, -17, -96, -9, -19, 82, 19, 68, 9, -44, 8, 77, -12, -26, -37, 36, -11, -19, -17, -7, -43, 22, 38, 65, -46, -42, -12, -71, 7, 70, 19, 0, 10, -48, -24, 17, 46, 30, -6, -30, -65, -30, 60, 19, -19, 46, -51, -46, 75, 31, 1, 9, -32, -46, -46, -59, -8, -12, 7, 94, 7, 29, 46, 20, -73, 41, 24, -21, -24, -38, -36, -34, -44, -2, 64, 25, 44, 5, -96, -55, 70, 93, -2, -45, 38, 6, -76, -29, 12, -63, 89, 57, -21, -5, -17, -20, 51, 34, -26, 34, -32, -21, -36, -4, 11, -39, 51, 41, -51, -81, 52, 47, 78, 36, -36, -64, 10, 32, -24, 3, 49, -21, -89, -41, 18, -39, 22, 93, -12, -39, -22, -47, -45, 0, -13, 20, 86, 26, 26, 37, 37, -58, -64, 22, -37, 6, -10, -41, 0, 35, -10, 36, 41, -60, -10, -53, 26, -27, 9, 40, 2, -41, 72, 38, -36, -23, -44, 21, 63, -7, -60, 72, -61, -19, 73, 58, 52, -6, -43, -22, -15, -62, -35, 6, 43, -20, 5, 66, -21, -18, 46, 52, -9, -51, -51, 3, 45, 24, -1, 96, -15, -37, -62, -41, -22, 54, -41, 10, -21, 41, 83, 30, -80, -8, 51, 0, -15, -3, 40, -23, -29, -63, 20, 38, 57, -32, 38, 18, -7, -4, 26, -22, -62, 9, 54, 1, -122, -23, 65, -22, -55, 10, -2, 41, 65, -2, -58, 19, -60, -20, 51, 58, 25, 74, -78, -20, -23, -37, -57, 37, -27, -26, -8, 10, -14, 62, 56, -91, 19, 69, -3, -3, 74, -32, -24, -36, -58, -29, 96, 55, 13, -14, -57, 2, -58, -8, 47, 58, 41, -23, -58, -48, -19, -13, 87, -29, -8, 30, 44, -7, -65, -86, 29, -47, -29, 127, 10, -37, 44, -9, -14, 49, -70, -88, 30, 6, 4, -36, -12, 0, 45, 27, 1, -13, -20, 46, 94, 34, -86, -18, -13, -74, 11, 75, -41, 43, 31, -17, 31, 28, -55, 52, -30, -78, 48, 21, -51, 42, 56, 8, 15, 1, -24, 15, -54, -51, -59, 41, -17, -4, -46, 106, -22, 23, -32, -45, -51, -12, 36, 91, 7, -19, 32, -29, 42, 63, -74, -56, 73, -32, 1, -42, 26, -63, 15, 27, 31, -65, 93, 0, -110, -30, 24, -6, 68, -19, 6, 29, 27, -54, 36, 17, -80, 25, 8, -61, -59, 6, 35, 27, 32, -27, -11, -5, 31, -15, -7, 58, -5, -11, -60, 23, -54, -6, 72, 96, -72, 2, 19, -43, -3, -3, -10, 54, 2, -48, -13, -45, -18, 41, -46, 15, 49, 51, -32, 22, -38, -35, 0, 53, 25, 87, -44, 29, -59, -52, 0, 62, -48, 47, 44, 0, -88, -86, 17, -12, 19, -36, 9, 25, 52, -12, -2, -28, -11, 52, 36, -32, -35, -13, -28, -72, 8, -40, 2, 34, 56, -36, -11, -39, 12, 59, 66, 43, 10, -14, 9, -56, -46, 7, 0, 41, 37, -20, -27, 47, 0, -40, -59, -34, -43, 81, 83, 22, -24, -49, 47, 59, -14, -63, -42, -52, 30, 124, 55, -47, -32, 23, -37, 41, 58, -4, 40, -30, -19, -19, -31, -34, 109, -76, -13, 0, -12, -39, 73, 54, -5, -99, -1, 40, -51, -5, 38, -70, -26, 90, 12, -83, 4, 40, 19, 28, 62, -66, -11, 5, -64, -22, 0, 5, 48, -2, -49, 21, -71, 48, 99, -34, 14, -13, -15, 25, 7, -79, 51, 7, -70, 19, -15, 15, -21, 45, -17, 19, -26, 29, 25, -24, 20, -6, -1, -19, 42, -15, 17, 19, -5, 11, -23, -23, -14, -41, 14, 6, 73, 37, 32, -82, 14, -74, 31, 27, -3, -59, -20, 30, 59, 32, 31, 73, -90, 3, -6, 42, -57, 0, -31, -28, -5, 115, 38, -25, -64, 14, -29, -39, 72, 40, -87, -8, -3, -29, 70, 94, -42, -20, 0, 9, -78, 23, -11, -8, -46, -43, 1, 44, 72, -36, 45, 35, 25, -73, -22, -1, 17, -47, 36, 104, -15, 18, -18, -45, -35, 55, -64, 34, -39, -44, 17, 66, 78, 37, -128, -39, 35, 38, 44, 59, -80, -61, 32, 0, -4, -18, -35, -40, 77, 10, 44, 31, -68, -40, -9, -53, 40, 61, -63, -29, 13, -43, 40, 85, 39, 63, -54, -40, -46, 20, 31, 53, 0, 1, -49, -61, -51, -70, 58, 66, 2, -8, 13, -43, -12, 1, -49, 21, 77, 60, 4, 13, 14, -53, 20, -30, -34, -42, -26, 6, 59, -18, 49, 71, -72, -47, 55, -49, -3, 45, -2, -37, 46, 22, 42, -26, -66, 52, 12, -107, 3, 36, 56, -3, -56, -49, -34, 42, 28, 48, -21, -56, -35, 52, -24, 79, 48, -43, -68, 48, 5, -4, -89, 12, 34, 78, 59, -23, -6, 26, 29, -65, -22, -109, -3, 44, 80, 13, 61, -62, -4, -15, -52, -45, 124, 13, -51, -8, 43, -11, -2, -18, 3, 19, -10, 15, -28, -1, 14, 2, -12, -18, 30, -34, 38, -6, 58, -2, 25, -88, 3, 47, -83, -26, 71, 81, -13, 22, -66, -60, -15, 99, 9, 27, -19, -51, -40, -11, 12, 24, -3, -69, -36, 15, -56, 46, 75, 14, 48, 11, -29, -37, 17, 5, 9, -20, 4, 22, -27, -34, -58, 82, -26, 41, 43, -13, -91, -21, -28, 31, 66, -18, -15, 8, 38, -20, -30, -28, -21, -44, 34, 34, 37, 49, -83, -42, 25, -47, -62, 51, 66, 10, 65, -7, -42, 19, -30, -48, 60, -17, 9, 19, -62, -68, 74, -21, 6, 48, 0, -112, -38, 21, 14, 69, 8, 0, -51, -60, -42, 26, -62, -6, 99, 53, -7, 19, -35, -27, 62, 3, -79, -6, 46, 45, -42, -11, 2, -10, -25, 8, -6, 54, 71, -19, -93, -13, 121, 29, -89, -20, -8, 55, 31, -43, -27, 27, -66, 38, 107, 18, -61, -73, 31, 46, -14, 23, 40, 10, -28, -76, -15, 24, 26, 0, 4, 39, 8, -77, 15, 5, -24, 53, 19, -45, -45, -47, 10, 53, 18, -10, 4, -73, 1, 28, -64, -37, 43, 32, 25, -10, -26, -25, -39, 57, 99, 13, -28, -83, 43, -20, 13, -37, -37, -14, 127, -23, -19, -34, -75, 12, 81, -3, -29, -49, -11, 17, -6, 52, 31, -51, 23, 86, -66, -10, 17, 65, -8, 47, -5, -3, -96, -39, 34, 48, -58, -48, -41, -15, 1, 60, -20, 1, 65, 38, -52, 22, -15, 1, 0, -17, 31, -21, -24, 9, -63, -68, 77, 52, 0, 8, -46, 57, -60, -8, 14, -6, -31, 0, 0, 39, 2, -32, -6, -85, 42, 45, -8, 45, 42, -38, 8, -61, 0, -20, -22, 56, 58, -100, 30, 10, -43, -63, 40, -39, 24, 19, 46, -43, 103, 24, -48, -108, 34, 71, 49, 29, 12, -53, -98, 72, 4, -35, -51, 17, -30, 35, 68, 57, -41, -69, 51, 14, -39, -59, 45, 52, -35, 13, -12, -36, 53, 75, -10, 43, -80, -60, 31, -32, -44, 72, 38, -35, -12, -43, -6, 31, 90, -3, 27, -44, 63, -21, -71, -41, -35, -10, -28, 38, 39, 41, -28, 112, 12, -97, -35, -36, -24, -34, 52, -8, 95, -8, 48, -34, 0, -41, 31, -27, -7, -1, -46, 22, 48, 19, -86, 31, 57, 27, -15, -9, -24, -38, -19, -5, -6, 52, 52, -11, -35, 65, -35, 35, -1, -72, -65, 99, 31, -6, 13, 25, 44, 8, 17, -46, -99, -98, 28, 36, 127, 26, -109, -57, 47, -31, 13, 60, 7, 44, 31, -102, -86, 66, -38, -37, 63, 76, -83, -8, -54, 21, 30, -30, -8, 39, -43, -45, 77, -31, 51, -18, 12, 34, 53, -128, -14, 65, -45, 23, 44, -24, -128, 52, -9, -23, 31, 59, -2, 0, -66, -27, 109, 22, -12, -6, 17, 4, -23, -40, 49, 2, -22, -4, -17, -36, 40, -19, -60, 38, 32, -35, 4, 24, -25, 14, 48, 52, 32, -13, -107, 4, 28, -78, -17, 74, 38, 36, -39, -34, -1, -23, -20, 56, -35, 8, -10, 18, -47, -45, -2, 93, 18, -4, 41, 60, -78, -19, 69, -52, -24, 23, -1, -94, 34, 49, 56, 17, -10, -55, -79, -57, -7, 91, 31, 14, 30, -75, -22, 47, 57, 46, 30, -100, -53, 42, -39, -34, 34, 38, -4, 61, -19, -65, -96, -41, 15, 78, 1, 64, 15, -117, 0, 64, -63, -34, 9, -8, 73, -12, 10, 32, -10, -28, 53, -31, -8, -24, -38, -10, 35, -4, -36, 20, 24, 20, 23, 52, -35, -7, 29, 24, -5, -1, 12, -18, 39, 43, 29, -94, -24, -22, -6, 20, -41, 2, 20, -17, 39, 68, -115, 8, 35, -22, -18, 10, -46, -41, 55, -1, 32, 75, 58, -18, -29, -36, 42, 53, 2, -4, -128, -42, 28, 92, 8, -39, 9, 18, -20, -2, -36, -10, 26, -66, -9, 72, 6, 29, 37, -31, -83, 14, 55, -11, 57, -4, -85, 7, 55, 38, -9, -49, -12, 35, 5, 72, -35, -77, -53, -32, 13, 8, -7, 39, 37, 2, -29, -38, -42, 29, 79, 46, -6, 64, -22, -27, -1, -23, -93, -4, -76, 44, 46, -27, -18, 29, -36, 51, 127, -1, -80, 8, -1, -49, 30, 17, -52, -17, -13, 45, -4, 10, 48, 42, -32, 87, -32, 8, -102, 35, -2, 15, -89, 35, 27, 0, 7, 94, 28, -90, -10, -5, -65, -25, 20, -26, 22, 91, 48, -44, -8, -56, 9, -7, 46, -26, 70, 42, 14, -92, -27, 10, 32, 58, 59, 5, -91, -60, 23, 56, -7, -30, -7, -6, -117, -38, 36, 48, 6, 40, 1, -56, -80, -27, 63, 19, 11, 17, 0, -25, 38, -27, -21, 116, 8, -52, -54, -22, -70, -19, 13, 53, 83, 51, 17, -7, -72, -78, 18, 52, 46, -29, -15, 26, 57, -9, 54, -37, -43, -31, 3, 0, 17, -63, 34, 38, -36, 41, 58, -15, 26, -27, -54, 1, -7, -43, 62, -8, -30, 71, 27, -55, -75, 1, -74, 73, 49, 28, -30, 17, -75, 100, 45, -46, -56, 43, -11, 72, 6, 40, -28, -9, -80, 46, 24, -1, -69, 55, 26, -11, 55, 66, -57, -55, -25, -22, 35, 32, 28, 55, -64, -28, 22, -10, -31, 36, -95, 36, 32, 4, 66, 20, -11, -19, 15, -93, 49, -22, 2, -17, 59, -19, -58, -23, 69, 77, -22, 48, 15, -28, -60, -34, -38, 61, 18, 38, 14, 4, -56, 46, -5, 15, -30, -39, -89, 34, -18, 52, 117, 9, -77, 36, 4, -86, -34, -6, -13, 91, 57, 3, 25, -20, 1, -41, 31, -21, -63, -96, 110, -6, -2, 3, -38, -91, 7, 102, 53, -25, -1, 62, -25, 59, -23, -30, -32, -2, -11, 78, 41, -11, -27, 37, -6, -83, -126, -9, 53, 65, 26, 89, 22, -125, -35, 37, 7, -66, 74, -53, 3, 21, 14, -60, -1, -70, 5, 7, -11, 69, -4, -27, 83, 37, -76, 28, 39, -93, -20, 58, 75, 55, 13, -71, -61, -12, -13, 26, 81, 4, -62, -20, -2, -42, 29, 27, -7, -75, -20, 74, 46, -41, -48, 13, 54, 46, -12, -29, -68, -19, 62, 10, 7, 0, -25, -52, -18, 19, 94, 28, 29, -40, -39, 8, 73, 37, 7, -37, -78, -59, 19, 0, -59, 10, 60, 20, 80, 22, -73, -95, 20, -41, 5, 100, -19, -30, 77, 5, -27, 78, -57, -83, 11, 2, -1, -36, -7, 35, 123, -17, 27, -20, -61, -128, 62, -5, -9, 6, 123, -2, -68, -37, 74, 12, -30, 78, -47, -69, 35, 31, -74, 63, 54, -34, -48, -86, 7, 13, 0, 26, 19, -55, -11, 22, -18, 43, 9, 35, 42, 57, -89, -10, 27, 6, 30, 52, -11, -77, -63, -42, -7, 34, 13, -62, -43, 29, 17, 21, 15, 13, 35, -17, 0, 82, 15, -78, 18, 26, -81, -8, 52, -22, 3, 31, -100, -17, 30, -1, 44, 3, -82, 19, 86, 55, -30, -32, -29, -37, 96, 40, -37, 0, -6, 22, 1, -5, 15, 18, -28, -1, -91, -82, -3, 89, 53, 25, 25, 22, 3, -9, -4, -23, -47, 4, -36, -30, 79, 5, 18, 0, -9, -47, -69, -40, 10, -20, 109, 99, -103, -9, -4, -20, 37, 68, -41, 57, -4, -80, -92, 18, 3, 83, -54, 10, 4, -43, -24, 86, -40, -34, 61, 43, 19, -40, -10, -61, 6, 28, -24, -54, 39, -37, -38, -34, 18, 94, 92, 70, -79, -61, 25, -7, -62, 63, -10, -36, -34, -1, -15, 47, 58, 4, -57, -23, 7, 36, 58, 60, -45, -9, 3, 15, -26, -24, -94, 17, -21, -14, 81, 60, -11, 30, -55, -88, 70, 52, -11, -11, 6, -82, -26, 57, 85, -14, -3, -110, -10, 43, 63, -58, 23, 14, 48, 29, -19, -34, 29, -5, 20, -53, -56, 64, -1, -97, 10, -39, -38, 28, -10, -24, 29, -49, 25, 76, 26, 24, 4, -62, 51, 45, -103, 1, 36, -92, 25, 75, 8, -30, 39, -46, -21, -65, 36, 20, 36, 38, 61, -72, -14, 25, 41, -15, -15, -37, -27, -26, 90, 17, 2, -43, -43, -58, 36, -49, 19, 80, 108, -32, -19, 0, -13, -57, 31, 82, -13, -29, -19, -58, -12, 24, -44, -39, 53, 10, 30, -41, 8, 85, 65, -76, 28, 34, -77, -41, 63, 63, -26, -6, -23, 13, -31, 13, 17, 10, -73, -42, 23, 51, -8, 14, 25, 2, -22, 1, -43, 48, 27, -3, -46, -45, -48, 20, 15, 40, 8, 7, 10, 27, 10, 32, -73, 24, 23, -52, -83, -38, 34, 56, -45, 24, 31, -60, -57, 37, -35, 41, 53, 20, 35, 35, -69, -45, 32, 72, 37, -58, -36, 5, 3, 14, -70, 30, 40, -23, -92, 46, -5, -12, -30, 32, -42, 95, 43, -42, -6, 77, 23, 81, -19, -10, -76, -76, -9, 122, 5, 0, -107, 2, 0, -9, -25, 49, 45, 21, -25, -62, 48, -28, 0, -7, 10, -61, 31, -5, 1, -5, 11, 86, -2, -40, 37, 0, -89, 62, -11, -23, -14, 42, -51, 43, 13, -40, -72, -20, -69, 70, 87, -25, -19, 72, 49, 55, -39, -65, -37, 0, 39, 30, -61, -47, -40, 10, 86, 80, -6, -72, -40, 20, 46, 15, 0, -37, -25, -32, -32, 46, 49, -23, -30, -35, -55, 58, 88, 68, 59, -8, -2, -14, -15, 5, 28, -91, -13, 6, -19, -83, -7, 46, 73, -30, -82, 26, -6, -13, 6, 8, 1, 42, -57, -39, 18, 92, 10, 32, -6, -25, -95, -5, -57, 22, -4, 11, -21, 96, 56, -35, -3, 49, -57, -61, 43, 54, 20, -76, 1, 29, 73, 57, -28, -85, -41, 30, 0, 7, 26, 127, -79, -3, -3, 42, 1, -42, -64, 36, 14, -36, -20, 36, -10, -19, 70, 72, -103, -18, -2, 49, 1, -80, 0, -13, -62, 75, 48, 0, 12, -19, -83, 3, -14, -11, 9, 65, 43, -12, 59, 31, 17, -43, -74, 14, -2, 34, -42, -5, -8, -11, -87, 36, -5, 45, 13, 35, -32, 20, -8, -5, -43, 76, -8, -41, 5, 38, 13, -25, -28, -63, -11, 2, -63, -3, 56, 62, 52, 91, -45, -72, -35, 51, -59, -42, 55, 71, -22, -37, -46, -32, -15, 37, -9, 19, 28, 30, 34, 83, 4, -79, -28, -58, -42, 15, 110, 95, 9, -54, -54, -1, 49, 26, -11, -31, -77, -41, 92, 9, -68, 13, 62, -36, 23, 78, -13, -70, 31, -10, -35, -70, 2, 93, 77, -87, 2, 27, -61, -5, 47, 35, 8, -6, -41, 51, -49, -46, -27, 26, -26, 24, 42, 83, -22, -23, 8, 42, -64, 25, -32, -124, -46, 90, 52, 26, 34, -40, 20, 21, -78, -47, -9, -76, 9, 31, -1, -12, 55, 3, 65, 13, 43, -56, 17, -42, -103, 11, 34, -43, 22, 109, -8, 17, -54, -58, -20, 10, -51, 26, 62, 42, -48, -31, 37, 56, -22, -23, 83, 39, -35, 9, 29, -24, 14, 40, -18, -60, -61, -88, 19, 81, 82, -9, 10, -51, -21, -8, 71, -5, -56, -12, 64, -92, 5, 32, -1, -25, 15, -54, 45, -15, 22, 80, 32, -19, -42, -74, 0, 72, -29, -17, -28, -3, 58, 59, -48, -88, -32, 29, 74, 1, 0, -55, 11, 69, 28, -99, -49, 7, 4, 0, -26, 19, 49, 106, 13, -70, -28, -26, 22, -15, 61, -28, 2, -6, 104, 31, -5, -39, -26, -77, -11, 22, 38, 2, -27, -2, 22, -17, -3, -40, -64, -17, 5, 80, 79, -23, 20, 24, 17, 0, -30, -72, 14, 26, 8, 60, 29, -122, -54, -6, 63, -51, 32, 5, 0, -2, 1, -55, 29, -8, -30, 17, -49, -30, 56, -1, 34, 42, 20, -27, 71, -78, 0, 66, 15, 17, 41, -70, -72, -11, 0, 23, 25, 52, 63, -63, -10, 24, -7, -24, 0, 14, -58, -7, -6, 17, -68, 8, 45, 28, -73, -49, 46, 26, -49, -9, -3, 41, 12, -24, 18, 51, -23, -38, -65, -29, 23, 58, 56, 22, -105, 2, 38, 37, -45, 30, 55, 1, -81, 4, 25, 14, 73, 19, -26, -24, -81, -15, 49, -48, 34, 77, -64, -30, 15, 59, 29, 58, 0, -125, -61, 43, 5, -17, 56, -56, 45, -23, 0, -21, 45, -48, 63, 53, -15, -23, 8, -48, -85, 56, 36, -65, 6, 15, -65, -76, 29, 42, 2, 36, 42, -47, 31, 18, -31, 19, 56, -96, 68, 26, -66, -40, 56, 7, -24, 28, 30, 114, 7, -56, -125, -30, 55, 90, -27, -35, -51, -58, -10, 87, -8, -28, -15, 58, 20, 0, 38, 37, -94, 15, 29, -74, -3, 53, -56, 43, 87, -37, -17, 26, -56, 24, 18, -85, -13, 93, -35, 12, 83, 1, -26, -69, -37, 69, -7, -1, -11, 41, -34, 65, -56, 2, -18, -35, -20, 30, 69, -18, 6, -51, 13, -77, -39, 35, 5, 63, 53, 106, -43, -18, -124, 0, 62, 127, -55, -1, -46, -30, 27, 55, -55, 66, 46, -81, -98, 12, 15, -5, 27, 1, 2, 26, 46, -24, 47, -25, -81, -43, 6, -19, -29, 75, 24, 21, -17, 13, 7, 32, -20, -53, 49, -8, 22, -45, 9, -36, 42, -52, 5, -48, 6, -51, 36, 90, 81, -1, -75, -77, -31, 70, 43, 15, 14, 2, -14, 88, 3, -110, -24, -31, -18, 30, 127, -63, -53, -5, 44, -6, 93, 12, -115, -54, -59, -37, 23, 96, 54, 22, -25, -74, -19, 48, -46, -32, 87, -3, -25, 56, -31, -110, -18, 91, 6, 7, 61, 14, 36, -34, -57, -70, -20, 7, 85, -26, 10, -13, -78, -19, 9, 22, -40, 53, -13, 24, -6, -24, -39, 96, 85, 7, -95, -38, -44, 20, -8, 45, 27, 77, -105, -13, -3, 95, 13, 14, -73, -42, -5, 119, 7, -21, 20, -42, -49, -19, 10, 20, -1, -82, 69, 28, -56, -6, 44, -74, 32, 49, -11, -117, 22, 24, -15, 64, 44, -13, -6, -3, -1, 44, -17, -37, -62, -20, 112, 20, -103, 25, 56, -24, -21, 68, -1, -54, 53, 48, -8, -65, 26, -35, 15, 12, 5, -66, -38, 25, 24, 55, 49, 0, -64, -6, -88, 64, 30, 15, 30, 31, -41, 59, -44, 4, 56, -4, -91, 27, -4, -99, -6, 66, 13, 59, 11, -89, -81, 24, 63, 4, -63, 37, -4, -59, -80, 24, 5, 92, -34, 53, 3, -39, -46, 35, 0, 22, -38, -56, -24, 32, 65, 43, -60, -5, 18, 20, -11, 37, 70, -23, -42, -41, 20, 0, 10, -53, 2, -25, 15, 21, 10, -18, 51, 26, 25, -41, -99, -28, -1, -53, 27, 49, -38, -20, -12, 19, 19, 71, 59, -12, -41, -5, -59, 68, 56, -47, -3, 46, -11, 54, 104, -13, -75, -42, -47, -21, 57, 13, 4, 21, -51, -12, 36, 11, -62, 35, -2, -10, 49, 90, -15, 17, -31, -31, -46, -5, 30, 1, -3, 35, 8, -9, 15, 13, -17, -83, -28, -18, -22, 44, 47, 30, 20, -45, -10, -12, -45, 76, 43, -99, 0, 37, -14, 25, 24, -82, -5, 24, 39, -6, 7, -27, -69, -31, 127, 25, -65, 1, -25, -30, 35, -28, -32, 124, -3, -14, 29, -39, -31, 77, 62, -37, 36, -65, 9, -48, 3, -1, 79, -88, -35, 27, -45, 49, 29, 0, -9, 18, -41, 11, 47, 34, 57, -79, -34, 62, 14, -72, -36, -91, -27, 127, 12, -6, 23, 20, -25, -47, -48, -26, 54, 11, 44, -4, -19, -85, 68, 23, 2, 25, -7, -51, 31, -17, -34, 36, 1, -22, 22, -29, -123, 10, 83, 47, 21, 47, -62, -93, 5, -2, 2, 43, 4, -8, 51, -24, -19, -9, -40, -39, 25, -5, 39, 108, 4, -26, -53, -34, 34, 42, -49, -7, -31, -88, 1, 121, 20, 32, 52, -94, -58, 66, -51, -38, 19, -10, 39, 60, 41, 5, -12, 6, -40, -29, -37, -85, 13, 81, 37, -24, -62, -31, 54, 58, 10, -80, -72, -44, -11, 127, 29, -40, -45, 57, 19, -28, -27, -14, -51, 3, 72, -15, -21, 62, -6, -4, 45, 102, -48, -66, -24, 40, -17, -15, -8, -59, 4, -2, 18, 68, 36, 12, -58, -30, -8, 28, -20, 7, -48, 48, 64, -49, -8, -68, -46, -12, 78, 54, 78, -89, -35, 4, 6, 26, 19, -72, -71, 31, 21, 14, -41, 12, -41, -19, -42, 9, 60, 109, -15, -51, -21, 80, -24, 46, 12, -86, -25, 35, 2, -3, -29, -60, 127, 9, -6, -3, -26, -42, 15, 17, 5, 7, 30, -56, -13, 41, 22, -105, 4, 58, 70, -46, 40, -13, -88, -45, -15, -1, 97, 83, -14, -40, -61, -23, 1, -38, 54, 72, 5, 28, 27, -82, -41, 54, 32, 127, -30, -80, -11, 46, 31, -22, -36, -23, 32, -63, 28, -29, -22, -125, 47, -19, 81, 23, -23, -1, 72, -64, -22, 24, 29, 18, -47, 22, -1, -6, 79, 56, -22, -1, -107, -10, 19, 0, -70, 51, -45, 5, 1, -6, 40, 57, -82, 1, 34, -46, -45, 41, 25, 93, -37, -8, 2, -5, -14, -19, -45, 31, 117, -14, 71, -22, -88, -128, 86, 15, -37, -14, 124, -27, -5, -34, -18, -55, -6, 26, 70, -19, 40, 37, 18, -5, -56, -8, 65, 32, -52, -36, -11, 9, -89, 5, 60, -9, 10, 2, 15, 30, 25, -81, -8, -12, -1, 42, -25, -25, 10, -12, -34, 77, 55, 39, 42, -26, -128, 18, 43, 69, -39, 51, -53, 17, 15, 20, -81, 6, 44, 35, -23, 20, 9, -13, -23, -31, 31, 29, -87, 13, 73, -35, 46, -20, -9, -18, -41, -58, 19, 10, 23, -18, -3, 51, 0, 17, -6, 30, 41, -1, -24, 44, 12, -87, -53, 74, -5, -94, 28, 53, 51, 5, -9, -31, -61, -53, -19, -3, 42, 57, 56, -8, -11, -10, 5, -89, -29, -27, 46, 41, 43, -12, -9, 54, -8, -26, 13, 6, -39, 45, -39, -29, -21, -43, -54, 69, 40, -14, 2, -8, -28, -1, 65, 25, -29, -73, 12, 65, 0, -51, 49, 2, -12, 20, -15, -42, 39, 15, -31, -30, -64, -39, 40, 54, -53, 2, 82, 6, 55, 61, -55, -6, -27, -22, 23, -28, 9, 35, -9, 1, -22, -21, 45, -40, -2, 27, -32, 9, 41, 54, 42, 26, -54, -44, -7, 19, 54, 21, -57, -41, -6, -23, 21, -25, 18, -40, -78, -21, 82, 18, -4, 79, -10, -15, 13, -39, -90, -30, 0, 15, 18, 9, 87, -3, -17, 23, 28, -30, 4, 48, -29, -82, -23, 66, 46, 5, 19, -60, -79, 34, 34, 19, 89, 43, -107, -53, -74, 15, 60, -1, -36, 68, 53, 31, -39, 6, -20, -65, -4, 75, 14, -21, 57, -21, -45, -31, 38, 47, 35, -47, -58, 22, -26, 10, 73, 83, 41, 28, -11, -41, -92, -107, 36, 43, 55, 30, 4, -63, -82, 8, 90, -5, -43, 65, -47, -43, 36, -9, -54, -14, 41, 45, 4, -80, -12, 2, 127, 7, -55, 41, 3, -58, 23, 26, -56, 45, 9, -71, 30, 10, -60, 45, 47, -128, 14, 52, -11, 46, 44, -65, -52, 0, -2, -41, 54, 87, -32, -63, 94, -17, 2, 36, -35, -9, 35, -8, -19, 35, 39, 37, -81, -62, -73, 4, 77, 25, 56, 12, -128, -39, 102, 6, -17, -40, 26, -14, 61, -13, -24, -61, 87, -37, 34, 82, 19, -92, -12, 3, -9, -21, -34, -31, 62, 61, 80, -4, -32, 4, -28, -20, 41, -78, -91, 59, 34, 5, 65, -35, -49, 4, 127, -49, -13, -81, 9, -45, 28, -23, 98, 3, -8, -49, -1, -31, -27, 9, 24, 57, 10, -12, 8, 57, 3, -66, 47, -8, -43, -31, 37, 2, 36, 7, 48, 29, -46, -95, 10, 14, -22, -41, 121, -5, -45, 70, -19, -54, 102, 52, -100, -20, 31, 12, -45, -41, 56, 63, -13, -96, 30, 21, -96, -1, 96, -73, 2, 80, -52, -20, 59, 4, -25, -14, -12, 8, 27, 45, 22, -57, -55, 34, 51, 18, 26, 10, -14, 6, 47, -7, -64, -122, 34, 52, 70, -39, -38, 34, -40, 0, 68, -36, -41, 3, -8, 20, 51, -18, 6, -27, 63, -29, 0, -23, -83, 31, 62, -81, -28, 86, -7, 44, 14, -14, -41, 5, 56, 11, -70, -88, 71, -37, 21, 61, 22, -102, 59, 11, -51, -48, -1, 55, 51, -23, 14, -29, -23, 14, 55, 14, 88, -6, -61, -93, -57, -38, 89, 66, 14, -30, -54, 15, 14, -24, 66, 4, -52, 25, 31, -36, -14, -47, 6, -52, 43, 60, 6, 7, 102, -6, -11, -111, 2, -15, 53, 6, 48, -87, -9, -57, 25, 29, 62, 26, 1, 19, -55, -99, 9, 32, -45, 40, 90, -103, -2, 29, -36, 2, 22, -47, 6, 9, -88, 94, 0, -12, 56, 68, -69, -46, -24, -27, 42, -5, 25, -13, -54, -45, 77, -21, -12, 72, 9, -57, 13, 14, -24, -53, 80, 17, 3, -3, 70, -38, -18, 28, -12, -91, 14, 79, -47, 21, 22, 12, -58, 30, -53, -5, -71, 30, 11, 28, -4, 71, -21, -27, 12, 44, 17, 23, -20, -20, 22, -11, -74, -5, 106, -40, -21, 76, 23, -4, 52, -28, 0, 2, -20, -59, -68, -32, 94, 40, -35, -32, -18, -70, -20, 57, 72, 52, 18, 11, 37, -64, -89, 13, 86, -25, -4, -17, 28, -70, 10, -19, 36, -11, -4, -44, 15, 76, 15, -8, 10, -25, -60, -7, -20, -13, 69, 14, -21, 1, -29, -27, 87, 76, -81, -21, 37, 31, 43, 11, 1, 26, -34, -54, -71, -32, 2, 63, 58, -17, -26, -30, -7, 17, 83, -10, 59, -24, -75, -36, -34, 6, -10, 55, -22, 47, -23, 31, -72, 77, 0, -9, 45, 30, -7, 46, -18, -61, 9, 40, 34, -70, -70, -53, -11, 14, 113, 6, -60, -40, 14, -31, -30, 69, 15, -15, -41, -39, 30, 87, 11, -92, 98, 0, 13, -36, 34, -36, 12, -20, 47, 69, 38, -69, -66, 31, 61, 43, 37, 2, -15, 18, -42, -34, -29, -45, -107, 32, 43, 107, -37, -1, 29, 37, -51, 46, -75, -9, 39, 32, -57, 13, -14, 36, 36, 45, -59, -32, 51, -38, -5, 12, -47, -108, 8, -9, 73, 46, 91, -19, -100, -128, -15, 69, 107, 37, -20, -47, 0, -26, -31, 18, -29, -37, -22, -22, 45, 72, 25, 56, -3, -93, -63, 29, 108, 29, -21, 56, -3, -95, -53, 23, 9, 53, 57, 60, -89, -68, -7, 3, 65, 5, -41, -82, -2, 22, 44, -54, 7, -46, -74, 48, 125, 31, -91, 1, 58, 12, 18, 10, -20, 5, -26, -86, -18, 69, 12, 40, 28, -32, -69, -29, 45, 2, 11, 0, 108, -15, -41, -111, 9, 72, 79, -26, 5, -45, 0, 13, 37, -89, -22, 28, 40, -9, -35, -53, -24, 56, 51, -25, 41, -18, 22, -19, 24, -76, 10, -74, 4, 18, 73, -3, 37, 14, -38, 13, 89, -53, -81, 87, 11, -78, -1, 97, -3, 6, -24, -36, 27, 34, 18, 38, 10, -87, -42, -24, 34, -39, 19, -56, 28, 45, -32, -51, 115, -17, -17, 99, 0, -114, 8, 70, 25, -58, -4, 31, -30, 5, 22, 0, -2, 10, -57, -15, -55, -21, -4, 82, 75, -54, 10, 27, -9, -85, 28, 56, 19, -115, 27, 49, 25, 35, -22, -45, 25, 11, 28, 11, -34, -4, 4, -76, -47, -10, 7, 72, 14, 28, -25, 5, -42, -27, -9, 48, 81, -5, 14, -22, 38, -74, -37, 34, 22, 17, -5, 5, -29, 5, -112, 0, 34, -2, -12, 125, 32, -71, -79, -11, -14, 55, 80, 40, -120, -2, 40, 0, 82, 34, -110, 2, 17, -64, -36, -8, 8, 56, 72, -5, -14, 8, -13, -59, 53, 36, 18, 4, -76, 3, 1, -43, -24, -32, -66, 58, 105, 13, -29, -42, -49, 2, 6, 45, 14, 5, 45, 92, -54, 1, -1, -22, -19, -39, 9, 70, -34, -45, 59, 0, -34, -9, -15, -17, 30, 95, 41, -54, -76, 9, -56, 46, 79, 29, -15, -3, -36, 23, 55, -51, -82, -10, 31, -11, 56, 81, -36, -92, -37, -53, -41, 46, 11, -42, 26, 95, 93, -18, -60, 18, 36, -31, 28, 34, -11, -90, -22, -9, -12, 18, -5, -12, 77, -3, 15, -9, -21, 5, 31, -4, 37, -28, 6, 20, -90, 32, 26, -2, -65, -9, -60, 35, 68, 15, -47, -12, -47, -19, 83, 58, -15, -7, 0, -37, 7, 45, 92, -9, -43, -31, -48, -64, 62, 23, 7, 18, -12, -54, 27, 40, 39, 49, -14, -39, -39, -42, -104, 56, 29, 1, -5, 48, 18, -23, 3, -31, 34, 1, 3, -128, 19, 20, 35, 37, 57, -93, 0, 32, -37, -55, 32, -38, -34, 88, 52, 1, -15, 29, -37, 70, 20, 1, -60, -76, 7, 64, 8, -40, 70, -42, -60, 37, 70, -60, 19, 36, 52, -17, 28, -24, -4, -27, 18, -57, -4, 29, -36, -43, 54, -7, 48, -14, 7, 46, 63, -110, -37, 49, 0, -81, 14, 44, -53, -24, 103, 0, 14, -18, -31, -11, 47, 55, -35, -18, -66, -41, 68, 31, -32, 95, 30, -103, 47, 51, -80, -4, -7, -7, -12, 6, -63, -11, -59, 20, 40, 10, 30, 39, 9, -5, 20, 40, -15, -42, 31, -21, -51, 17, 31, 98, 22, -19, -19, 15, -23, -47, -62, 30, 19, 69, 18, -17, 3, -27, -47, 39, -53, -9, 41, 20, -12, 7, -26, 72, 31, 18, -57, -61, -21, 9, 59, -7, -69, 0, 55, -12, -2, 53, -31, 41, -41, -54, 12, 56, -21, 91, 28, -106, -39, 12, -6, -52, 46, -7, 2, -21, 0, -96, -4, 37, 70, -6, -27, -7, 29, -20, 53, 24, -91, -23, 92, 20, -17, 7, -42, -45, -44, 28, 30, 98, 20, -108, -53, 29, 43, -6, -2, -8, 6, -46, 27, 69, -17, 14, -6, -7, 36, -1, -70, 19, -54, -88, 65, 55, 53, 40, -89, -49, 9, 61, -23, 37, -40, 1, -128, 58, -10, 21, 35, 51, -111, 9, -39, 60, 45, 56, -36, -29, -109, 86, -12, 13, 60, 111, -90, 21, 8, -11, -102, 30, 28, -36, -20, 81, 31, -51, 26, 0, 21, 1, 80, -59, -94, -17, 78, -69, -18, -19, -68, 38, 69, 26, -4, -11, -47, 11, -1, 71, 44, -66, -10, -51, 19, -21, 17, -7, 79, -43, 28, 36, -17, -19, -62, -41, 17, 98, -15, -14, -86, -3, 11, -1, -65, -41, -10, -3, 48, 52, -28, 3, 102, -7, -23, 5, 25, 42, -45, -52, 21, -62, 0, 120, 26, -87, -6, 12, 3, -46, 24, 46, 28, -66, 21, -55, -15, 15, 91, -45, 3, -25, 19, -104, 28, 8, -2, -22, 1, -32, 41, 112, 18, -5, 11, -7, -38, 56, 28, -63, -37, 37, -32, -12, 75, 0, -20, 18, -60, -29, 54, 6, -42, -9, 5, 40, 60, 43, -73, -7, -13, 1, -46, -27, 36, 125, 48, -37, -92, -19, 9, 42, -24, 10, 0, 61, 20, -39, -48, -4, 72, 24, -61, -18, 58, 5, -23, -39, -96, -23, 61, 127, 23, -44, -86, -80, -38, 85, 104, 34, 41, -32, -57, -93, -28, 12, 96, 15, 3, 52, -13, -7, 5, -25, -91, 4, -5, 73, 40, -1, -46, -22, 9, 29, 24, -23, -36, -5, 26, 97, -42, -51, 12, 48, -39, -21, -69, 6, 0, 0, -64, 62, -3, 65, 24, 19, -34, 81, -45, -47, 32, 9, -18, -6, -29, 5, 102, 17, -58, -98, -42, 22, 48, -24, 29, 27, -89, -5, 83, 17, 3, 99, -13, -80, -92, -19, -39, 18, 25, 61, 46, 73, -27, -49, -4, -28, 0, -46, 57, -19, 5, 68, 39, -66, 26, -35, -45, 30, 37, -14, -31, 39, 69, -98, 0, 8, -53, -8, -26, 23, 61, -34, -1, 75, -81, -5, 75, -52, -19, 72, -12, -45, 3, -64, 36, 68, -26, -12, 62, -66, 43, 59, -43, -37, 55, 44, 55, -19, -34, 54, -40, -34, 54, 42, -68, -64, -14, 82, -12, -1, -4, -42, 36, 26, -72, 40, 61, -31, 3, -38, 39, -17, 25, 18, 94, -78, -7, -74, 3, 8, 97, 57, -21, -66, -20, 32, 42, 3, -37, -90, -7, -10, 2, -18, 64, 12, 57, -68, 2, -29, 0, -28, 26, -12, 6, -47, -10, -5, 12, 12, -58, 57, 74, 11, -31, -5, 47, 38, -41, -24, -60, -32, 127, 49, -45, -48, 30, 9, 66, -31, 15, -73, -15, 21, 55, 25, 4, -93, -35, 29, 58, -2, 54, -54, 3, -47, 49, 17, 63, -73, 35, -42, -49, -25, -69, -55, 90, 15, 38, 66, -8, -36, -30, -76, 10, 6, -4, 39, 113, -21, -26, -35, -58, -1, 60, -18, 27, 29, -35, -60, 46, 41, 41, 0, -31, 7, 4, -17, 19, 55, -75, -69, -8, -18, 95, 53, -3, -42, 42, 6, 28, 54, -72, -39, -74, -7, 34, 86, -56, -20, -39, 72, -6, -1, -10, -26, 17, 61, -87, -45, 20, -49, 69, 80, -17, -72, 19, 66, -7, -3, 66, -34, -77, 55, 32, 28, 19, -91, -71, 15, 29, 29, 26, 55, -11, -9, -15, -17, -20, -18, -25, 37, 0, 54, -37, -29, -36, -2, -99, 36, 25, 47, -47, -39, -19, 44, 64, -25, 10, -7, 11, 8, -31, -41, -28, -34, 34, 95, -71, 31, 9, 0, 11, 47, -87, -37, 52, 4, 7, 45, 42, -100, -3, 4, 22, -30, 51, -2, -5, -37, -32, -76, -24, 36, 87, 53, -77, -73, 43, 42, -4, 1, 22, 22, -6, -48, -90, -32, 0, 49, 89, 47, -66, 41, -3, -60, 55, 3, -32, -31, 7, 45, 32, -124, -20, 45, 54, 17, -10, -23, -89, -61, 8, 64, 54, 47, -2, -86, -22, 60, 2, -46, -49, -43, 81, 96, 34, 76, -37, -71, -89, 40, 6, -25, -32, 15, -87, 30, 82, 63, -19, 28, 12, 55, -12, -4, -71, -69, -82, 30, 92, 45, -2, 27, 41, -13, -43, 11, -31, -82, 31, -18, 23, 7, 34, 17, 58, -75, 63, -41, -63, 30, -30, -18, 87, 0, -31, 20, -68, -1, -15, 18, 51, 44, -8, -2, -85, 76, 20, -77, -57, 58, 47, 82, 34, -27, -10, -6, 23, -26, -34, -88, 40, -24, 4, -81, 46, -42, 17, 81, 64, -96, -29, -36, -9, 23, -49, 45, 117, -7, -19, -22, 0, -13, 80, -15, 14, 19, 76, -20, 0, -77, -15, 38, -4, 15, -9, -85, 40, 26, -62, 14, -9, -29, 41, 127, -14, 1, 14, -18, -95, 40, 62, -9, -44, -32, 30, 12, 4, 34, 99, -91, -18, -66, 3, 29, 18, -76, 25, -26, 20, 29, -26, -6, 7, -21, 76, -30, -22, 6, 5, -18, 61, -38, -39, 28, -1, -69, -12, 9, -77, -41, 87, 45, -26, -47, -39, -12, 91, 74, 22, -14, 9, -31, 28, -26, -40, -57, -30, -25, 53, -59, -44, 44, 35, 112, 58, -88, -69, 64, 8, -74, -6, 35, -6, -73, 43, 24, 2, 29, 8, -34, 70, 9, -26, 28, 24, 21, -43, -10, 0, -64, -60, 6, 9, 78, 91, -34, -40, -17, -31, 12, 32, 2, -61, -15, -73, -26, 46, 127, 94, -43, -9, -31, 14, 17, 28, -39, 12, -39, -75, -4, 64, 90, -2, 43, -36, -108, -98, 61, 63, 25, 40, -4, -79, -60, 43, 32, 14, -31, 32, -44, -13, 25, -42, -7, 12, 4, 59, 76, -83, 9, -78, -56, 72, 105, -12, -48, -51, -14, 11, 30, 78, -3, -31, -6, 9, -44, 0, -51, 25, -32, 28, 98, 46, -30, 25, 40, -32, -10, 48, 24, -95, -98, 18, -43, 35, 35, 8, -111, 83, 46, -4, -85, 59, 45, -43, -9, 87, 10, -69, -49, 41, 8, 29, 9, -28, 18, 51, -73, -65, -9, -25, 97, 43, 17, -82, -17, 23, 57, -6, 20, 10, 12, -72, -37, -46, -39, 81, 74, -94, -63, -1, 31, 80, 68, 24, 18, -75, -38, -15, -65, -25, 41, -2, -49, 73, -12, 39, -36, 1, -37, -35, 0, 63, 60, -51, -14, -4, 28, -47, 40, -66, 8, 18, 22, -1, 71, 5, -29, -47, -29, 64, -62, 34, -12, 46, -109, 27, 53, -1, -26, 79, -22, -34, 6, -1, 17, 19, -64, -41, -41, 46, 100, -3, -54, 38, -8, -25, 49, -37, -100, -13, 25, 18, -2, 19, 88, -42, -23, -7, 19, 61, 5, -56, -91, -18, 11, 72, -75, 7, 18, 9, -71, 31, 78, 7, -75, 24, 27, 61, 24, -104, -57, 60, 28, -8, -43, -53, 5, -25, -15, 73, -18, 9, 89, 69, -60, 1, 26, -10, -115, -14, 87, 45, -37, 23, 40, -34, -40, -12, -62, 5, 73, 23, -47, -49, 47, 62, -69, -1, 65, -66, 12, 107, -14, -9, 70, -26, -10, 53, -63, -71, 70, -29, -28, -10, 2, 20, 47, 4, 35, -51, -37, -22, 34, -45, 8, 7, 25, -42, 72, -11, -11, -78, -6, 4, -10, -2, 98, -60, -47, 40, -43, 1, 14, 19, 8, 81, -78, 0, -28, -1, -44, -18, 35, 86, 39, -7, -18, 6, 28, 39, -9, -114, -44, 0, 34, 17, 64, -28, -40, -119, 2, -4, 71, 52, -14, -55, -3, -51, 12, 116, -18, -90, 11, 56, -58, 11, 77, -2, -12, -62, -28, 44, 4, -85, 14, 31, 13, -51, 62, 51, -82, -12, 73, 15, -52, 29, -9, -7, -11, 127, 21, -29, -105, -31, -26, 8, 53, 47, -88, 15, 35, -1, 69, 61, -24, -13, -25, -72, 55, 6, -1, -30, 70, -23, -19, -49, -11, -102, 39, 111, 55, -32, 43, 17, 6, 96, -19, -108, -49, 15, 13, 20, 52, -41, -28, -20, -28, -88, 77, 23, 32, -25, 28, -11, -53, -94, 37, 62, 42, 52, -13, -88, -36, 22, -27, 46, 32, -14, -36, -26, 3, 36, -7, 9, 40, 44, -52, -89, 20, -1, 13, 70, 52, -44, 39, 31, -102, -39, -25, -74, 8, 88, -39, 57, -14, -17, -21, -5, -25, 102, -60, -64, -11, 23, 12, -19, -12, -17, 18, 10, 13, 34, 7, -28, -7, 71, -71, 38, 42, -48, -19, 65, -72, -8, -20, 31, 63, 94, 28, -58, -56, -6, 0, -30, -1, -27, 113, -10, 30, 24, 4, -76, 18, 39, -25, 5, -35, -36, 15, 74, -75, 22, 21, 51, 2, -80, -18, 62, -34, -90, 0, 44, 10, -46, 70, -9, 0, 7, -29, -46, 68, 44, 41, 26, -21, -38, -7, -68, -31, 13, 8, -89, 58, -41, -18, 75, 81, -70, -17, 14, 15, 24, -32, -98, 2, 66, 72, -30, 54, -57, -22, 1, 65, -77, 47, 20, -6, -47, 11, -26, -22, -1, 60, 49, -62, -7, 56, -10, -52, 95, -7, -9, 22, -4, -79, -56, -10, 79, 68, -20, -114, -25, 35, 4, 41, 99, -77, -44, 52, 15, -109, 41, 22, -94, -17, 64, -26, 21, 43, -39, 71, 52, -73, -60, 4, 45, 4, 86, -52, -25, -79, 22, -3, 127, -51, 18, -43, -47, -26, 75, 27, -40, -19, -2, -72, -54, 71, -44, -25, 2, -35, 36, 48, -34, -1, 11, 17, 30, 42, -68, 30, 18, 4, -34, 18, -35, 37, -53, -25, 49, 38, 39, -2, -5, 14, 58, 64, -6, -22, -41, 1, -37, -3, -65, -23, -25, 49, 17, -3, 20, 8, 61, 53, -68, -112, -5, 82, -1, -4, 40, 19, -20, 23, 5, -19, -106, -52, 49, 81, -12, 8, -69, -6, -20, 72, -9, 53, -32, -63, 22, -26, -76, 31, 75, -73, 11, -46, 7, -20, 58, 25, -38, -63, -58, -27, 66, 127, -19, -44, -60, 26, 26, 23, 14, -20, 22, -6, -69, -95, -1, 9, -37, 48, -24, 2, 45, 83, -36, -13, -2, -36, 6, 28, 39, -58, -57, -13, -9, 28, -20, 41, 21, 58, -68, 76, -14, 1, 7, 8, -1, 26, -111, -63, 51, 71, 37, -11, 1, -39, 25, -7, -4, -80, 19, 2, 41, -23, 0, -29, 80, 48, -89, 4, 22, -64, -26, 47, -40, -8, 26, 27, 74, 51, -31, 43, -9, -81, -46, 18, 6, 65, 44, 78, -93, -79, 6, 31, -20, -21, -76, 39, 14, -58, 52, 79, -85, -22, 42, 7, -58, 14, 6, -21, 2, 17, 35, 29, -37, -24, -22, 5, 18, 12, -68, 51, -17, 23, 30, 72, -46, 4, -21, -35, 41, 81, -41, -9, -52, -17, 23, 23, -69, 45, -22, -6, 4, 40, -23, 5, -53, 74, 49, -48, -44, -34, -69, 3, 30, 39, -22, 44, 53, 11, -68, 45, -36, -59, -14, 43, 42, 69, -12, 31, -63, 15, -51, 46, 48, 69, -122, -13, -70, -31, 91, 39, 0, 45, 23, -37, 14, -86, -51, 6, 91, 47, 51, 28, -44, -9, -3, 6, -65, -89, -61, 65, 99, -10, -37, 29, 9, -80, -27, -62, -2, 43, 53, 64, 5, -58, 60, 4, -62, -40, 6, -18, 29, -22, 56, -18, 20, 45, -12, -71, 120, -1, -46, 52, -36, -58, -32, -46, -19, -14, 31, 98, 39, -102, 32, 44, -5, -28, 5, -7, -41, 42, 59, 99, -24, -47, -63, -31, -66, 11, 76, 42, 81, 32, -102, -66, 37, 0, 4, -18, -91, 42, 91, -3, -26, 47, -47, -21, 73, 83, -13, -90, -40, 4, -45, 12, 97, -11, -30, 44, -48, -7, 25, 47, -48, -15, -17, 56, 4, 38, 7, -47, -5, -19, -46, -27, 7, 3, 15, -28, 54, 54, 5, 29, 59, -66, -85, 3, 88, -24, 14, -37, -6, -15, 74, -64, -55, -30, -7, 3, 44, 41, 24, 19, -103, -15, 47, -11, -22, 6, -20, 4, -22, 6, 11, 76, 64, -14, -53, -65, 24, 65, 20, -52, -11, -10, -30, -1, 3, 2, 36, 89, 14, -6, -73, -39, 30, 97, 2, -6, -53, -2, -5, 69, -18, 12, 40, -6, -4, 29, -28, -12, 35, -34, 61, 30, -77, -8, -1, -5, -17, 13, -74, -32, 20, 29, 36, 30, -68, -64, -2, 27, 26, 7, 47, 59, -21, 36, -28, -18, -52, -80, -34, 42, 25, 110, 20, -51, -90, -37, 29, 38, -3, 44, -4, 3, -20, -86, 65, 24, -96, 51, 10, -54, 53, 102, -23, -61, -71, -46, 2, 70, 21, -64, 52, 44, -42, -87, -2, 6, -12, -9, 62, 94, 10, 17, -7, 21, -91, -1, -26, 35, -43, -19, -56, 21, 60, -5, 27, -4, 5, -21, 47, -19, -27, -5, 41, 15, 2, 60, -13, -23, -39, -82, -14, 36, 70, 30, 39, -86, -65, 26, 18, -41, -53, 4, 52, 59, -28, 54, -38, -39, 20, -61, -44, 89, 45, -62, -73, 17, -3, 40, 94, 5, -57, 60, -38, -45, -38, -35, 60, 89, -10, 6, -19, 27, -10, -76, -52, -24, 15, 4, -36, 55, 32, -49, 15, 58, -5, 12, -32, -7, 13, -37, -52, 93, 52, -65, -9, 39, -92, 44, 51, 68, 1, -8, -88, 47, 4, 66, 52, 19, -52, -85, -23, 9, 26, -74, -9, 74, 57, -41, -36, -46, -54, -54, 74, 77, 29, 11, -21, -86, 46, 63, 18, 56, 6, -51, -70, -1, 45, 56, -62, -97, 2, 14, -62, 3, 41, 25, 42, 41, -3, 41, -48, -79, 29, 0, -18, 13, 0, -87, 61, -3, -29, 70, 59, -80, -11, -15, -102, 31, 8, 36, 37, -32, -48, 111, -43, -21, 39, -65, -46, 113, 10, 29, 15, -44, -89, 25, -15, -10, 5, -26, 10, -3, 102, 0, 39, 7, 61, 9, 32, -99, 15, -35, -71, 15, 71, -18, 43, 64, 10, -98, -72, 47, -19, -55, 14, 78, -2, -21, -47, -42, -38, 61, 94, -8, -3, 52, -21, -109, -8, 28, 39, 24, 9, 8, 27, -25, -42, -47, -82, -47, 98, 18, 19, 49, -17, -55, 99, -31, -14, -29, -28, -18, 76, -8, 6, -56, -105, -23, 106, 31, 18, 14, -42, -31, 12, -45, -15, 15, -4, 77, 18, -39, -36, 96, -60, 10, 31, -27, -95, 76, 32, 9, 19, 7, -78, -40, -63, 41, 95, 88, 25, -12, -85, -19, -12, -52, -49, 30, 34, 69, 37, 22, -8, -22, -17, -52, 6, 19, 49, 23, -6, -80, 6, -13, -51, -31, 75, 29, 39, 102, 7, -68, -3, -9, -11, 5, -38, 91, -10, 0, 0, -29, -75, -12, -69, 74, 40, 38, 59, -9, -63, 27, -14, 23, 42, -59, -96, -22, 21, 3, 3, 66, 14, 8, 34, -48, -3, 34, -98, 31, 54, -109, 24, 31, -41, 2, 81, 9, 26, -38, -45, 36, -30, -14, 80, 41, 17, -17, -12, -89, 3, -4, 43, -38, 82, -3, 31, -20, -114, -29, 31, -25, -8, 35, -54, 49, 38, 58, -59, 11, -51, -70, -11, 59, 32, 80, 38, -75, 32, -4, 8, 37, -39, -22, 58, -35, -100, 30, -14, 19, -4, 79, -38, -48, -123, 9, 75, 71, -15, -74, -39, 52, 45, -32, 86, 40, -120, -12, 5, -45, 39, 104, -20, 15, -32, -58, -61, 44, 70, 36, -27, -32, 4, -58, 27, 72, 26, -90, -13, -37, -3, 49, -49, -76, 87, 39, -47, -47, 56, 11, 75, -6, -7, 45, 10, -127, 3, 47, -24, 23, 21, 17, -46, -21, -20, 52, -28, -15, -22, -47, 22, 88, -11, -32, 5, -20, 51, 30, -24, 97, -11, -85, -61, 18, -18, -18, 14, 43, -30, -48, 42, 11, -6, -23, 53, 45, 15, 11, 43, -40, -57, 69, 44, -20, -36, -20, 32, 59, -39, 1, -54, 11, 23, 7, -72, -7, -65, 32, 25, 35, 46, 20, 5, 54, -47, 4, -2, -5, 29, -12, -86, -9, 29, -3, -38, 22, 69, -64, 26, 36, -38, 28, 43, -56, -46, 71, 6, -81, -23, 14, -8, -23, 44, 61, 20, -7, 19, -85, -74, 45, 9, 80, 21, -4, -32, -45, -15, 117, -3, 7, 25, 17, 6, -47, -42, -26, 42, -2, -12, -68, 26, -74, -12, 92, 77, -40, -5, 25, 11, -3, 45, -55, 11, -48, -2, -43, 31, -11, 36, 11, 41, -75, -46, 25, 41, 30, 70, -39, -63, -86, 9, -15, 37, 25, 47, 4, -24, -17, -10, 25, -6, 18, -39, 47, -30, 40, -26, 18, -15, 3, -61, -1, -100, 21, 10, 35, 51, 85, 43, 15, -65, -39, -39, -52, -13, 23, 25, -11, 3, 29, 69, -23, -17, 34, 64, -36, -23, -46, 26, 59, -52, -35, -13, 81, -38, -13, -15, 54, 14, 58, -98, -26, 1, 1, 26, 46, -15, -26, -40, -8, 34, -46, -58, -45, 13, -3, 24, 28, 18, -9, 35, 3, -41, -51, -8, 41, 89, 46, -11, -4, -28, 28, -14, -75, -80, 0, -10, 96, 63, 12, -62, -45, -30, -21, 70, 5, -5, 25, 76, -112, -8, 21, 110, -19, -4, -52, -6, -68, 47, -21, -26, 8, 46, -77, 34, 17, 59, -25, 4, 28, 32, -112, 56, -14, -22, 59, 2, -41, 29, -94, -17, 28, -32, -6, 26, -82, 24, 22, 9, 48, -26, 15, 12, 22, -22, 58, 40, 51, -29, -46, -13, -35, 17, -44, 18, 0, 34, -55, 0, -39, 2, 25, 42, 18, 76, -12, -28, 10, 74, -35, -23, -88, -44, -10, 80, -29, 24, 34, -15, -11, -38, -31, 17, 44, -30, 49, -108, -14, 57, 12, -72, 1, -7, 5, 35, 0, -18, -55, -22, 20, 103, 53, -19, -10, 51, -8, -68, 0, 9, -35, 85, 14, -47, 20, 48, -122, -13, 92, 28, -28, 51, 25, -35, 4, -1, -77, -61, 17, 1, -10, -31, -12, 49, 48, 66, 27, 8, -51, -58, -13, 54, -34, 53, 77, -23, -25, 51, -55, -3, -1, -22, -42, 65, -40, -32, 10, 46, 7, 34, -73, -8, 34, 24, -128, 47, -22, 8, 61, 80, -105, 32, -37, -20, -4, 92, -28, 38, -34, -69, -70, 45, 39, 52, 17, -93, -7, 27, 1, 6, 89, -28, -25, -8, 51, -82, 9, 7, 12, -64, -10, 58, 42, -26, 1, -69, -36, 72, 48, -47, 43, -42, 43, -10, 63, -15, 29, -49, -17, -8, -7, -44, -21, 5, -32, 0, 79, -27, 0, 90, 0, -18, 105, -13, -115, -13, 46, 13, -65, -25, 66, 20, 37, 1, -76, 1, 66, -62, -18, 8, -73, -19, 103, 82, -38, 53, -52, -30, 45, 8, -38, 70, -29, -103, -3, -11, 24, 68, 52, -53, 11, 6, -88, -72, 48, 28, 30, 57, 17, -94, -63, 30, -24, 37, 85, 48, 19, -30, -70, -37, -3, 40, 51, -15, -8, 10, -41, 15, -31, 20, -8, 22, 19, 71, -95, 1, -49, -34, -12, 70, 4, -2, -8, -2, 38, -63, 20, 59, -49, -37, 121, 31, -71, -7, -77, -22, 51, 127, -38, -34, 28, 18, -66, 38, -11, -15, 31, 23, -17, -34, -9, -20, -46, 14, -41, -46, 87, 14, -30, -27, -3, -47, 14, 5, 27, -48, 35, 24, -1, -44, -47, 41, 110, 36, -20, -46, -55, -86, 29, 12, 45, 27, 103, -45, 10, -41, 17, -34, 24, 44, 2, -8, -31, 10, 66, 6, -69, -26, -37, -17, 92, 54, -43, -23, 9, -1, -65, 20, -56, 10, 25, 10, -42, -9, -82, 9, 14, -3, -21, 24, 17, 40, -31, 12, 85, 120, -24, -68, 17, -9, -89, 31, 81, -47, 18, 45, -75, -1, 4, 6, -81, 22, 54, 86, -80, -74, -52, 52, 87, -14, 41, -4, -47, 7, 11, -95, 9, 31, 36, 31, 98, -69, -32, 32, 14, 11, -12, -34, -2, 19, -53, 25, -120, -3, 40, 53, 5, 14, -46, -8, -12, -11, -10, 47, 58, 27, -7, -6, -35, 32, -32, 4, 15, 11, -28, -11, -71, -38, 2, 4, -27, 46, 43, 54, 37, 26, -78, -1, 61, 21, -79, -34, 55, -36, -13, 60, -19, -3, 75, -9, -21, 15, -80, -73, 38, 70, 59, 10, 24, -40, -46, -58, 18, -38, -1, -11, 30, -26, 90, 15, -10, -12, 18, -65, 77, 65, -60, -10, 46, -2, 38, 54, -93, -23, 14, 7, 31, 18, -36, -19, -55, -78, 0, 77, -4, -8, 0, 45, -17, 56, 0, 78, -70, -7, -2, 14, -1, 52, -98, -29, 21, -60, -72, 59, 34, -37, 21, 123, -27, 14, 38, -87, -18, 27, -13, 46, -41, -26, 105, 21, -15, 4, -14, -43, 12, -6, -20, -13, 6, -17, 92, 53, -37, 6, 1, 0, -11, -19, 2, 14, 38, 61, -87, -3, 14, -55, 31, 41, -88, -74, 3, 25, 56, 48, 71, -15, -117, -42, -37, 18, 72, -12, -23, -12, -28, 0, -24, -62, 96, 71, 5, 7, 32, -22, -45, 29, 41, -39, -9, -15, -73, 4, 73, 11, -44, 49, 0, -79, -63, 47, 38, 95, 13, 19, -17, -60, -116, 10, 5, 9, 64, 15, -71, -11, 119, -28, -72, -12, -14, 8, 18, 52, 15, 12, 5, 8, -89, -51, 54, -39, 74, 7, -75, 26, 34, -62, 8, 61, 0, 2, -13, -46, -4, 3, 61, -6, 48, -14, -78, -25, 51, -48, 5, 114, -28, -128, 18, 25, -26, -51, -1, 10, 73, 104, 3, -73, -34, 82, -22, -1, -43, -39, -77, 63, 5, -18, 52, 60, -107, 5, 24, 8, 64, 17, -6, 10, 10, -53, 32, -48, 8, -4, 19, -115, -14, -29, -3, 57, 114, -43, -23, 4, -3, -8, -19, -87, 57, 37, 51, 29, -73, -24, 1, 58, 15, -40, -29, 59, -71, 19, 120, -55, 5, -13, -20, -26, 1, -10, 42, -24, -19, -11, -49, 66, 72, -17, 37, -4, 6, -39, 70, -46, -55, -6, 69, 51, -22, -42, 24, 18, -34, 2, -71, -37, 22, 23, 21, 13, -37, -77, -46, 63, 22, -45, 56, 52, -48, -22, 90, 24, -51, -45, -43, -32, 0, 1, -20, 78, 88, -27, -31, -30, -28, -6, 48, 54, 113, -22, 18, -66, -39, 39, 17, -103, 44, 41, -88, 40, -14, 0, 36, 43, -91, -34, -12, 39, -24, 8, 22, 60, -25, 18, 19, -32, -53, 53, 26, -78, 13, 0, 62, -12, 14, 12, -43, -107, 9, 58, -11, -35, -59, 25, 19, 27, 88, -10, -128, 22, 8, -42, 1, -13, -53, -4, 64, 73, 46, -47, 7, -20, 45, -4, -2, 21, 30, -74, -6, 59, -21, -65, -3, 5, 7, 61, -42, -65, 4, 61, 23, -58, -21, 58, 37, -41, 38, 47, -56, -25, -44, -12, 11, 40, -73, 91, -17, -7, 36, -25, -53, -5, -36, 35, 23, -25, 51, 38, -47, -21, -8, 31, -9, -20, 58, 7, 11, 22, -77, -88, 63, 69, -53, 32, -24, -6, -62, 2, -3, 34, -15, 20, -68, -6, 52, 6, -21, 61, -14, -21, -53, 3, 2, 96, 4, -9, -21, 66, 12, -23, -5, 44, -3, -42, -28, -14, 18, -86, -15, 103, 62, -60, -24, 71, 6, 1, -7, -55, -79, 35, 60, 54, -5, -3, -38, -53, 17, 36, 21, 48, 104, -36, 3, 19, -17, -128, 51, 13, -26, 44, 61, -23, 42, 12, -79, -30, -15, 48, -21, 18, -40, 11, 56, 49, -96, 6, 51, -31, -2, 8, 23, -57, 40, -19, 73, -51, -35, -11, 21, -71, 37, 28, -69, -12, 102, 0, 12, -18, -39, 12, 70, 2, 43, -8, -74, -10, 5, 22, -42, -28, 23, 71, 21, -25, -28, -2, -22, 17, 24, -39, 17, -34, -21, 23, 31, -26, 63, -6, -42, -7, -9, -23, 11, -9, -124, 54, 9, 45, 51, 48, -94, -68, -2, 38, 4, -6, -7, 10, 42, 5, -62, -7, 24, 65, 65, 39, -79, -57, 98, -15, 27, 13, -63, -24, 78, -69, 48, -22, -44, 63, 18, -62, 56, -15, -91, 31, -15, -3, -24, 28, -9, 77, -51, 9, 55, 51, -64, -20, -24, -10, 69, 37, -24, 30, 58, -55, -36, -17, -8, -11, -22, -3, 6, -13, 82, 109, -41, -94, 19, -19, -36, 92, 40, -28, 6, -13, -122, 34, 74, 23, -1, 11, -93, -19, 86, -54, 25, 97, -38, -31, 80, 12, -128, -15, 44, -14, 43, -19, -32, 13, -25, -66, 38, -54, 31, 83, 7, 32, -11, -15, -22, -69, -89, 29, 46, 105, 75, -47, -38, -38, -77, -36, 100, 15, -60, 34, 29, -69, 9, 89, 34, 18, -26, 9, -14, -80, -28, 90, -42, -9, 88, 24, -21, 15, -80, -74, 93, 21, -39, -4, -1, 52, 8, 34, -51, -6, -81, 26, 20, 61, -55, -17, -37, 61, 36, -63, 29, 31, -81, -4, 77, -60, 6, 38, -19, -57, 58, -59, 5, 58, 20, 17, 42, -17, 22, -22, -121, -14, 79, 12, 12, 12, -38, -48, 31, -6, -43, -39, 74, 74, 9, -30, -1, -47, -5, 17, 127, -7, -74, -26, 52, 24, -36, -55, 31, 14, -91, -12, 46, 78, 39, -30, -91, -36, -100, 47, 80, 42, 48, 61, -41, -40, 44, -31, -3, -9, -21, -58, -5, 59, 11, -7, -14, -8, 0, 62, -23, -68, -53, -47, 107, 60, 42, -37, -6, -21, -6, -108, 64, 29, 60, 17, 9, -23, -13, -80, 44, 80, -3, 15, 1, -9, -25, -8, -28, -13, -13, 27, 32, 29, 49, -80, -54, 32, 83, -36, -44, -12, -41, 6, 6, 11, -12, 69, 37, 70, 21, -29, -77, 0, 44, -80, -27, 1, 31, -29, -61, -11, 25, 10, 21, -2, -60, 45, -31, 0, 34, 63, 35, 59, 13, -57, -122, -9, 62, 36, 54, 12, -29, -45, -48, -34, -14, 13, 78, -10, -42, 64, 100, -8, -44, -115, -48, 32, 78, 14, 61, -21, -46, -46, 59, -41, -15, -44, 71, 15, 46, -63, -89, 7, 11, 43, 49, -1, -60, -28, -9, 46, 0, 8, 31, 28, -54, -32, -23, 17, 53, 46, -93, -72, 5, 30, 92, -2, -25, 22, 5, -5, 36, -89, -54, 8, -89, -10, 126, 55, -36, -43, -21, 46, -22, -17, 63, -26, -55, 82, -2, -42, 27, -58, -66, 95, 63, 76, -38, -56, 52, -4, -90, 53, -48, -57, 108, 4, -23, 82, -20, -128, -29, 55, 23, -26, -37, -20, -81, 27, 102, 111, 65, -54, -38, -32, -24, -42, 34, -64, 11, 58, 76, -14, -20, -46, -57, 6, 59, 68, -14, -57, 31, 72, -78, 41, -6, -58, -10, 85, 32, 15, -49, 22, 43, -109, 18, 1, -120, -1, 62, 7, 71, 70, -98, -29, 29, -42, 22, 31, 26, -15, -60, -43, 53, -68, -31, 43, 23, 36, -8, -6, -26, -31, 65, 79, -2, 72, -43, -48, 26, -31, -36, 69, -41, -60, 42, 30, 107, -1, -41, -71, 25, -42, 28, 12, 8, -20, 3, -36, -52, 97, -4, 25, -73, 42, -44, 22, -18, 127, -62, -8, 44, 56, -60, -28, -66, -55, 66, 38, -2, -6, -28, -8, 65, 112, -17, -87, -25, 37, -75, 1, 58, 61, -39, -21, -62, -26, -15, 41, -51, -15, 5, 93, 54, -20, -31, -11, -100, 14, 121, 30, -20, 29, -57, -38, 52, 73, -35, -17, 30, 24, -53, 42, -31, 38, -15, -58, 36, 43, -123, -12, 14, -1, -36, 36, -25, 40, 19, 87, -58, 3, -14, 10, 22, 49, -97, -30, 38, -31, 26, 64, -12, 8, -25, -110, -6, 80, 53, 3, 35, -2, -43, -70, -28, -18, 22, 98, 55, -80, -29, -37, -39, 2, 38, 38, 85, 29, -23, -11, -40, -38, 27, -43, -8, 27, 34, 35, 5, -93, 44, 14, 20, 26, -9, -91, -23, 58, 5, -55, 41, -18, -44, 49, -3, -25, -14, -61, -62, -5, 104, 95, -23, -41, 46, -7, -75, 32, 18, -10, 12, 11, 18, 32, -25, -56, 17, -30, -9, -36, 26, 36, 10, 32, 35, 26, -64, -25, -51, -3, 65, 46, 32, 0, -3, -109, 59, 7, -37, -27, 73, 0, 55, -3, -61, -22, 44, 22, 23, -24, 15, 17, -72, -9, -25, -26, 38, 12, -18, 24, -43, -82, 70, 0, 85, -36, -18, 19, 57, -94, -39, 30, 0, -59, 34, 21, 0, -37, -38, 21, 55, -82, 52, -8, -38, 3, 77, -81, 49, 5, 20, -24, 59, -36, 23, 0, 46, -38, -28, -42, -71, -73, 78, 42, -17, -25, -46, -1, 96, 45, 49, -3, -103, -15, -30, 13, -12, 62, -7, -12, -26, 87, 2, 35, -28, -41, -61, 35, 38, 62, 25, 32, 12, 8, -91, 6, -12, -66, 37, 5, -28, 77, 12, -94, -53, 13, 27, 48, 43, -58, -89, 63, 24, -77, -17, -4, -49, 2, 88, 29, -47, 44, -19, -41, 13, 76, -4, -13, -65, -34, 17, -3, 61, 65, 31, -35, -7, 0, -7, 23, -37, -59, 32, 42, -97, 38, 25, -37, -27, 35, 28, -4, -27, 79, 23, -111, 5, -41, -51, 37, 59, -74, -22, 64, 20, -10, 54, 14, -24, 42, -20, -11, 8, -26, -46, -23, -27, 77, 64, 21, -29, -23, 86, 37, -39, 14, -3, -93, -4, 48, 8, 21, 73, -48, -122, -54, 17, 65, 0, -4, -8, 45, 35, 37, -71, -95, 2, 47, 48, 2, -24, -44, 75, 22, -51, 29, 20, -64, -34, 13, -6, -4, 29, 29, -15, -87, 66, 18, -24, -1, 66, 5, -12, -107, -20, 56, -3, 0, 18, -11, 63, 13, -31, -14, -68, -26, 127, -2, 5, 82, -77, -53, 27, -46, -39, 39, 7, 12, 53, 18, -39, -89, -21, -12, 28, 39, -24, -25, -37, 28, 49, 20, 48, 3, -43, -68, 24, 73, 51, -52, -30, -47, -10, -43, 49, 55, 5, -58, 17, -34, 45, 85, 45, -35, 1, 0, -74, -9, 0, 39, 39, 4, -106, 55, 15, -30, -31, 81, 45, 26, -43, -58, 39, -24, -36, -49, 9, -1, 80, 15, 54, -15, 63, -35, -45, -82, 9, -17, -14, 55, 6, -28, -27, 11, -57, 10, 3, -15, 1, 65, -13, -54, 97, -12, -22, 62, -13, -39, 69, 4, 6, -18, -14, -9, -10, -19, -10, -107, 8, 6, -37, 12, 99, -8, -13, -13, -53, -7, 34, 30, 37, 72, -13, 48, 14, -85, -56, -4, -11, -7, 83, 13, -11, -64, -66, -1, 20, -74, 22, 32, -43, 12, 90, -32, 2, 26, -20, 1, 61, 23, -30, -54, 2, 43, -54, 19, 70, -14, -75, 6, 19, 75, 99, 13, -54, 27, -18, -120, -20, 18, 47, 69, -38, -34, 23, 4, 35, 14, -66, -40, 46, -34, 60, -26, 45, -6, 15, -27, -13, -21, 0, 38, 8, 126, -46, -93, -31, -30, -53, 34, 27, -44, -20, 29, 55, 102, -9, -25, 14, -47, -76, 83, 7, -47, 57, 1, -22, 36, -54, -46, -8, -6, 28, 10, -53, -11, 12, -72, 52, 29, 32, 19, -8, -34, 100, -78, -34, 109, -1, -57, 43, -15, -27, 4, 10, -31, 5, -69, 27, 62, 44, -51, 31, 2, 63, -12, -23, 17, 31, -54, -49, -5, 27, 1, -19, 44, -38, -25, 97, -29, -27, 0, 37, -53, -10, -22, 54, -89, 0, 86, 39, -29, -25, -44, -54, 27, 81, -6, -44, 20, 55, -11, -21, -9, 76, 20, -10, -18, 13, -20, -86, -53, 42, 23, -7, 14, 80, -22, 6, -49, 2, -35, -5, -10, 74, -3, -69, -24, 26, -54, -36, 81, 5, -76, 32, 63, 39, 39, 0, 4, -8, -51, -41, -18, 9, 37, 12, -20, -28, 9, 26, 17, 41, -46, -59, 56, -49, 7, 127, -2, -20, -90, 0, -10, 43, 2, 93, -61, -8, -2, 26, 28, 87, -79, -86, 27, 6, 26, 24, -37, -61, 18, -85, 20, 19, 12, 60, 119, -38, -53, 3, 23, 12, -69, 3, 3, -76, -36, 113, -18, -3, 35, 12, -58, 12, -49, 56, -30, 38, -56, 66, -1, -34, -55, 76, 59, -4, -6, 10, -7, -53, 56, -32, -59, 36, -7, -128, 15, 48, -60, 15, 58, 22, 7, 72, -89, -9, -10, -13, -44, -37, -2, 91, -21, 3, 82, 40, 0, -17, 15, 0, 5, -69, 5, 6, 4, -77, 86, 46, -30, -25, 28, -2, -76, 10, 35, 0, 0, -28, -68, 22, 14, 3, -8, 58, 21, 39, 13, 23, -108, 29, 9, -42, -30, 27, -92, 58, 111, -15, -35, -34, -6, 95, 51, -70, 46, -6, -35, -51, -13, 17, 25, 62, 29, -52, -54, 88, 18, 53, -10, -69, -18, 14, 17, 5, 9, 2, 105, -37, 0, -34, -43, -128, 52, 43, -10, 18, 57, 8, 26, 56, -10, 21, -93, -58, -35, -37, 36, 21, 19, -43, 30, 19, 56, -56, 25, -89, -12, 70, 113, -25, -54, -45, 80, -53, 22, -46, -28, -12, 6, -27, 62, -40, 0, 56, 23, 37, -29, -114, 75, 11, -13, -22, 49, -44, 5, 51, 60, -57, -32, -5, -42, 0, -9, -7, -35, 0, 85, 58, -41, -1, 27, -56, 62, 63, -70, -28, 38, 71, 7, -58, -93, -2, 20, 110, 31, -72, -93, 85, -11, 19, 0, -20, -24, 109, -57, 26, 25, -56, -28, 115, -13, -73, -70, 0, 29, -23, 24, 121, -12, -70, 6, 60, -19, -58, 20, -14, -32, 48, 23, -59, 36, 24, -23, -9, 68, -48, -8, 21, -14, -39, 114, -30, 19, 0, -57, -87, 47, -31, -10, -46, 40, 39, 47, 27, 12, -58, -40, -13, 21, 31, 9, 1, -52, -54, -19, 51, -15, 40, 36, -15, -63, 107, -8, 0, 1, -32, -5, -13, -37, 91, -14, 3, -14, 11, -95, 58, -43, 6, -62, 35, -15, 36, 13, -39, -2, -35, 70, -20, 55, 0, 5, -42, 8, -26, 42, -4, -64, 10, 41, -14, 27, 86, -22, -52, 74, -9, -82, -31, -25, 21, 81, -48, 0, 62, 14, -49, -2, -44, -88, 38, 70, 5, 32, 36, -66, -25, 12, -53, -19, 62, 35, -15, -31, 36, -39, -21, 79, 14, -97, 26, 38, 39, 63, -47, -100, -7, 41, -30, -26, -78, 5, -1, 45, -23, 53, -29, 56, 7, 77, -25, -48, -40, 25, -58, -69, 100, -7, 14, 12, -7, -119, 54, -4, 71, -27, -21, 14, 96, -3, -86, -6, 14, 105, -25, 36, -56, -17, -95, 68, -10, 28, 47, -11, -77, 11, 31, 0, 6, -1, 38, 3, -46, 37, -71, -9, 10, 9, -36, 35, -49, 57, 14, 25, -2, 18, -48, -53, -90, 43, 9, 58, -28, 24, -19, 25, -23, 56, -64, 21, 6, 30, 53, -7, -79, -92, 29, -9, 2, 15, -14, -15, 24, 42, 0, 7, -62, 116, 6, -49, 8, -39, -44, 39, 22, 27, 8, -35, -69, 49, -38, 71, -74, -3, 39, 69, -91, 0, -3, -26, -27, 52, 25, -28, 22, 12, 7, 8, -25, -56, 19, 35, -22, 2, 4, 88, -68, -32, -9, 80, -95, 3, 0, -46, -93, 34, -30, 35, 83, 59, 1, 71, -72, -62, 5, -9, -51, 17, -51, -22, 61, 89, 2, -94, -19, 47, -12, -37, -42, -37, 74, 76, -5, -81, 9, 22, 56, -37, 0, 4, 51, 14, -6, -15, 9, -30, 0, 73, 26, 8, 68, -66, -77, 36, 7, -21, 60, -55, -83, 46, 40, -39, -28, 25, 27, -30, -21, -61, -28, 32, 21, -7, 70, 23, -30, -14, -25, 8, 14, 47, -26, -96, -71, 73, -8, -22, -42, 8, -3, 49, -6, 26, 12, -24, -8, -57, 28, 11, -37, -37, 72, -37, -19, 11, -37, -1, -30, -6, 103, 74, -59, 30, 40, -70, 7, 37, 1, 62, -7, -55, -21, -37, 44, 95, 60, 4, -29, -62, -9, -44, 31, 7, 69, -47, 3, -53, -12, 38, 3, -21, 75, -26, -66, 25, -4, 71, 35, -20, -52, -19, -75, 60, 13, 10, -46, -4, -38, 54, 53, -25, -26, -37, 37, -13, 7, 5, 44, 3, 42, -29, -44, -24, -61, 59, 64, -4, -7, -9, -38, 65, 79, -22, -21, -6, -36, -14, 37, 22, -80, 39, 77, 25, 7, -60, 7, -8, 11, -48, -9, -20, 81, -8, 59, -23, -53, 38, 24, -26, 32, -27, -21, 25, -31, 40, -2, 3, -1, -2, -102, -14, 22, 40, -66, 0, -48, 37, 0, 21, 46, 56, -46, -8, -76, -60, 104, 11, -6, 71, -24, -78, 37, -15, -48, 24, 53, -23, -93, -8, 109, 20, -74, 0, 46, -11, -82, 20, -23, 31, 43, 13, -98, 41, 44, 51, -11, -12, 0, 59, 5, -98, -59, 17, -61, 12, 110, -32, -27, -32, -34, 27, 94, 42, 11, -94, 15, -23, -70, 14, 24, -77, 4, 66, -31, -2, 59, -10, 13, 7, -7, -64, 55, -15, 78, -44, 45, 31, -6, -66, 9, -52, -87, 38, 90, 34, -56, -78, 41, -8, 14, 82, 4, -29, 53, -56, -22, 15, -17, 20, 38, -104, -1, -73, 36, 65, 29, -61, 93, -9, 10, -46, 62, -53, 13, 2, 85, -17, -51, -35, -28, 24, 8, 46, -69, 0, -45, 35, 46, 63, 11, -31, -94, -25, 61, 73, 43, 69, -104, -48, 5, 52, -46, -49, -5, 9, -35, 70, 4, -29, 0, -4, -57, 2, 59, 21, 17, -8, 32, -55, -15, -11, 32, 24, 17, -49, -35, 98, -42, -48, 36, 70, 10, 45, -14, -27, -18, 64, -40, 10, -60, 9, -47, 46, 18, -38, -106, 81, 56, -21, -15, -4, -44, 15, 64, -36, -37, -29, 20, 7, 6, -20, 32, -3, 61, 41, -19, -102, -39, 32, -19, -20, 13, -27, -25, 69, 28, 42, 36, 76, -61, -18, -74, 42, -53, 19, 49, 53, -116, -4, -28, 39, 12, 3, -26, 75, -27, 42, 17, -24, -53, 89, 13, 22, 9, -25, -55, 8, -37, 41, -7, 1, -28, -21, 30, -5, -6, 0, -30, -77, 111, -29, 56, 24, -77, -83, 115, 6, -36, -30, -23, 11, 116, 23, -7, -54, -38, -1, 113, -57, 0, 13, -3, -7, 18, -98, 17, 29, 24, 28, 32, -71, 5, 18, 59, 36, -64, -54, 13, 34, -63, -25, 27, -6, -2, 21, -14, -72, 81, -70, -18, 63, 70, 27, 71, -25, -108, -94, -15, 85, 20, -58, -63, 19, -1, -30, 13, 0, -60, 8, 127, 53, -4, 24, 0, 29, 11, -80, -15, 6, -106, -26, 89, 48, -34, 15, -48, 47, -37, 38, -119, 29, -6, 22, -5, 55, 0, -31, -44, 40, 22, -53, -7, 71, -54, 28, 51, -45, -24, 22, 13, -48, 76, -20, -18, -44, 41, -38, 58, 19, -97, -55, 69, 78, 35, -64, -46, 42, 13, 64, -1, -56, -123, 27, -13, -3, 2, 64, 56, 1, 1, -95, -2, 57, 71, -88, 27, 25, -64, 10, 20, 1, 9, 18, -27, 9, 22, -58, -32, 7, 34, 21, 13, -64, -15, -37, -45, 37, -38, 11, 22, -5, -55, 61, 47, 124, 32, -69, -39, 9, -20, -65, 34, -68, 42, 32, -3, -18, 54, -85, 10, 80, 15, -21, 53, -68, 0, 49, 53, -28, 13, -25, 35, -24, -80, -53, 15, -2, 62, -3, -39, 55, 8, -74, -95, 22, 41, 22, -13, 13, -59, -38, -4, 41, 117, 7, 32, 20, -86, -27, 55, -14, 18, 71, 4, -32, -102, -8, 40, 27, 42, 10, 6, -92, 6, -51, 4, 39, 63, -11, 58, -26, -128, -31, -38, -42, 35, 104, -11, 19, -24, -47, 38, 56, 6, 53, 1, 13, -25, -63, -39, -68, -66, 127, 53, -71, 6, 17, 19, -18, 49, -46, -10, -31, 111, -21, 13, -64, 1, -49, 27, 32, 47, -73, -6, -24, 43, 53, 40, 17, -15, -63, 0, -13, 7, 28, -13, 15, 29, -51, 71, 23, -23, -7, 90, -51, -34, -70, 76, 22, 27, 19, 7, -100, 25, 12, -18, 18, 10, -72, 0, 26, 37, 57, 49, -32, -86, -36, 75, 39, -56, -10, -20, -28, 59, 39, -68, -58, 56, -24, 38, 14, 32, -24, 122, -21, -107, 1, 34, -103, -4, 90, -39, 0, 1, -41, -25, 65, 53, 23, 18, 5, -104, -68, 121, 24, -37, -56, 8, 61, 1, -48, 0, -47, -76, 45, 95, 36, 46, 20, -22, -42, -43, -22, 22, 22, -38, 43, -47, -32, 17, 59, -100, 9, -47, -2, 41, 127, -8, -53, -98, -25, 45, 77, -30, 10, -35, -97, 31, 97, -58, -18, -18, 29, 52, -3, -66, 31, -24, -36, 44, 64, 9, -36, 53, -14, -64, -58, -34, 5, 112, 55, -44, 0, -5, 18, -35, -8, 53, 43, -97, -27, 92, 20, -62, -59, -44, 13, 75, 62, -27, -41, 14, 52, 32, 30, -105, -7, 18, -91, -10, 81, -28, 10, 18, -57, -42, 55, 29, 66, -23, 3, -2, 87, 17, -23, -29, -23, -52, -49, 39, 37, -18, 0, -32, 0, 45, 31, -85, -56, -2, 69, 11, 32, 24, -95, -49, 53, -7, -7, 35, 3, 54, 9, 19, -44, -79, -38, 60, 53, -28, -62, 26, -44, -19, -2, 32, -7, 59, -112, -10, 29, -9, -53, 29, 42, 13, -3, -66, 0, 15, 9, 40, 17, -28, -34, 80, -29, 27, -38, 98, -30, -49, -22, 66, -56, 8, 56, -24, 24, 28, -18, -28, 18, 13, 11, -85, -24, -51, 8, 60, 93, -83, -5, 12, 30, 36, -28, -38, 12, -64, -54, 29, 6, 28, -31, -57, -6, 20, 31, 115, -37, -34, -111, -2, 51, 47, -69, 4, -21, -55, 2, 54, 64, 61, 44, -87, -41, 39, 13, -70, -24, -60, 3, 102, 32, -2, -32, -18, 18, -2, -48, 73, -35, -6, 25, -11, -94, 72, -17, 51, 42, 34, -117, -18, 15, -17, 6, 66, -57, -38, 44, 4, 9, -32, -19, 59, 3, -56, 89, 1, -28, -9, 10, -66, -12, -30, 51, 14, -34, 12, 96, 28, 69, -18, -47, 21, -17, -49, 4, -52, -41, 107, 8, -37, -17, -12, -3, 93, 64, 32, 7, -27, -52, -22, 10, 41, -95, -29, 93, 11, -104, 13, 26, -24, -70, 61, -5, -1, 63, 20, -38, -3, 20, 30, 13, -18, 28, 7, 0, 19, -21, 12, 24, -48, -18, 40, 0, -13, 30, -70, -86, 23, -35, -15, 46, 103, -7, 13, 18, 20, 38, -6, -113, -49, -61, -12, 68, 11, 19, 37, -31, 5, -8, -85, -48, 0, 110, 49, -26, 4, 28, 22, 23, 43, -12, -119, -59, 18, -29, -38, 86, 21, -27, -13, 34, -43, 8, 71, 55, -59, -35, 94, -17, -93, 26, 8, -90, 17, -12, -1, 97, 56, 2, -21, -12, -37, -19, -89, 19, 40, 95, 0, -41, 5, 23, 43, -35, -72, 9, 1, -25, 44, 38, -88, -20, 76, 30, -40, -36, 54, 31, -1, -28, 29, -32, -6, 12, 15, 24, 31, -22, 60, -35, -100, -28, 24, 47, 45, -70, -49, -74, -27, 59, 36, 45, 53, -85, 2, 37, -24, -31, -47, -51, 78, 15, -28, 34, -42, -72, 74, 8, -13, 80, 51, -73, -12, 39, -15, -22, 24, 11, -21, 45, -14, -103, -14, 54, -23, 17, -9, -30, 26, -2, -42, 20, 11, -29, 74, 5, 0, 25, 115, -30, -52, -53, 35, -55, 12, 71, 35, -19, 7, -60, -30, -1, 40, 85, 8, -39, -34, -30, 20, 28, 49, -4, -40, -13, 29, 7, -36, -12, 0, 7, -72, 15, 36, 53, -2, -46, -38, -29, 9, 46, 30, -54, -91, 20, 107, 0, -43, 7, 41, 6, 83, -27, -35, -24, -38, -63, 31, 10, -41, -8, 69, 3, -38, -62, 21, -8, 92, 11, -19, -25, 6, -54, 21, 14, -1, -1, -18, 3, 28, 0, 2, 31, 12, -36, -77, 92, 6, -23, 14, 62, -72, 9, 41, 15, -37, 1, -47, 21, 108, 58, -62, -5, -10, 20, 34, -11, -40, -49, -46, -10, 43, 80, 80, -17, -12, -30, -77, 3, 35, 40, -5, 49, -53, -71, -34, 64, -48, -25, 98, 7, -25, -19, -34, -13, 117, -63, 11, 56, -1, -76, -30, -1, -40, 7, 31, 86, 26, -1, -110, -48, -9, 42, 68, 25, -100, -8, 29, -43, -17, 6, -46, -22, 22, 54, 71, 24, 11, -5, -102, -30, -27, 36, 72, -1, -88, 61, 7, -23, -10, 113, -32, -14, 73, 29, -116, 8, 26, 30, -11, 25, 14, -39, -98, 65, -20, -21, 45, -17, -86, 56, 74, 20, 58, -43, -128, -56, 99, 30, -65, -2, 0, 26, 34, 0, 4, -5, -22, -35, 1, -19, 10, -46, 21, -26, 35, -47, 19, 71, 39, -60, 13, -31, -42, 46, 24, 49, -11, -10, 14, 4, -106, -6, 45, 25, -13, -5, 77, 8, -59, -58, -9, 53, 5, -25, -64, -10, 8, 22, 14, 77, 14, 1, 25, -79, -62, 59, 14, -53, 46, 25, -74, 21, 42, -38, -2, -35, -40, 46, 52, -1, -7, 34, 18, -37, 21, -13, -64, 5, 105, -43, 25, 12, -41, -78, 120, 12, -36, -93, 5, -10, 45, 14, 41, -19, 12, -98, 12, 34, 52, 37, -56, -81, 46, 34, 13, 29, 27, -56, -20, 7, -35, -111, -4, -30, -15, 36, 102, 19, 15, -4, -68, -30, 9, 43, 23, 15, -43, -28, 11, 53, -19, 10, -29, -52, 26, -11, -36, -29, -48, 22, 83, 83, 69, 4, -65, -88, -22, 95, 24, -18, 63, -39, -70, 76, 7, 6, -15, -1, -37, -40, -65, 69, -6, -46, -9, 43, 80, -14, -12, -68, 18, -31, 71, -15, 41, -56, -23, -41, -55, -2, 66, 54, -22, -44, -57, 53, -25, 8, 22, -54, 3, 115, -3, -68, 88, -15, 7, 15, 39, -10, 42, -89, 17, -11, -49, -42, -20, -7, 55, 44, 77, -12, -11, -28, 59, -32, 38, -10, 82, -69, 3, 14, -58, -49, 35, 1, -25, -3, -69, -34, 34, 95, 61, -21, 45, -44, -7, -31, -57, -25, 109, 90, 1, -3, -7, -21, -119, -39, 70, 81, -49, -24, 57, 52, -41, -8, -91, -18, 41, 86, -18, 69, -34, -32, -58, -22, 35, 29, -9, -6, 34, -55, -24, -86, -12, 95, 66, -30, -79, 48, 3, 58, -45, 47, -22, 74, -45, -6, 7, 42, -20, 52, -47, -77, 71, -28, -37, 28, 0, -9, 24, -94, 32, -7, -30, 65, 75, -83, 7, 37, -64, -30, 66, 58, 2, 29, -43, -75, -70, 55, 79, 41, -7, -88, -39, -9, 11, -24, 37, 40, 35, -51, 10, 4, 12, 81, 12, 10, 15, -61, -98, -40, -91, 47, 73, 94, 35, -11, -105, 51, -41, 5, 6, 35, 19, 21, -71, 21, -8, -12, 14, -49, -18, 68, 29, 54, 54, -59, 0, -12, 2, 35, -30, -82, 22, -7, -52, -58, 12, 121, 75, -110, -23, 58, 44, 40, -3, -61, -14, -26, -78, 29, -3, -8, 55, 72, 7, 45, -15, -13, 40, -11, -17, -72, -21, -34, 52, -52, 53, 8, -51, -92, 59, 40, 13, 45, 0, 35, -56, -20, -71, -18, -28, 86, 17, -45, 36, 36, -25, -35, -2, -27, -46, 30, 74, 0, 2, 57, -76, -75, 48, 41, -49, 18, 64, 42, 6, -40, -64, 12, 1, 21, 39, -62, 7, 2, -47, -3, 91, 13, -9, -65, 17, 15, 30, 9, 70, -94, 14, 71, -6, -43, 110, -21, -64, -11, 18, -39, 57, 7, 27, -95, 29, -35, -30, -6, 38, -79, -23, 5, -4, -25, 64, 29, 35, 2, 42, 14, 44, -29, 70, -42, -18, 49, -24, -57, -5, 15, -11, 15, -57, -38, 10, 37, 24, 14, 18, 38, 10, -104, 19, -2, -87, 48, 7, -44, 47, 31, -2, -8, -3, 51, 66, -119, 12, -25, 40, 0, 26, -53, -18, -59, 49, 34, 57, 44, 9, -39, -117, -31, 48, 20, -64, -17, 76, 44, 25, 41, -17, -12, 43, -2, -89, -5, -74, 3, 22, -32, -24, 64, 31, -5, -3, 9, 28, 4, 24, -89, -85, 40, -37, 23, 27, 20, 40, 13, -104, 42, -9, -31, 60, 108, 4, -34, -3, -64, -15, 37, 45, -61, 31, -38, -42, -25, 34, 5, -68, 5, 41, 52, 56, 17, -17, 46, -22, -86, -5, -14, 30, -24, 29, -32, 49, -13, -30, -38, 56, -56, 42, 45, -18, 9, 114, 11, -22, -87, -57, -39, 46, 38, 0, -71, 55, 11, 38, 47, 66, -45, 42, 12, -116, -41, 30, -13, 22, 56, 32, -10, -6, -43, -78, -76, 47, 51, 53, 75, 37, -79, -59, -1, 5, -25, 23, 23, 6, -25, -92, 9, -19, 28, -48, 6, -64, 38, 77, 71, -36, 0, -77, -36, 19, 51, 24, 18, -94, 0, 32, 26, -27, -57, -31, 18, 5, 23, 10, -19, 17, 11, 0, -44, 1, 81, 26, -4, 49, 32, -2, 54, -73, -70, -36, 20, -39, 5, -37, 35, 71, 80, -43, -17, -35, -15, 32, 42, 37, 20, -36, -64, 24, 6, -18, -14, 11, -20, -20, -23, -24, 65, 65, -6, 12, -6, -111, 24, 96, 18, -75, 14, 2, 28, -2, -25, -38, 74, -17, -2, 49, -45, 2, 19, 9, -43, 51, -61, 78, -39, 5, -5, 109, 9, -11, -128, -41, 75, 54, 36, 19, -89, -62, 22, 15, 55, 12, -10, -10, -8, 65, 10, -3, -19, -58, -28, 71, -10, 66, -62, -34, 62, -17, -83, 20, 59, 39, 9, -91, -48, -48, -25, 51, 40, 38, 15, 2, 42, -14, -79, -8, 87, -21, -22, -36, 29, -96, 35, 15, 39, 56, 59, -128, -25, 13, -42, -45, -2, -22, 46, 44, 100, 12, -34, 2, 31, -41, -21, -64, -10, 29, 36, 68, -12, -57, 18, 41, 27, 86, -44, -61, 40, -39, -74, 48, 1, -73, 42, -22, -54, 79, 32, -19, -28, 5, -12, 40, -34, -49, 23, 62, 11, -64, 43, -4, -4, -9, 73, -4, -14, 57, 66, -48, -55, -46, -69, 51, 42, 0, 20, -10, -15, 95, 21, -44, -4, -36, -36, -40, 8, 51, 78, 68, 1, -37, -56, -6, 10, 89, 5, -1 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
