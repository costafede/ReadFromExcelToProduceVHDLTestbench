-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            -24, 102, 106, 65, 35, 103, 7, -104, 80, 85, -1, 98, 30, -125     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( 40, -96, -53, 104, 32, 71, 36, -92, 79, -81, -125, -38, -23, 123, 74, -108, 92, -6, -14, -85, -65, 104, 59, 14, 34, 60, 21, -118, 108, 37, -69, 0, -27, -31, 64, -53, 127, -78, -118, -23, 56, 87, 115, 93, 104, 107, -62, -92, 57, -117, 102, -86, 46, 94, -100, -89, 101, -102, 16, 113, -117, -73, 79, -32, 4, 48, 92, -101, -23, -86, -37, -15, 14, 43, 66, 23, -36, 112, -58, 40, -124, 114, -62, -59, 17, 29, 10, 27, 107, 69, 97, 49, 98, 114, -108, 42, 93, -57, 99, -6, 93, 30, 89, -49, -123, 16, 33, -1, 121, 126, 58, -42, 74, 93, -15, -52, -14, 98, 47, 26, 59, -68, -101, 50, 8, -22, -37, -52, -94, -85, 31, -27, -65, -79, 24, 88, -33, 89, -126, 110, 123, -90, -121, 30, 86, 20, 35, -51, -8, -128, 86, 46, -57, -12, -62, 36, -119, 93, 11, -56, -49, -119, -25, 96, -7, 117, 16, -85, -61, -44, 31, 116, -64, -87, 33, 21, 58, -120, 112, -52, 106, -66, 59, 88, -90, -85, -46, -57, -76, 21, 63, 86, -105, 63, -91, -120, 53, 121, -15, -25, 59, 110, -49, 72, -47, 82, 43, 3, 96, 43, -121, 86, 106, 57, 68, -55, -60, 18, -4, -56, 66, -96, -64, 116, -114, -102, 66, 18, 53, 20, 13, -120, 21, 100, 78, 29, 97, -4, -58, -90, -49, 25, -8, 119, -63, -22, 14, -112, 29, -103, -106, 124, -15, 119, 94, 4, 102, 20, 15, 52, 83, -22, -38, 110, -95, -18, -51, -33, -108, 32, 116, 23, 9, 40, -121, 73, -91, -121, -19, 49, -115, -120, 94, 1, 27, -121, -86, -1, -107, 94, -25, -43, 1, 60, 124, -39, -116, -117, 86, 58, -125, -89, -20, 101, -99, 52, 98, -113, 15, 14, 73, -35, -124, -36, 97, -16, 120, -8, 106, -105, 29, 103, 5, 34, 56, -54, 5, -61, -22, -24, -8, 114, -11, 123, -13, 116, 84, -58, 124, 126, 11, 71, 91, -121, -32, 77, -97, -97, 126, 15, 44, 121, -87, 122, -127, 100, 41, -95, 78, -3, 36, 11, 102, -78, 91, 106, 94, 85, 101, -77, 59, 6, 91, 91, -98, -120, 67, -50, 85, 66, -105, -118, -41, 62, 37, -106, -51, -57, 101, 125, -117, 67, 42, -59, -58, -32, -65, 39, 89, -112, -36, -68, 57, -48, -109, -43, -88, -33, 97, -46, 82, 88, -123, 89, -126, -72, -45, -118, -64, -127, 63, -110, -117, 36, -78, -112, 76, 107, -101, 113, 89, -74, 103, -116, 66, -29, 105, 3, 51, 13, -41, 84, -22, -72, 3, 68, -9, -80, -4, 126, -109, 107, 34, 19, 108, 52, 74, 50, -76, 68, 96, -37, -114, -85, -53, -82, -63, -9, 23, 21, -125, -118, -62, -61, -103, 11, -83, -4, -46, 8, -80, -91, -128, -75, -74, -20, 58, 58, -64, -100, -93, 102, 102, 4, 98, 24, 13, -13, -24, -23, 22, 102, 60, 42, -97, 96, 55, 70, 28, -9, -48, 21, 97, 91, 117, -124, 123, -90, -34, -36, 97, -117, 44, 116, -30, 67, -69, -72, -79, -31, -80, -33, 108, -99, -21, -24, 72, -66, 12, 41, -118, -98, 39, 88, -84, -61, 91, -115, -104, -67, 115, -8, 49, -8, -92, 34, -49, -35, 76, -41, 123, 34, 49, 39, -80, -77, 58, -1, 37, -33, 78, 41, -88, -93, -91, 86, 20, 117, 53, -37, 62, 121, 112, 11, 19, 81, -41, 79, 0, -12, -87, 30, 90, -85, 82, 81, -72, 78, 51, -93, 51, 82, 21, 35, 18, -126, 75, -74, 24, -98, 21, -48, -118, -107, 37, 87, 76, 114, -12, 13, 106, -41, 117, 52, 69, -110, -103, -106, -43, 65, -48, 98, 31, 124, 34, -25, 28, 39, 116, 56, 2, 35, 91, 78, 80, -87, 15, -40, -24, -11, 107, 123, 19, 39, 26, 56, -95, -103, 10, 53, -33, 115, 39, -52, -109, -125, -12, -11, -18, 71, 104, -36, -12, 118, -88, 119, 115, 72, 57, -103, 4, 51, 120, -25, -7, 116, -50, -3, 13, -96, 15, 0, 28, 109, -123, 107, -123, 100, -88, 99, -36, -73, -24, -79, -103, 77, 28, 16, 111, 25, 45, -9, 26, -62, 22, -63, 122, -10, -86, -65, -31, 84, -71, -119, -99, -93, 35, -22, 51, 124, -106, 38, -36, 33, -67, 11, 98, -10, 84, -85, -70, -113, -122, -109, 83, -10, 89, 102, 7, -46, -25, -106, 62, 47, -77, -103, -25, 41, 80, 37, 41, -61, -58, 73, -5, 82, -48, 79, 104, 17, -23, -84, 98, -13, -93, 1, -69, 52, 90, 45, 38, 58, 16, -58, 118, 72, -113, -80, 111, -96, -27, 45, -117, 24, -26, -73, -73, -31, -68, 100, 76, 107, 38, 24, 124, -22, -23, 38, 4, 29, 29, 107, 102, 99, -76, 73, -120, -93, 91, -62, 9, -111, -100, -36, 20, 69, -54, -94, 85, 102, -99, 93, 116, 51, -56, 41, 82, 110, 102, -32, 45, 23, 72, -127, 32, 105, 21, -68, -86, 26, -1, 3, -92, 43, 30, 124, 126, -32, -41, -103, 3, 0, -81, -78, 75, -72, 89, -40, -124, -24, -109, 104, -107, 18, 2, 23, 123, -18, -61, -80, 120, -31, -72, 17, -106, 34, 104, -37, -101, -9, -63, -74, -11, 83, -48, 41, 95, 46, -8, 115, -120, -24, 0, 28, -14, 43, -5, -97, -49, -12, -43, 6, -123, -126, -68, 6, -69, -115, -103, 3, 69, 101, 3, 96, -75, -45, -81, 40, -29, -97, -74, -67, -82, -72, 120, 86, 106, 100, -34, 99, 117, -91, 57, -8, 22, 118, 48, 11, 118, -38, 8, 82, -93, -20, -78, 45, -15, -102, -108, -121, 113, -123, -35, -60, 11, -128, 104, -4, 87, 31, -44, -81, -120, 113, -115, 11, 100, 37, -50, -114, 58, -14, 29, 125, -64, -56, -40, 42, 31, 65, -117, 107, 81, -42, -66, -93, -12, -3, 69, -5, 28, -24, -79, -61, -94, 110, 36, 15, -10, 117, -30, 122, -14, 105, 81, -27, 55, -105, -77, 96, 75, -108, 1, 55, -29, -51, 83, 17, -81, 90, -58, 3, -14, 77, 49, 65, 119, -32, 102, 3, 31, -70, 62, 94, 34, -25, 124, 5, 66, -32, 79, -122, 47, -29, -108, -19, 82, 17, 104, 49, -13, -14, 75, -12, -112, -27, 18, -65, -113, -52, 33, 87, -27, -90, 97, 64, -71, 20, -8, -59, -37, 104, -105, -128, -121, -61, -31, -91, 104, 116, 40, 74, -63, 23, -116, 76, 112, 15, 60, 30, -79, -120, 125, 127, -30, 10, 37, -64, 58, -15, 63, 11, 46, -70, -128, 92, -83, -14, 7, -107, -31, -126, -107, 24, 59, -43, -105, 15, 49, 44, 37, 3, 3, 45, -38, 115, 19, 118, -125, 121, 51, 116, 81, 93, -14, -38, 24, -63, -16, -29, 72, -16, -10, -52, -43, 127, -128, -86, -96, -7, 117, -26, -95, 50, 43, -37, 100, -57, -100, -14, -27, 37, -32, -27, 102, -117, -54, 55, 33, 58, 24, -46, 49, 106, 50, -17, 105, 37, 17, -54, 60, 65, -56, -57, 37, -78, -122, -30, -72, 48, 64, 54, -84, -93, 31, 14, 96, 47, 68, -18, 46, 21, 124, -58, 88, 50, -21, 16, 8, -34, -49, -113, -24, 8, 47, 65, 30, 57, 20, -118, 18, 27, 63, 122, 27, 126, 116, -104, -107, -12, -101, -24, 10, -14, 15, -32, -119, 21, 93, -115, 3, -21, -113, -110, 46, -90, 90, -5, 114, 57, -89, 25, -107, 108, 66, 44, 58, 112, 114, -96, -91, 13, -63, -17, 5, 60, 8, -95, -48, 101, 7, 24, 23, 2, -56, -50, 114, 115, -7, -84, -96, 19, 49, -60, 56, -22, -123, 102, 97, 71, 104, 115, 127, -125, -16, -96, 113, -2, -108, 118, 62, -31, 79, 114, 66, -99, -69, 127, 43, 113, -11, -35, -3, -59, 85, -100, -101, -84, 29, 107, -47, 4, -12, 21, 84, 127, 101, 1, -5, 97, -72, -75, 29, -67, -25, 112, 59, -65, 68, 93, -21, -32, -111, -44, 35, 85, 38, -21, -78, -60, 32, -69, -26, -93, 10, 50, 95, -110, 31, -79, -13, 69, 127, -124, 25, 127, 15, -42, -76, 57, 102, 6, -22, 80, -77, -76, -98, 47, 105, 32, -38, 2, 48, 127, -54, -39, 44, 17, -97, 65, 113, -29, -21, -98, -37, -1, 49, 65, 99, 84, -47, -72, 43, -112, -96, -59, 50, -97, -35, -13, -126, -3, -105, 87, -55, -49, -101, 24, 81, 52, 91, 45, 84, -84, 64, 82, -73, 33, -1, -5, 49, -61, -19, -16, 23, 125, 31, -58, -23, 27, -99, 94, -105, -124, -55, 21, -110, -28, 125, 73, -29, 32, 84, 75, 40, 79, -40, 63, 27, 52, 39, -33, 102, -41, 75, -21, 107, 65, 76, 0, -103, 14, -28, 52, -60, -5, -56, -27, 108, -111, -99, -24, -112, 27, -52, -56, -98, 58, -91, -24, -106, 60, -117, 124, 123, 68, -24, -88, 21, -51, 85, -90, 114, -2, -121, 79, -88, -101, -37, -3, 45, 40, -85, -56, 76, -41, -75, 91, -67, -55, -74, -12, 26, 52, -39, -32, -48, 31, -71, 32, -43, -104, 20, -32, 59, -49, 69, 31, -41, 6, -114, -101, -2, -93, -20, -53, -96, -76, -37, -54, -123, 35, 59, -22, -30, -3, -59, 108, 77, 95, 41, 127, 104, -24, -10, 73, 84, -39, 25, -17, 34, -125, -102, -33, 46, 73, 16, 108, 34, 50, -14, -28, 124, 34, -128, 106, 73, 96, 47, 33, 120, 6, 111, 14, -46, -53, -70, -55, 123, -80, -106, 100, -29, 73, -51, -115, -24, -50, 35, 56, 74, 67, 33, 66, -31, -6, 115, 105, -71, 61, -128, 97, -72, -72, -119, -40, 89, 105, -4, -15, 50, 79, -15, 56, -18, 55, -90, 104, -109, -38, -79, -80, 21, 33, -80, 107, -64, 12, -63, 111, 37, 1, -66, -37, -15, 20, 93, -49, 90, 115, 10, -114, 79, 45, 30, 59, 92, -84, -60, -2, 78, 15, 16, 45, 85, 24, -50, 36, 94, -9, -61, 99, -67, 119, 75, -78, -47, 55, 30, 73, -110, -54, -1, 67, 35, 86, 75, -15, -38, -117, 5, -57, 57, -120, 91, -110, 14, -125, -113, -35, -117, -27, -34, -77, 90, 38, -103, -102, -5, 122, 36, -20, 19, 118, 0, 73, 80, -127, -65, -39, -76, -3, -64, -1, -66, 126, -120, 9, -125, -27, -113, 7, 126, -47, -64, -94, 18, -74, 1, -6, 16, -25, -39, 83, -8, -63, -101, -126, 114, -104, 75, -52, -87, 114, 37, 74, 78, -40, 100, -120, 4, 46, 45, -9, 42, -20, -88, -121, -65, -58, -40, -76, 13, 84, -103, -124, -125, 2, -82, 39, -41, 26, -11, -124, -90, -126, -116, 98, 22, -2, -76, 1, -96, -128, -53, -97, 9, 87, -71, -116, -11, 67, -15, -41, 28, 99, 111, -98, -110, 60, -81, 16, -25, -75, 79, -8, 109, 65, 68, -94, 54, -110, -58, 80, -5, -69, 23, 124, 62, -85, -31, -115, 78, 122, 36, 41, -116, 45, -92, 91, -85, 57, 124, -20, 4, -71, 94, 81, 47, -14, -39, -74, 81, 96, 123, 58, 63, -10, 116, -112, 10, 37, 13, 64, -65, -37, 109, 89, -103, -83, 28, 88, 50, 4, -115, -54, -61, 106, 33, -100, -57, -58, -17, 99, 23, 67, -33, -38, 100, 120, 56, 27, -56, 79, -124, -120, -41, -117, -10, 39, -44, -98, 108, -124, -42, 7, 46, 65, -51, -17, 92, -26, 121, 125, -67, 78, 28, -44, -63, 89, 120, 82, 6, 74, 19, 18, -58, 26, -73, 4, 123, -86, -46, 27, 24, -123, 25, 66, 73, 71, 57, -10, -3, -10, -92, -58, 48, 19, -81, -121, 12, 109, 85, 46, 83, -15, -42, 97, -114, -121, -128, 63, 23, -76, -69, 17, 86, -61, 1, -46, -27, 80, 8, -77, -4, 2, 81, 116, -31, 125, -55, 3, 109, 2, -40, -123, 74, -46, 3, 122, -64, 77, 108, -49, -53, 37, -62, -125, -127, 12, 114, -85, -28, 36, 19, 45, -127, -72, 89, 119, -84, -46, -124, 39, -122, -119, 13, 38, 100, 50, -70, -31, -106, 86, 7, 67, 108, -44, 18, -118, -39, -15, -100, -87, -95, -45, 42, -66, -108, -122, 31, -103, 51, 29, 117, -94, -56, 111, -70, 113, 94, -5, -87, -123, -90, 10, -39, 82, 23, -119, -40, -95, -47, 94, 32, -5, -55, 21, -90, 107, 40, -113, -31, 92, 61, 105, -37, -83, 2, 36, 6, -7, -102, -5, -44, 23, -108, 104, -15, 113, -28, -44, 47, -13, -88, -2, -115, 55, -117, 102, -50, 8, 114, 110, 12, 73, 35, -16, -127, -37, 115, 3, 120, -57, -45, -21, -36, -42, 84, -68, -62, -25, -84, -25, -98, 12, 74, 13, -11, -104, -19, 51, -88, -1, -112, 73, -49, 100, -56, 20, -16, -71, 0, -29, 59, -19, 5, -88, -21, 59, 109, 112, -6, 36, 42, 72, 26, -61, -80, -2, -95, -57, 88, 16, 13, -85, 64, 61, 34, 9, -89, -110, 72, -8, 123, -28, -38, -42, 104, 111, 111, -41, 71, 63, 68, -55, -1, 20, -50, -47, 43, 76, -103, -4, 44, -35, -38, 78, 43, -102, -23, -77, 94, 111, 101, -86, -84, 122, -70, -106, -3, 24, -62, -48, 97, -117, -30, 65, 16, -52, 84, -48, -10, 30, -38, -90, 72, 57, 96, -8, 5, -20, -46, -23, -122, 91, -105, -99, 75, -94, -54, 12, 126, -115, 16, -126, 99, -49, 14, 9, 96, 102, -102, -108, -111, 52, 77, -6, -70, 83, -62, -70, -72, 83, 49, -54, 45, 9, 83, 3, 16, -97, -81, -119, -25, 115, -96, 31, 81, -6, -116, 121, -23, -65, -56, 20, -16, -20, 45, 95, -96, 88, 43, 56, -94, -78, 80, 110, 66, -35, -55, 113, 40, 80, -95, -80, -126, 73, 76, -6, 75, -49, -71, -14, -63, -33, -79, 97, -102, 13, 47, -66, -59, -79, -18, 39, -17, 101, -37, -113, 112, 58, -63, 98, -72, 64, -116, 103, 42, -22, 65, -7, -84, -121, 61, -89, 12, 65, 32, -111, 52, -52, 25, -111, 102, 89, -77, 109, -47, 122, 60, -25, 22, 30, 73, -46, 97, 25, 121, -114, 104, 125, 52, 104, 4, -6, 46, -1, -41, -65, -62, -44, -13, 21, -62, 71, 49, -32, -33, 125, -100, 117, -104, 120, -117, -4, 19, 8, -116, -104, -52, 13, 20, 40, 20, 5, -113, 25, 108, -57, 89, 126, 72, 91, 55, -107, 102, 63, -88, -38, 97, -84, 112, -22, -122, -19, 14, -68, 63, 114, -80, -102, -16, 78, -66, 44, 114, 107, 72, -66, -7, -118, -19, 91, 76, 60, 125, 38, -38, 52, -14, 48, -119, 98, 91, 2, -91, -70, -89, -23, -91, 114, -107, 61, -22, 10, -3, -8, -97, 5, 120, 86, -82, -69, -102, 11, 53, 106, -84, -32, -62, -7, -117, -61, 92, -88, -68, 29, -107, -35, 120, 17, -26, -50, -106, -44, 70, 30, -115, 60, -93, 39, 90, -70, 125, 48, 44, 17, -9, 102, -69, -50, -2, -38, 29, -4, -53, -126, -87, -59, -80, 55, 95, -98, -107, 9, 15, -8, -76, 37, 40, 2, 60, -53, -25, -112, -79, -22, 55, -14, 35, -58, 108, 64, -97, -106, -105, 85, 85, -13, -115, -56, -51, 5, -16, -108, -41, 16, 40, 46, 55, -15, -14, -72, 115, 61, -51, -54, 100, -37, -44, 105, 28, -21, 0, -51, 103, 6, 117, -125, 97, -72, 32, -88, 111, -25, 95, 107, -121, 86, 76, -106, -123, -115, -10, 34, -123, 98, -99, 104, 16, -102, -49, -71, -10, -42, -75, -28, -114, 10, 98, 34, -1, -9, 73, -92, 121, -62, 32, -98, 119, 91, 58, 123, -111, -70, -25, 96, 104, 57, 120, -63, 70, -38, 67, 6, 95, 106, -100, -26, -117, 84, 116, -105, 10, -91, 15, -20, 47, 40, 56, -84, -87, -48, -12, -27, -119, 117, -31, -87, 33, 37, 32, 116, -2, -80, -89, -66, -2, -23, 103, 42, -73, -91, -46, -82, 82, 52, 97, 60, -126, 91, -34, -93, -43, -53, 26, 1, -50, 4, -80, 20, -112, 74, -91, 23, -11, -12, 17, -19, -21, 93, -89, -119, -63, -69, -92, -61, 91, -108, 71, 84, -99, -76, -75, 119, 64, -3, -52, -87, -85, 57, -26, 109, -108, -23, -25, -81, 91, -63, -29, -71, 52, -19, 80, 41, 85, -117, 40, 110, -69, -6, -6, 22, 24, 86, 10, -128, -59, 73, -33, 85, 107, -45, -68, 83, 33, -97, 63, -41, -1, 118, -14, 87, 103, 53, -49, 104, -105, -88, -29, 44, 35, 45, 39, -5, 38, 6, 96, -24, -13, 43, 77, 8, 31, 121, 72, -89, 85, -96, 93, 97, -121, 79, -21, 34, -19, 52, -53, 57, -118, -74, -60, -63, -12, -42, -51, 28, -15, 27, -92, -67, -106, 127, -63, -2, 107, 68, 43, -107, -119, -52, 69, -32, -37, 46, -76, 20, 120, -71, 2, -104, -125, -79, -60, 4, -59, 15, -106, 127, 3, 69, 48, 103, 59, 55, -46, 54, -79, -70, 123, 60, -89, -64, -97, 0, -123, 42, 56, 67, -40, -108, 108, 67, -17, 118, 4, -79, -34, -69, -77, 8, 49, 63, 40, 104, -99, -23, -51, -62, -115, -105, -116, -27, 15, 83, 110, -119, 91, 72, 51, -55, 9, 78, -118, -125, -80, 0, -53, -51, -73, 35, -88, 1, 92, -11, 45, 113, -64, -33, 47, -38, -82, -32, 58, 80, 87, 88, 26, 103, 34, 104, 111, -107, 40, 45, 28, 41, 22, 118, 78, -42, -77, 17, 26, -107, -78, 53, -79, 114, 16, -3, 47, 64, 95, -64, -32, -97, 87, 96, 37, -71, -9, 17, 91, -99, 110, 108, 68, -73, 5, 31, -39, 63, 26, -110, -66, 111, -87, -104, -101, 118, -95, -30, -36, -59, 49, -6, -2, -12, -114, 65, 20, 40, 120, -81, 59, -62, -125, -125, 68, 93, 13, -111, -13, 39, 89, -42, -111, 52, -15, -100, 42, -95, 57, 105, -31, -61, -49, -40, -67, -63, -47, 126, 92, 32, 20, -50, 37, 122, 58, -1, 53, 111, -12, -95, 64, -96, 68, -103, -77, -49, 10, -58, -66, 78, -83, 42, 78, 62, -117, 66, 84, 54, -55, 54, 62, -35, 76, -94, 34, 58, 51, 62, 124, -103, -125, 88, 54, -36, 31, -86, -41, -101, 69, -61, 12, -25, 88, 79, 15, -107, 83, 55, -125, -30, 18, 87, 102, 111, -33, 113, -92, 20, -12, 44, -60, 109, -117, 49, 121, 5, 81, -54, -33, 30, 15, -50, -20, -108, -28, -25, -24, 87, 81, -32, 119, 125, 35, 125, 76, 121, 49, 119, -122, -40, -17, 92, -124, 117, 61, -115, 120, -43, -81, -19, 3, 57, 111, -67, -77, -99, -105, -78, -66, -21, -11, 49, 81, -11, 52, 35, -25, 109, 23, 37, 62, 99, 24, 78, -38, 126, 77, 109, 101, -15, 104, -27, -110, -94, 102, -6, -24, 30, -49, 84, 58, -11, -53, -63, -49, 103, 13, -6, -95, 79, -16, -63, 37, -11, -60, 100, -52, -61, 43, 96, -118, 77, -43, 108, -126, -15, -23, -43, 63, -23, -72, -124, -25, -95, -19, -7, -76, 119, 121, 36, -67, 14, -19, -21, -10, -58, 43, -4, -18, -101, -85, 37, 8, -2, -123, -55, 96, 57, -103, 90, 60, 71, -118, 115, -59, 62, 34, 42, -76, 3, 91, 121, -112, -94, -7, 10, -22, 66, 32, -49, 60, -128, 118, -125, 106, -23, -20, 11, -37, -54, -119, 120, 48, -47, 72, 57, -58, -12, 64, -90, -3, -64, -73, -119, -17, 93, 14, -69, 53, 85, 22, -127, -102, 83, -94, -107, -119, 44, -24, 74, -68, -9, -2, 41, 105, -25, -98, 114, -81, -84, 89, 37, -124, -76, -68, 38, -94, -107, -87, 84, -97, 109, -76, -6, 125, -62, 109, 117, 84, 66, -77, 51, 122, -126, 98, -31, -17, -34, -14, 55, -26, 109, 61, 26, 26, 53, 16, 48, -7, -70, 125, -107, -75, -83, 45, 52, -2, 80, -28, 16, -55, 16, -77, -124, 6, -92, -12, -35, 13, 90, 72, -9, 66, -125, -59, -24, 11, 50, 87, 86, -3, 19, -122, 51, 60, 62, -113, -118, -45, 113, 55, -29, -17, 20, -15, 37, -53, 118, 124, 113, 58, 26, 108, -106, -25, 97, -128, 5, -74, -110, -69, -41, -120, -6, 103, 84, -45, -26, -8, -77, 97, -99, 57, -61, 121, 33, 20, 1, -9, 115, 126, 109, -86, 5, 122, -44, 14, -125, -126, -82, 33, 122, 16, -6, -49, -76, 60, -56, 62, -60, 9, -109, -42, -46, -113, -65, -99, -55, -45, -111, 103, -101, 120, -125, -101, -11, -92, -32, -121, -98, -63, -73, 52, 25, -87, -14, -35, 95, -79, 63, -128, 85, 116, 91, 23, -65, 111, 78, -91, 110, 113, -24, -1, -111, 96, 101, -47, 20, 84, 90, -66, -48, -29, 38, 20, 109, 50, -110, -93, -99, -102, -26, -124, 127, 14, -122, 91, -20, 108, -82, -10, -55, -15, 61, 60, -6, -49, -6, 44, 0, 64, -101, 113, -108, -61, -42, 23, 12, -31, -91, -35, 58, -9, 12, -22, -4, 52, -91, -59, 19, -19, -57, 27, -72, -112, -1, -126, -108, 39, -91, 116, 28, 63, 123, -40, -56, 4, 47, -12, 31, 49, 2, -45, 94, -79, 97, 103, 59, 28, -97, 102, 61, -39, -91, -104, 71, -24, 75, -45, 44, 60, -14, 24, -6, 94, -67, -87, -73, 60, -111, 17, -86, -113, -11, 10, 80, -109, -106, -14, 40, -100, -27, -39, -113, -97, 26, -92, -58, 37, 118, 123, -75, 100, -111, -106, -2, 39, 16, -8, 102, 69, 4, -128, -122, 4, 61, 22, 70, 67, 12, -82, 74, 22, -100, -112, 60, 71, -14, -88, 32, 19, 2, -89, -15, -73, 48, -91, -121, 95, -61, 122, -115, -80, -90, -35, -87, 60, -6, -94, 85, -13, 97, 30, -30, -25, -95, -113, 82, -27, 85, -21, -30, 101, 26, 104, -104, -31, 1, 53, 21, -52, 28, -14, -127, -95, -91, 118, -123, 120, -24, -19, 124, 121, -11, 66, -74, -122, 47, 5, -38, -91, -95, -18, 59, 58, 127, 124, 85, -35, -83, -72, -52, 37, -107, 113, -109, 93, 54, 112, -121, 116, -104, -104, -108, 121, 125, 29, 18, 50, -2, 67, -109, 81, -27, -44, -58, -98, -73, 34, -47, 84, 100, -61, 104, 23, 1, 100, -76, -46, 67, 105, -103, 14, -4, 117, -15, 122, 89, -117, -34, 90, -58, 85, 90, -61, 73, 41, 18, 53, 14, -70, -81, -39, -96, 117, 23, -2, 25, -28, 4, -119, 28, -53, -116, 69, 3, -47, 46, 48, 36, -110, -23, -70, -52, -76, 49, 79, -98, -73, 2, 51, 1, -92, 39, 80, 2, 34, 106, 69, 3, 34, -60, -48, 57, -36, -16, -6, -48, 122, -128, 112, 3, -79, -48, 14, -4, -102, -68, 59, -27, 32, 82, -126, 90, -17, 12, 63, -39, -88, 19, 16, 122, 22, 99, -119, -1, 117, 103, -57, -81, 121, -69, 17, -67, 72, -98, 35, -59, 91, -83, 42, 31, -3, 120, -82, -100, 75, -73, -76, -69, 112, 10, 0, -56, -47, 107, -118, 16, -97, -56, 22, -119, 64, 82, 32, -114, -125, -102, -19, 37, -2, 6, -13, 73, 87, 45, -63, -1, 39, -41, 87, 116, 43, -9, 108, 7, 21, -45, 7, 6, 117, -110, 17, -113, 58, 21, 10, -116, 106, -82, -37, 84, 0, -127, 101, -103, 9, -76, -125, -95, 42, -1, -45, 10, -117, -120, -39, -123, -14, 43, -97, 69, -78, 38, 115, 105, 110, 31, -16, 16, 11, 25, 9, -5, -119, -74, -10, 104, 70, -88, -63, -105, 21, -2, 116, -30, 25, -80, -49, -79, 123, -104, -43, 43, 117, 67, -128, 119, 37, 4, -121, -90, -115, 37, -91, -7, -74, 48, 56, 14, 84, -14, -8, 27, 83, -84, 57, 94, -98, -45, 110, -23, 60, -63, 4, 42, -96, 44, 17, -127, 4, 11, 84, 10, 12, -63, -109, 74, 15, 62, 33, 81, 27, 38, 114, 9, 25, -56, -128, 125, 61, -120, -77, -76, -57, -46, 104, -8, -22, -73, 79, -15, -115, 10, 100, -84, 18, -106, 37, -42, -43, 125, -71, -69, 68, 35, -99, 25, 22, -67, 2, -72, -55, 117, 60, 13, 84, -116, -128, -77, 80, -41, -110, 100, 127, -13, -22, -104, 37, -37, -1, -40, -116, 98, -38, 96, 109, 124, 7, 93, -95, 16, 8, -26, 67, 26, 121, -68, 66, -16, 115, -92, -93, -64, 79, -77, -5, -125, -38, 76, -116, -56, -127, -68, 16, 5, -17, 32, -62, -8, -2, -58, -91, 61, 100, 73, -87, 47, 26, -111, 7, 84, 47, 88, -54, 65, -30, -117, 115, 38, 8, -41, -75, -89, -75, 10, -91, 31, -13, 125, -111, -63, -86, -35, -39, 7, -5, -111, -120, 97, -58, 23, 7, -32, 4, -63, -34, 33, 60, 96, -38, -53, 66, 102, -91, -50, -42, 96, 21, 41, -45, 72, 95, -58, 68, 66, 5, 53, 121, 15, 9, -122, 67, 22, 78, 97, 77, 63, 62, 32, -81, -105, 37, -65, 120, 22, -77, -2, 9, -124, 27, 107, 73, -100, 93, 95, 79, 1, -57, 25, 27, 124, -107, 80, -99, 74, -102, -22, -15, 99, -14, 30, 82, -41, -57, -11, 79, -82, 56, 6, -103, 48, 19, -5, 62, 29, -111, 104, -34, -85, -98, -50, -110, 11, 113, 3, -22, 25, -63, 110, 116, -98, 28, -82, 122, -29, -117, -58, -68, 60, -48, -10, -45, 89, -66, -74, 90, -115, -3, 43, -39, 123, -38, -109, -125, -113, -26, 29, -49, -32, -71, -22, 62, 78, 67, 10, -44, -116, -80, 40, 86, 56, 108, -80, 43, 99, -48, -36, 75, 24, 37, -58, -65, -13, -106, -93, 5, -98, -73, -66, 21, 1, -82, 1, 124, -15, -84, 99, 80, -50, -79, -93, 34, -6, -26, -5, -95, -112, -73, 36, -119, 35, -13, 108, -86, 16, -45, 93, -20, 27, -28, -83, 36, -86, -95, 62, 38, -54, -21, 54, 34, 105, -31, -96, -63, 24, -76, -111, 14, -49, -48, -52, -92, -103, 58, -44, 118, -114, 49, -43, 105, 59, 100, -46, 125, 45, -20, 25, 13, -115, 126, 28, 27, -62, 40, 89, -107, -26, -7, 35, 68, -21, -6, -107, 31, -19, 64, 122, 111, 49, 85, 15, 34, 120, -111, 70, -67, -38, 84, -28, -24, 22, 30, 34, -44, 16, -5, -5, 79, 24, -62, 59, -105, -64, -50, 84, 64, 83, 3, 118, 43, 0, -47, -32, 38, -101, 32, -124, 97, -65, -71, 27, -51, 94, -16, -7, 33, 0, -27, 83, 64, 109, 110, 18, -28, 44, 46, 43, 38, -82, 2, 119, 23, 52, -16, 26, -57, 124, -25, 36, 70, 61, -53, 109, 45, 85, 14, -52, -110, 32, 68, -107, -51, 75, -124, -10, -79, -60, -72, 119, -62, 18, -34, -82, -110, 98, -83, -51, 43, 6, 91, 103, 91, -28, -20, 23, -109, -23, 121, -59, -113, 23, -68, -107, -53, -62, -22, 58, -124, 51, 32, -36, -71, -20, 81, -67, 70, -86, 102, -80, 91, -59, -89, -116, -45, -27, 4, -95, -21, -65, 57, 73, 59, 19, -104, 67, -1, 37, -112, 83, -65, 117, 22, -18, -118, 87, -101, -75, -125, 114, 52, 117, -17, 9, 24, 41, -103, -111, -63, 17, 45, 16, 110, 119, 22, -6, 111, 72, 56, -44, -55, -42, 60, 109, 15, 35, -8, 20, 15, -28, -67, 37, -116, -40, -34, -116, 34, 112, -12, -93, 11, -101, -108, -29, -21, -36, 27, -53, -43, 41, -99, 106, -115, 42, -22, -14, -103, -70, -45, 41, 89, -71, -20, -62, -58, 62, -92, -68, -83, -16, 124, -29, 17, 10, 99, 106, -73, 58, 115, -125, 38, -18, -27, 82, -87, 94, -115, -64, 45, 73, -62, 74, 112, 11, -66, -3, -30, -40, -83, -15, -84, 12, 95, -121, -81, -121, 116, 10, 39, -23, 47, 12, -62, 8, -18, 26, 42, 74, -14, -77, -126, 31, -93, 30, 75, -6, 113, -107, -41, -14, -63, 70, 85, -63, 82, -120, 85, -25, -91, -8, -126, 126, 41, 94, -16, -74, 53, 49, 55, 41, -58, -55, 77, -41, 52, 11, -41, 55, 106, -66, 71, 0, 17, -125, -125, 53, 21, -109, 76, -88, -118, -105, -84, -64, 102, -31, -58, -115, -36, -19, -48, -92, -61, -24, 88, 62, 113, -17, 115, 11, -103, 5, -44, 38, -120, 50, 26, -101, 80, -56, 17, -94, -69, -31, 0, 107, -45, -41, -116, -65, -14, 115, 73, 117, -20, -25, 47, -116, -114, -49, -106, -108, -66, 92, 81, 23, 4, 24, -26, -36, -115, 29, -54, -5, -35, 69, 59, -61, -115, 7, -22, 69, -5, 19, -53, -101, 35, 30, -110, -41, 87, -56, -98, 13, -122, -45, 100, 65, 9, -19, -125, 108, 111, -116, 0, -112, -28, -3, 7, 99, -10, -126, -4, 1, -8, -50, 24, -60, 55, -9, 42, -82, 47, -4, -74, -82, 46, -33, -110, -113, 26, 106, 93, 17, -44, -24, 99, -54, 87, -71, 7, -57, 127, 15, -6, -62, 109, 8, -82, 41, -123, 56, 88, -34, -85, -7, -9, 123, 19, 93, 121, -46, -75, -80, -10, 114, 39, 71, 114, 121, -106, -105, -125, -98, 63, 28, -60, -27, 27, -78, -84, -128, 125, -10, -70, -123, -124, -101, 95, 67, -123, -97, -96, -45, 72, 84, -87, -115, 56, 38, 52, -61, 3, -83, 75, 64, -90, 126, -120, -47, -51, -114, -114, -69, 78, 39, -12, -48, 39, -105, 42, -103, -102, 18, -12, -54, -29, 2, -10, 99, 30, -25, 112, -65, 30, -110, -44, -46, 28, 23, 89, -118, -24, -9, -50, -84, -89, 43, 3, 26, -50, 15, 56, -37, 2, -51, -119, -97, -121, -84, 3, -30, -88, 14, 82, 12, -116, 32, 47, -98, -60, 44, -78, -1, -100, 104, -80, 20, -86, -90, 91, -8, -128, -3, -59, -82, 15, 25, -81, -94, -35, 2, 116, -65, -58, 18, -21, 57, 75, 122, -128, -57, 105, -6, -111, 115, -77, 90, 53, -56, 108, 52, -82, 66, -36, 102, 31, -60, -57, 69, -10, 8, 81, -56, -24, 17, -42, 125, -110, -116, -95, 43, 93, -76, 32, -20, 19, 117, 104, 84, 21, 119, 16, 58, -79, -22, -103, -98, -18, -25, -50, 81, -58, -117, 72, -41, -39, 16, 61, -5, 102, 124, -121, -15, -35, 113, 113, 47, -49, -57, 21, 0, -80, -124, -111, 53, -5, -108, -41, 81, -37, -52, -35, 47, 53, 78, 78, -76, -93, 28, -81, 10, 102, 124, 55, -23, 108, 83, 40, -42, 21, -103, -74, 38, 56, 21, -60, -87, -37, 5, 96, 112, -1, 39, -46, -13, -26, 9, 49, 14, -18, 17, -4, -52, 71, -68, 88, 35, 91, 124, 0, 36, 124, 99, 16, 44, 98, -48, 109, 37, 89, 96, -78, 37, 111, 34, 121, 46, 120, -26, 3, -13, 118, 105, -96, -80, -38, -30, 40, 119, 101, -128, 113, 44, 96, -45, 112, 63, -83, -48, -88, -13, 83, 46, 41, 89, 22, -87, 106, 31, 120, 26, -62, 108, -106, 66, 97, 2, 62, 75, -62, -96, -53, 126, 120, -14, -44, -75, -106, -33, -66, -108, -84, 78, 46, 13, -59, -54, -101, -42, -1, -28, -113, -122, -125, 62, -60, 16, 95, -83, -25, -111, -103, -62, 39, 40, -61, -31, 9, -24, -54, 122, -76, 24, 59, -121, 113, -25, 75, 58, -121, 45, 123, -123, 42, -42, -125, -35, -65, 29, 87, -19, -119, 2, -46, 108, -10, -13, 104, 27, 99, 113, 69, -85, -12, -112, -74, -39, 61, -103, 57, 65, 86, -65, -7, 72, -94, 55, -100, 85, -19, 15, -62, 74, 95, -112, -100, 124, -47, 65, 113, 14, 93, 121, 5, 72, -36, 115, 113, -105, 63, 19, 43, -51, 13, -56, -47, 45, -117, 64, -91, 0, -38, 37, -82, 9, -116, 116, 68, 19, 127, -63, -54, 5, -116, -59, 102, 25, -13, -31, -81, 70, 53, 82, 38, -118, 33, -16, 15, 100, -16, 47, -29, -11, -39, 70, -30, -70, -79, 24, 85, -6, 4, -72, -3, 9, 98, -83, -65, -124, 85, 66, 117, -103, -61, 88, -11, -61, 81, 118, 31, 118, -27, 55, 60, 16, 4, 42, -69, -119, -124, -112, -74, 108, -112, 106, 20, -74, 99, -53, -54, -89, -113, -108, 54, -60, -110, -84, 45, -51, 20, -53, -41, -23, 103, 61, -3, -120, 25, 88, 29, 104, 49, -9, -75, -105, -97, -127, 92, -115, -39, -58, -22, -60, 109, 17, 40, 114, -102, -123, 104, -25, 90, 30, -4, -118, -32, 54, -92, -13, -13, -83, -79, 83, -49, 22, 115, -49, -53, -85, 74, 91, -127, -31, 65, -74, -49, 59, 82, -127, 25, 76, 121, -63, 55, -105, -21, 34, -88, -8, 69, -17, -120, 83, -26, 78, -36, 32, -4, -122, -22, 117, 74, -76, 48, -126, -30, 29, 47, -15, -48, 89, -39, 100, 8, 102, -16, 94, -4, 67, 124, -53, -113, -112, 50, -128, -110, -53, -82, -124, -37, 57, -12, 34, -26, 91, 7, 29, 54, 21, -55, -83, 37, 20, -52, 42, -105, 91, 85, 117, 90, 121, 49, 56, -118, -100, -87, 21, -49, -103, 21, 82, -47, -43, -1, -37, -85, -114, 6, -70, 63, -71, 124, 4, 71, 50, 87, -124, 106, 70, 45, 108, 93, 31, 101, -95, -101, -8, -27, -1, 105, 50, 93, -64, 55, -50, 33, 124, -4, -74, 116, 84, 81, -74, -66, -56, 57, -67, 68, -39, -54, -101, 90, -112, 72, -122, -3, -16, 6, 52, 70, 27, -127, -110, -48, -36, 124, -71, -102, 107, 126, -121, -50, 70, 0, -18, 118, -3, 105, -79, -85, 46, 121, 38, 120, -122, 117, -14, 59, 103, 49, 16, -77, 13, 40, 44, 42, 57, -1, 62, 88, -74, -113, -119, -56, 59, -25, 42, 119, -74, 15, -43, -26, -60, 114, 33, 65, -123, 13, 107, 66, -24, -120, 93, -110, -34, 97, -31, 80, 119, -126, -87, -37, -61, -123, 111, 16, -102, -34, 18, -13, 30, -58, -30, 52, 79, -17, 56, 51, 118, -80, 49, -106, 47, -71, -8, 94, -66, -76, 103, -32, -74, 64, -30, 80, 47, -40, -46, -11, -20, 61, 114, 67, -68, -7, 33, 21, 112, 85, 15, 0, 1, 113, 17, -81, 13, -95, 88, 2, -60, -17, 48, 107, 27, -53, -73, -34, -4, 34, -86, -94, 127, -86, 89, 109, -103, -113, 46, -43, 105, 74, -66, -123, -75, -38, -58, -73, -23, 123, -74, 119, 22, -32, 66, -78, 72, -119, -63, -108, 2, 59, 73, -39, -7, 30, 88, -14, -95, 104, -80, 7, 11, -112, -120, 41, -93, 102, -101, 63, -35, -38, -2, -101, 92, -68, -64, 101, -27, -101, 69, 96, 90, 124, 16, 42, 95, 65, -31, -69, 60, 97, -97, -2, 42, 102, -41, 110, 107, -46, 82, 33, 123, -94, -15, -89, 68, 110, -104, -120, -5, -115, 108, -125, -1, 1, -10, 53, 40, 28, 52, 125, 106, 50, -108, 94, -107, -51, 35, 26, 123, 117, -19, -10, -3, 50, -110, 96, 34, -6, -93, 119, 19, 97, 120, -64, 74, 87, -121, 104, 120, -77, -82, 96, -33, 28, 85, -81, -2, 32, 6, 86, -5, 120, -3, -109, 109, -61, 46, -106, -35, -63, 54, 27, 9, -115, 27, -84, -46, 53, 87, 48, -115, 101, 81, 118, 13, -123, 100, -3, 22, 4, -87, -2, -20, -63, -29, -46, 29, 48, 45, -12, 67, -78, 3, 24, 72, 46, -50, 12, -128, -86, 34, -89, -114, 104, -112, -56, 86, -85, 99, -108, 111, 116, -64, 96, 90, -121, -99, -21, -99, 48, -37, 105, -106, -42, 42, 6, -35, -103, 79, 68, 46, 69, 30, 45, -93, 75, -18, -14, -62, 111, 126, 47, -42, -27, -84, -17, 9, 37, 56, -23, 93, 106, -60, -71, -58, -100, 20, 84, -36, -22, -51, -18, -70, -75, 109, -39, -61, -53, -25, 71, 9, -127, -15, 111, -24, 58, -126, 79, 114, 46, -31, 117, 6, -32, 20, -83, 118, 115, -77, 27, -40, 67, 34, 80, -123, -101, 41, 103, -57, -33, -109, -20, -29, -124, -126, -41, 15, 10, -82, -24, -77, -97, -44, 65, 114, -100, 59, 88, -33, 93, 120, 65, 29, 38, -95, 95, -23, -25, 20, -79, -75, -95, 90, 78, -106, -72, -17, 31, -49, 47, -76, -91, -99, -44, 24, -11, -64, -119, -47, 97, 38, -54, -14, -11, -112, -90, -73, 16, 19, -64, 48, -23, -111, -11, -94, 100, -89, -53, -48, 13, 4, -91, 59, 37, -41, -111, 112, -71, -9, -74, 42, -64, -26, 53, 34, 27, -25, -51, 74, 123, 37, -121, -40, 72, 116, -58, 119, 122, -2, 20, 91, -109, -78, -127, -38, -40, -86, 58, 26, -34, 90, -60, -120, 88, -80, -41, 45, -59, 57, -114, -114, 25, 71, 99, 103, 7, 16, -66, 122, 110, 0, 57, -3, 8, 31, -117, -39, -86, -7, 72, 39, -106, -77, -118, 87, 97, 17, -22, -53, -111, -3, 66, -57, -57, 39, -43, 103, 21, 50, -36, 51, -43, -10, 109, 99, -26, -85, 27, 25, 34, 120, -83, 73, 88, 79, 50, 32, 67, 0, -98, -48, -40, -90, 5, -107, 11, -35, -125, -7, 120, 0, -13, 99, 77, 14, 17, -98, -28, -13, 95, -116, -22, 120, -2, 6, -89, 47, 45, 16, 126, 99, 32, -41, 103, -32, 124, 81, -3, 110, -62, -54, -110, -111, 69, 83, 96, -43, 71, -47, -115, -106, 36, 107, -1, 60, 37, 36, -128, -33, 121, -56, 0, -34, -35, -65, 91, -30, 1, 41, -107, 22, 67, -90, -50, -126, -16, 57, -38, 103, 35, -61, 15, 104, 92, 114, 126, 49, -74, 72, 21, -95, -2, -64, -4, -33, -57, 81, -60, -114, 73, -109, -55, -98, -82, 82, -20, 84, -72, -73, -101, 90, 6, -90, 99, 80, 46, 105, 57, -26, 65, -109, -4, 116, -1, 23, -62, -43, -41, -90, -76, -43, -101, 125, -120, -71, 117, 32, -43, -125, 87, -82, 57, 16, -47, 87, -10, -113, -77, -115, -91, 85, 95, -46, 89, 84, 81, 43, -7, 16, -75, 91, -124, 120, 90, 54, 27, 119, 96, 100, -36, 60, -76, -76, 26, -83, 39, 8, -102, -71, -84, -40, 53, 58, 82, -54, -3, 124, 45, 119, 37, -57, 78, 114, -101, 100, -112, -46, -19, -119, 123, 38, -93, 105, -65, -43, -66, -77, 26, -21, 105, 47, -78, -29, -80, -117, 59, 12, 12, 70, 64, -35, -12, 98, -125, 111, -77, -79, -19, -27, 77, -3, -47, -70, -56, -83, -101, -83, -46, -24, 108, 20, -90, -53, -26, -70, -12, 104, -114, -45, -86, 40, -42, -118, 74, -35, -73, 28, 29, 52, -120, 114, 70, -47, -33, -33, -101, -61, -53, 61, -95, 101, -52, 9, -58, 26, 122, 42, -14, 22, 14, -5, 126, -117, 39, 31, 113, -104, -10, -57, -4, 117, -103, 9, -109, -60, 113, 65, 32, -72, 118, 7, -68, -21, -50, -65, -125, -119, 82, 5, 46, 69, -71, 68, 81, 37, 66, 59, -101, -90, 8, -13, 13, -106, 101, -7, 6, -20, -41, -121, -4, 48, -88, -17, -79, -97, -79, 63, 89, -46, -77, 65, 6, -26, -92, -118, 71, -127, 10, 109, 109, -101, -114, -122, 35, -44, -22, 12, 83, -93, -102, -28, 28, 86, -71, -77, 57, 20, 123, -104, 15, 84, 8, 42, 13, 127, -72, 8, -52, -42, 88, 28, 67, 67, 117, 15, 11, 16, -31, 106, -113, -111, 40, -101, -81, 71, 29, 6, 61, -101, 111, 114, -111, 53, 113, 123, -46, -77, -15, 111, -30, 63, -78, -111, 41, -8, 34, 121, 95, -56, 30, -97, -121, -105, 48, -41, 32, -14, -54, -100, 99, -100, 111, 10, -77, 4, 54, 126, 10, 73, -103, -122, 37, 33, 98, 13, 92, 40, 21, -70, -24, -15, -2, 114, -23, 52, 90, 47, -58, -93, 125, 126, 30, -41, 96, -17, 104, 114, 95, -106, 21, 112, -92, -48, 9, -30, -19, 77, -87, 27, -6, 46, -37, 19, -66, 6, -93, -105, 18, -40, 20, 43, 64, -73, -33, 22, -93, 52, -21, -98, -113, -117, -44, -40, -20, -104, 44, -44, 84, -113, -92, 109, 44, 69, 14, -80, -16, 73, -42, -1, 77, 5, -52, 13, -2, -55, -54, 6, 92, -32, 88, -76, -18, -116, -84, 109, 28, 106, -41, -47, -10, -75, -29, -4, 92, -53, -51, -87, 55, 21, -102, 6, -52, 62, -80, 32, 97, -12, -5, 64, -127, 109, 114, 19, 96, 89, -8, -112, 39, -14, -5, -23, -75, -48, -38, 59, -79, 27, 97, 82, 100, -66, -84, -29, 55, 56, 60, 91, 87, 110, -82, -31, -57, -93, -101, -100, 119, -82, -101, -110, 38, 24, 77, -120, -21, 111, -47, 83, -88, -78, -27, 115, -35, -67, -27, -66, 92, -25, 118, 111, -93, 23, 122, 14, -41, 103, -11, -98, -110, 4, -26, 119, -92, -26, -94, 41, 71, 109, -61, -86, 80, 35, 117, 79, 96, 52, 102, -39, -56, -21, 125, 93, 22, -122, -109, 32, -54, 56, -96, -49, 110, 93, -39, 13, 104, -17, -119, 65, 108, -82, -125, -118, 95, -80, -41, 102, 53, -32, -50, 58, 56, -49, 52, -16, 7, -96, -36, 50, -123, 112, 87, 26, 106, -74, -86, 83, 67, -16, 71, 117, -15, 14, 19, -36, 120, 89, 94, 77, -7, 90, 88, -126, -76, -125, 74, 89, 76, 97, -4, 79, -112, 18, 5, -127, -86, -101, -101, -84, -91, -116, -57, 77, 56, -26, 41, 38, -124, 61, -53, -92, -43, 117, 100, -116, 9, -15, -20, -102, -14, -108, 96, 106, 94, 63, 109, -3, -27, -17, 127, -126, 93, -57, 33, 45, 12, -77, 76, 87, -30, -57, 95, -11, 8, -1, -119, -54, 87, -128, -95, 101, 74, -96, -110, 13, -111, 60, 83, 65, 78, -108, 3, -56, 71, 56, 6, -6, 49, 123, 22, -99, -120, -68, 54, 31, 44, 26, 62, 111, -109, -107, -128, -75, -53, -33, -25, 115, 53, 55, -94, -105, -105, 97, 95, -69, -27, -23, 73, 85, -76, -45, 3, -65, 27, 120, -107, -57, 55, 7, -128, -97, -76, -35, -63, 36, 1, -19, 122, -5, 102, 122, 14, 60, -64, 56, -37, -97, 12, -63, -11, 3, -62, 73, 106, 103, 91, 105, 25, 108, -117, -95, 98, -56, -26, 30, -111, 111, -60, 75, -2, -29, -120, -127, 60, -98, -110, -59, 21, 126, -102, -90, 20, 65, -11, -103, 25, 16, -30, -14, 81, 15, -105, -110, -8, -44, 39, 24, 80, -97, 75, 121, 8, 66, 54, 122, -30, 114, 92, 1, -51, -28, 95, 38, -20, 2, -104, -39, 73, -99, 11, -94, -98, -115, -6, 101, 30, 31, 75, -101, 57, 85, 31, 80, 39, 47, -33, 42, -104, 92, 48, -82, -21, -71, -94, 61, -5, -46, -26, -38, 38, 58, 35, 112, 81, 9, 35, 92, -37, 13, 67, -83, 121, 58, -41, 18, -43, -121, -88, 29, 95, -68, 16, 52, 59, 23, 16, -20, -31, 69, 8, 101, -113, 72, 100, 52, 89, -125, 76, -60, 24, 123, 40, 65, 5, 127, 55, -119, -91, 32, -42, -118, 44, 119, -82, -49, -22, -52, -53, 80, 81, 55, 108, -65, -99, 13, 90, -74, 0, 64, -68, 23, -111, -71, -59, 21, 33, -19, 98, 2, 120, -90, 80, -83, -65, 46, 29, -90, -14, 26, -8, -84, 66, 54, -66, 54, -52, -89, 54, -11, 3, 107, 14, 71, -8, 37, 124, 91, 92, -59, -44, 105, 51, 35, -92, -103, -121, 84, 10, 46, 123, 45, 42, 8, 62, -97, 74, 42, -59, -98, -76, -30, -101, 114, -15, 54, 105, -42, 66, -36, 26, 100, 126, -2, -95, 78, -23, -8, 5, 67, -38, -86, 46, 52, 97, -47, 12, 40, 112, 12, -50, 77, -72, 32, 97, -18, 68, -91, -44, -54, -27, 122, 40, -52, 26, 110, 116, 90, -67, 110, 53, -118, -4, -50, 20, -50, 35, -40, 125, 28, -96, 102, 71, 86, -36, 31, 9, 77, 16, -45, 22, -121, 58, -7, -113, -69, 88, -98, 106, -60, 27, -106, -104, 87, 34, 95, 8, 120, 100, -7, -55, 109, 84, -82, -114, 72, 126, 55, -123, -100, -93, 102, -81, 91, -77, -22, 5, -57, -44, 65, -73, -34, -33, -53, 113, 29, 67, -10, 36, -6, -86, -91, 113, -50, 47, 48, -86, -30, -7, 9, -41, -124, -92, -49, -58, -50, 76, 16, 91, 77, -13, -105, -115, 51, 69, -85, -29, 66, 127, 17, -125, -112, -15, -109, 14, -58, 0, -113, -99, -69, -16, -65, -11, 5, -90, 119, 82, -111, 9, -68, 85, -103, 6, 88, -55, 85, 11, -119, 51, 122, 82, 68, 78, -106, 51, 37, -21, 115, 93, -82, -104, -6, -100, 76, -41, 125, -59, 21, -58, 120, 115, 90, 16, 118, -20, 40, -116, 53, 69, -96, -83, 109, -57, -53, 12, 44, 4, -33, -29, -87, 15, -92, 56, -93, -30, 91, -9, -5, 119, -86, -96, 34, -49, -82, -38, -60, 18, 90, -41, -83, 90, 46, 38, -59, 125, -99, 67, -18, 121, -81, 92, 61, 123, 69, 32, 48, 41, -63, 112, 80, 75, 15, -45, -105, -70, 47, -18, 103, -30, 65, 90, 45, 108, -10, -23, 103, -68, 21, 74, -116, 46, -117, -22, -88, -71, -27, 123, 42, -111, 9, 39, 95, 34, 86, 76, -128, -116, -81, -124, -84, 92, 27, 64, -107, 104, -109, 98, 2, -114, -78, 118, 85, 46, -38, -4, 10, -107, -102, 13, 31, -108, -83, 86, -51, 0, -45, 5, -92, 89, -61, -79, -42, 4, -37, -122, 73, -5, -35, -81, -72, -46, -37, 84, -117, -90, 121, 70, -21, 53, -123, -48, 103, 10, 13, -115, 73, -39, -40, 90, 106, -64, -76, 113, 24, 18, -29, -91, -106, 113, 5, -35, -123, -23, -62, -98, 121, -38, 102, 59, 97, 15, 51, -89, -119, -69, -106, 108, 36, 87, 62, -6, -13, -7, 87, -89, 73, -17, -32, 72, 124, 77, 44, -118, -65, 124, -31, 122, 123, 65, 89, -13, -55, -128, -11, 57, 95, 21, 112, 37, 74, -119, 103, -23, 14, -50, -103, 46, 18, 82, -55, -48, -5, -16, 116, -107, -90, -14, -35, 16, 57, 49, 28, -54, 5, 61, 76, 113, -17, 74, -16, -98, 22, 41, -86, -106, 77, 19, 6, 6, 34, -78, 77, 13, -102, 84, 9, 38, 4, 74, 81, -110, -96, -21, -79, -23, -27, 48, -10, 5, -58, 105, 28, 33, 45, 99, -110, -6, 8, -112, 122, -63, -48, 118, -55, 99, -41, 110, -123, 102, 116, 1, -44, 122, -99, 77, 65, 28, -108, -110, 63, -74, -92, 86, -106, 109, -108, -17, -23, -61, -115, -60, 52, -113, 111, 115, -44, 37, 28, 114, -25, 87, -44, 10, -24, -86, 48, 36, -14, 38, -98, 120, -85, -56, -35, -118, 62, 98, 100, 88, 65, 52, -98, 73, -91, 43, -112, -13, 96, 74, 23, -89, -79, 16, -107, 14, -119, 6, -82, -85, 25, 2, 107, 49, 70, 37, -53, -49, 100, -104, -21, -6, 119, 40, 57, -100, 6, 75, 81, 30, -21, -23, -49, 107, -1, 8, -67, 57, 28, 2, 116, 11, -47, 121, -94, 14, -63, -29, -6, -65, 60, -112, -126, -61, 14, 44, 122, 42, -90, -55, 34, 110, -9, -119, -6, 66, 108, -38, -104, -127, -44, 111, -65, -14, 53, 38, 46, -4, 40, 97, 88, 125, -68, -40, -31, 30, -62, -72, 17, 32, -11, 1, 121, 9, -96, -56, 43, -65, 45, 23, 2, 99, -92, 29, -84, -4, -59, 67, 37, -128, -109, 44, 32, -20, 34, -29, -37, -11, 72, -101, -2, 65, -88, -85, 124, 108, -49, -80, -85, 76, -23, -35, -23, -65, 70, 88, -80, 91, 81, 121, -32, 62, -60, -2, -85, 62, 61, -15, -29, -79, 51, 24, 97, 82, -57, -85, 18, 21, -10, -109, 55, -45, 54, -120, -124, -69, 7, 25, 86, -38, -13, -125, 104, -88, 12, 6, 41, -113, -93, 90, -99, -14, 90, -120, 117, -99, -11, -110, -20, 98, -99, 89, -115, -49, -11, 111, -95, 65, -100, -91, 24, -2, 51, -92, -127, 111, -10, 12, 34, -17, 91, 98, -43, 72, -28, 105, -53, -103, 56, -105, -22, 61, 19, 86, -23, 114, 50, -40, 104, 118, -25, 105, -124, -89, -5, -25, 33, 118, 60, 0, 96, -16, -91, 2, -9, -58, -3, 126, 27, -83, -3, 31, -100, -23, 16, 109, -87, 29, -74, -13, 19, -42, 69, -88, 55, -116, -44, 98, 119, -105, -105, 6, 24, -14, 121, -107, 76, 4, -67, 79, -102, 41, 17, -105, 60, -23, 125, 78, 127, -25, -55, 100, -20, -61, -17, 124, 108, -42, 80, 123, -86, 66, -49, -8, -92, 25, 24, 74, 62, -38, -47, 4, 35, 48, 44, -80, -10, 83, 35, -45, -116, 0, 50, 14, 69, 12, 67, 70, -98, -2, -21, 110, 79, -113, -119, 97, 110, -91, 17, -75, -39, -85, 87, -48, 83, 41, -82, 32, 18, 54, -10, 1, 24, 3, -63, -88, -115, -61, 35, -60, 103, 63, 5, -43, 6, 16, -102, 98, 126, 2, 107, 100, -62, 25, 78, 119, -64, 94, -62, -102, 44, -40, -74, -125, 46, -110, 111, 8, -98, -124, -98, 8, -95, 91, 69, -30, 44, -111, 59, 78, 109, 9, 62, -101, 43, 45, -100, 17, -87, 75, -102, -96, 66, 42, -93, -19, 40, 117, 4, 68, -15, -44, -87, 20, 94, 34, -83, -83, 11, 93, -125, 61, -24, 107, 69, 66, -114, 39, 48, 108, -107, -98, -59, -83, -97, -33, 86, -28, 52, 92, -97, -76, 71, 79, 33, 101, -109, 6, -21, 0, 25, 61, -102, 104, -14, -29, 76, -7, -9, 69, 56, -15, -91, 110, 73, 0, -11, 90, 39, 92, 91, -33, 126, -101, 15, -51, 83, 94, 104, -81, -127, 74, 30, 116, 16, 11, 93, 32, -99, 124, -95, -70, 92, 79, -34, -98, -18, 122, -5, 102, 4, -42, 5, 88, 65, -119, -3, 96, 89, 90, -59, -41, -37, -44, 22, 45, 36, 107, 43, -98, -7, -50, 77, 116, -102, 74, 0, 113, 90, -101, -38, -35, -78, -60, -44, 82, 69, 97, -39, -80, 57, 46, 118, -41, -3, 63, -67, 74, -80, 116, 93, 69, -107, 67, 68, 48, -106, 91, -91, 18, -110, 4, -84, 112, -25, -9, 69, 69, 58, -6, -45, -42, -57, 44, 20, 20, 104, -101, 50, 78, -82, 53, 69, 119, -71, 51, 20, -123, 120, 117, 112, -53, -54, -70, -106, 4, 91, 104, -33, 122, -56, -94, 42, 16, 63, 28, -18, 46, -99, 70, 48, -91, -50, 60, -31, 30, 48, 64, -41, -44, 58, -81, 81, 0, 108, -102, 123, 98, -27, -122, 7, -78, 96, -106, 40, 62, -50, -4, -113, -37, 95, -82, 66, 52, 85, -54, 124, -77, 36, 32, 68, 79, 86, -21, -121, -15, -70, 123, 113, 77, -42, -43, 79, -14, -107, 93, 18, -68, -77, -41, -59, 32, 56, 77, 10, -50, -23, -119, 11, -57, -33, -63, -92, 76, 81, -84, 18, -127, -79, -125, 24, -124, -87, 59, -83, 27, -57, -108, -54, -90, 86, 62, -56, 115, -29, -100, -120, 68, 91, -42, 98, -84, -52, -29, -113, 40, -56, 94, -21, -85, 19, -81, 105, -114, 92, 114, -87, 118, -20, 113, -44, 66, 104, 9, 117, -26, 56, -116, 20, 85, -83, -21, -80, 4, 14, -73, -119, 46, 12, 89, -56, -88, 33, -42, 20, -47, 57, -90, -1, -90, 3, 49, 125, 109, -111, 4, 37, 81, -120, -7, -123, 64, -25, -115, -80, 31, -91, 1, 18, 118, -47, -38, -112, -108, -17, 70, 109, -128, 56, 10, 28, -78, -113, 56, -124, -25, 83, -124, 81, 0, -89, -25, 4, 101, -114, -2, 81, 46, -15, 104, 127, 62, 26, 70, 37, 69, -68, 97, 52, -78, -125, -1, 67, 41, 4, 107, 61, -60, 21, -66, 27, 19, -44, 49, -69, -53, 26, -21, 8, -53, -124, 88, 9, -14, -53, -73, -41, 48, -77, 4, -44, 39, -115, -2, 113, -64, -105, -125, 88, -74, -25, -60, 35, 54, -1, -47, 121, -118, 67, 32, 50, 21, 60, -66, -19, -27, -79, 126, -122, -29, -47, 28, 62, 55, -123, 120, 37, 53, 81, 121, 51, -20, 38, 5, 80, 122, -6, -112, -82, -29, 105, 118, 118, 71, 66, 11, 37, -42, 59, -49, -105, 97, 73, -48, 44, -13, -78, 79, 93, 31, -33, 101, 111, -69, 70, -66, -84, -37, -91, 51, -111, -46, -114, -12, -60, 34, 49, -115, 32, -12, 96, -1, -16, 30, 22, 97, 59, -38, -6, -95, -28, -92, 5, -126, -46, -34, 43, 110, 49, 42, -17, -60, 61, -11, -7, 13, -77, 126, 86, -24, -79, -32, -87, -102, -119, -27, 41, -127, 119, -47, -87, -105, 45, -34, -108, -3, 124, 102, -128, 100, -6, -51, -44, -80, -2, 93, -91, -115, 50, -103, 80, 108, -23, -31, -33, 5, -40, 113, 111, 56, -74, -106, -39, -102, -78, 24, -39, -42, -102, 120, -8, 92, -85, -46, -81, 81, -66, -26, -28, 24, 33, 100, -27, -34, -119, 7, 86, 86, -24, 35, -121, -26, -1, -50, -48, 49, 93, 3, -30, -118, -96, -106, 18, -70, 109, 3, 100, 23, 88, -67, 111, -34, -82, 35, 104, 85, -127, 50, 71, 117, 56, 93, -8, -93, -88, 119, 16, 68, 106, -66, 68, -38, -126, 17, -83, -116, -87, -7, 0, 28, -35, -4, -110, -112, 0, -30, 62, -89, -100, 53, 49, 49, 33, 21, 119, 118, 124, 10, -82, 20, -100, 109, 86, -5, 96, 68, -89, -54, 0, 90, 19, 58, 58, 103, -8, 124, 23, -88, 96, 74, -60, 121, 62, -111, 124, 97, 65, 122, -53, -24, -107, -28, 38, 70, 112, -115, 108, -98, 120, -83, 74, -75, -39, -67, -103, 100, 85, 25, -118, 57, -123, 124, 115, -87, -89, -92, 70, 75, -121, -116, 36, 118, -115, -117, 98, 89, -45, 73, -7, -80, -71, -84, -12, 98, -14, -126, -35, -78, 53, -58, 122, -46, -14, -114, -115, 52, -21, -37, -38, -30, -78, 22, -124, 62, 65, 39, -1, -21, -44, -17, -92, -23, 26, 118, -123, 15, -121, 14, 61, -15, -7, -74, -11, -24, -8, -12, 2, -105, 24, -27, -15, 45, -11, 52, 41, -82, -47, -70, 44, 126, 114, -18, -83, -54, -122, -118, -110, 71, -70, -72, 107, -4, 2, -23, 116, 15, -90, 73, -118, 39, 1, 47, 84, -92, 16, 26, -98, 47, 28, -25, 91, 77, -33, -89, 2, 127, 64, 98, 59, -126, 10, -19, -65, -106, 12, -122, -4, 110, -20, 72, -125, 37, 32, 68, 53, 42, 110, 28, -112, 80, 40, 117, -8, 10, -94, 18, -13, 97, -48, 71, 121, -44, -118, -26, 94, 8, -59, -75, -5, -44, 101, 12, -81, 51, -85, -55, 118, 51, -94, 60, -126, -119, -61, 6, 79, 5, 82, -110, 5, 6, 31, 48, -21, 85, 23, -108, -69, -14, -45, 12, 65, 96, 6, 37, 43, 35, 119, 97, 11, -67, 53, 63, 104, 35, 68, -10, 74, 125, -21, 22, 25, 78, 61, -95, -103, 103, -2, 71, 124, 80, -46, 64, 0, 122, -37, -69, 125, 58, 118, 70, 33, -120, 127, 57, 59, 86, 85, -25, -94, -43, 79, -38, 60, 1, 53, 87, -112, 1, -5, 15, 42, -77, 38, 84, 43, -92, 14, 14, -77, 83, 9, -96, -66, -4, 91, -65, -64, -84, 98, 71, 66, 101, -72, -83, 48, 24, 60, 78, -77, -19, -81, -110, 63, 120, 79, 112, -97, -61, -20, -95, 59, 116, -110, -40, 48, 75, -97, -108, 54, 28, -104, 125, -7, -9, -3, -44, -18, 49, 6, -49, 118, -124, -97, 16, 8, -75, 3, 99, -53, -93, -60, -21, 36, -45, 63, -46, 120, -42, 16, 63, -79, -3, -93, 89, -117, -12, -116, -32, -76, 9, 100, -35, -93, -52, -97, -73, -105, 93, -100, 79, -31, 25, -100, -113, 83, 96, -51, -1, 0, 83, 50, -67, -57, 127, 105, -19, -25, 87, 36, -42, -103, -97, -20, -48, 19, 78, -125, 103, 67, 20, -24, -78, -118, -2, 97, -28, 5, -35, -65, -128, -56, -99, 125, -121, -25, 23, -41, -32, -84, 6, 41, -128, -16, -24, 25, -13, -103, 67, -122, -73, -46, 1, 46, -78, -32, 124, -69, -128, 15, -41, 124, 41, 35, 40, 26, 109, -6, 14, 55, 33, 10, 58, -93, -102, -105, -56, 57, 13, -19, 52, 65, 90, 64, -33, 56, -30, 116, 91, 32, 98, 102, -69, -13, -54, -15, 87, 19, 119, 54, 60, -35, 0, 24, -41, 86, 25, -87, 53, -107, 76, 32, -52, 88, 30, 91, -47, 110, -84, -115, -88, 102, -7, 29, 22, 17, -60, -81, -6, 99, -99, -69, -53, 109, -7, -21, -30, -98, -81, -54, 9, -75, 101, 126, -33, -29, -110, 61, -33, 77, 83, -123, -117, 66, 22, -47, -95, 54, -86, -97, 109, -35, -122, -94, 22, 64, 86, -66, -91, -78, 4, 95, 79, 99, 55, -125, -60, -119, -33, -10, -71, 121, 88, 26, -64, -30, -14, 111, -27, 115, -3, 16, -28, 46, 19, -75, -104, -113, 14, 14, -1, -83, -125, -111, 8, -65, -34, 34, 4, 88, 120, 19, 83, 82, -112, -12, 26, 89, -34, 8, 16, 54, -34, -125, 90, -49, 0, 55, -18, 96, 112, 112, -31, -57, -121, -104, 109, 8, -91, -2, 30, 98, -13, 104, -16, 10, 13, -52, 13, -66, -57, -56, 121, 18, 8, 89, -13, -66, -25, 99, -45, -27, 89, 80, -108, 19, 75, 104, -55, 19, 71, -59, -96, 30, -61, -122, 76, 89, -124, 30, 13, -97, 117, -57, -99, -95, 53, -114, -92, -85, 82, -75, -114, -105, 66, -95, -51, -41, -42, 106, -15, 67, 119, -7, 24, -85, -59, 82, 6, -125, -29, 2, 46, -103, 73, -108, -100, -103, 67, -29, -1, 43, 24, 98, -38, 88, -3, -125, 23, -109, 102, 124, 121, 16, 35, 99, 60, 0, -27, 71, -69, 45, -115, 31, 9, 74, 117, 49, -128, 2, 7, 81, -22, -49, 125, 126, 94, -18, -89, 97, 91, -78, -29, -34, 60, -41, -4, 121, -74, -72, -75, -104, 66, -40, -27, 62, -99, 98, 114, -124, 44, 3, -93, 45, 67, -78, -49, -22, -8, 109, -85, -96, -59, 0, 74, 93, -64, 87, 112, 61, 125, 73, -127, 97, -101, 13, -120, -100, -81, -22, -123, 90, -70, -110, 21, -118, 123, 121, -62, -116, 5, 93, 78, -16, 79, -66, -124, 40, -13, -113, -55, 34, -57, -40, 72, -128, 71, 107, -21, -66, 5, -93, -95, -18, 65, 51, -39, -61, 119, 114, -76, -46, 64, -74, -14, 37, -23, -128, -18, -43, -117, 65, -43, -128, -64, 21, 106, 9, -33, 102, -18, 121, 74, 112, -116, 106, -29, -69, 15, 5, 127, -93, -69, -84, 49, 105, -104, -110, 91, 40, 54, -17, 104, -119, 102, 36, 99, -106, 102, 60, 52, -61, 33, -69, 115, -34, -94, 67, 40, -9, 4, 82, 113, -64, 0, 110, -82, -54, 78, 81, 49, 101, -21, -89, -117, 49, 102, 20, -61, 80, 71, 40, -11, -92, -23, -30, 79, 92, 114, 84, -7, -120, -63, -3, -114, -98, 34, 118, 96, -96, -68, 0, 120, -61, -81, 108, -115, 93, 106, -115, 69, 6, -2, -8, -74, 29, -91, 62, -53, -67, -85, -127, -109, 65, 103, -44, 83, 2, 25, 31, -119, -20, -32, -110, 82, 51, 70, 71, 12, -121, -31, -26, -93, 102, -28, -65, -108, 114, -67, 44, -53, -61, -95, -63, 77, -68, -7, -83, -10, -66, 125, 15, 64, -84, 82, -7, -103, -3, 72, -50, 48, -72, -123, 16, -78, 35, -123, 126, 25, -82, -87, 107, -15, -107, 71, -67, 14, 127, 116, -7, -86, 57, 56, 88, 104, -113, -57, -55, 28, -6, -74, -70, -16, 123, 23, 81, 1, 125, -14, 98, 106, -66, -12, -77, 29, 21, -52, 72, -11, 78, -123, -117, 93, -92, -31, -20, 39, 24, -6, 101, -15, -26, 68, 53, -61, -76, -16, -95, 38, -126, -96, 82, -33, -87, 26, 127, 38, -39, -74, -3, 21, -85, 32, 2, 37, -56, -72, 81, -6, -92, 56, -74, 16, -17, -82, 78, -6, 49, 108, -98, -36, 95, 87, 95, -58, 36, -116, -25, 52, 82, 2, 112, 16, 88, 39, -63, 40, -65, 18, -74, 106, 107, 65, -65, 32, -55, -5, -90, 13, 79, 117, -127, 122, -62, 0, -12, -4, -1, 58, 19, 123, 99, 105, 45, -108, -114, 60, -99, -46, 121, 107, -12, -56, -61, -28, 105, -35, -55, 56, 55, -112, 24, 9, 85, 111, -103, -6, 47, 45, -57, -124, 113, -14, -110, -7, -117, 126, 68, -6, -110, -26, -62, 12, 40, -79, -45, 62, 14, 81, -64, -29, -128, -37, 44, 100, -113, -125, -105, 48, 37, 41, 100, 17, 74, 113, -62, -37, -118, -113, -61, -119, -82, 31, 39, -52, -50, 127, -121, 15, 90, -124, 21, 2, 15, -95, -46, -85, 100, -12, 1, 93, -105, -87, -25, 104, -86, -121, 6, 79, -110, 119, -110, -40, 33, -102, 54, 85, -32, -99, -75, 15, 124, -6, 69, -69, 114, -74, -42, 97, -20, 38, -96, -123, 87, 9, -38, -57, 104, -55, 22, 59, -101, 10, 117, -13, -23, 42, -101, -63, -19, -74, -119, -117, 111, 49, -26, -49, 108, 47, -103, -78, -126, 98, -93, -80, 21, 47, -58, -85, -127, -124, 93, 5, -19, 108, -22, 54, -112, 7, -11, -21, 114, -75, -58, 117, 112, 127, -69, -119, 90, -107, 116, -36, -9, 124, 121, 98, 73, 13, -108, -23, -81, -30, 40, 113, 50, -39, 119, -51, 43, 5, -91, -44, 105, -32, 112, 29, 118, 97, -15, -39, 68, 26, -11, -111, -56, 63, 78, -50, 113, -117, -82, 85, -48, 29, 5, 66, 54, 48, 35, 26, 4, -87, -17, -101, -39, -103, -126, -38, 98, 80, 0, -74, 107, 112, 6, -117, 36, -28, -73, 93, 91, 80, 68, -17, -118, -83, 30, 86, -95, -48, -107, 86, 90, -108, 57, -12, -104, 18, 78, 18, -115, -7, -106, -108, 16, 39, 95, 11, 117, -46, -44, -77, 47, -119, 37, -96, 42, -42, 88, 120, 75, -30, 51, 66, -110, 87, 22, -34, -93, -43, 61, -69, 45, -53, 101, 54, -35, 17, 111, 21, -127, 87, -68, -52, 28, 38, 104, -104, -23, -109, 66, -127, -89, 68, -124, 120, 116, 91, 92, 56, 14, -17, 48, -58, -54, -95, -61, -104, 100, 30, 8, 86, 21, 50, 115, 117, 96, 6, -19, 124, -92, -63, -17, -105, -15, 114, 91, -85, -60, 63, -9, -18, 1, -35, -1, -66, -31, -60, 71, 100, -32, 10, 114, -68, 52, 55, -100, 3, -46, -76, -123, -100, 92, -65, -87, 60, -120, 77, -104, -114, 61, -49, 6, 48, 105, 88, -43, 50, 50, 55, 92, 116, -69, -110, -72, -61, 111, -116, 124, 16, -60, -111, 14, -24, 73, -6, 13, 16, -125, 55, 26, -116, -26, -114, -56, -35, 12, 25, 74, -93, -110, -43, 70, -107, -114, 22, 72, 68, -98, 90, -12, -98, 101, -63, -104, -112, 29, 44, -2, -12, 93, -107, 114, 98, 83, -12, 72, 57, -63, 41, -33, 125, 91, -19, -96, -94, -66, -65, 77, 8, -114, -29, 80, -17, -109, -47, -31, -64, 0, 100, -107, -92, -1, -84, -30, -23, -46, 64, 87, -17, 126, 114, 98, 92, 20, -27, 14, -5, 57, 92, 6, -33, -39, 123, 31, 96, -69, -18, 67, 41, -32, -104, 61, 34, 8, 86, 102, 79, -105, -106, 47, 61, -54, -111, 19, -82, 65, -87, -113, 106, -50, 98, 4, 20, -68, 81, -60, -15, 87, -104, 87, -40, 46, 49, -65, -116, -33, 125, -57, -10, -35, 53, 79, 17, -10, -107, 42, -107, -73, 47, -13, 66, 95, 89, -49, -109, -71, -8, -42, 78, -3, 70, -34, -67, 101, 121, -101, -83, -122, 24, 84, 99, 2, -60, 42, -38, -98, 92, 42, -58, 116, -114, 119, 91, 127, -31, 42, 25, 60, -115, -110, -47, 57, -110, 77, 30, -104, -16, -32, 70, 26, 15, 0, -67, 59, -47, 81, -72, 3, 108, 90, 33, 62, -113, -98, 67, -17, 42, -48, -84, 42, -49, 37, 53, 63, 33, 78, -93, -66, -46, 127, -105, -51, 104, 34, -118, -39, -68, -13, -64, -93, 119, -1, -84, 42, 124, 47, 37, -37, 80, 89, 37, -93, -102, 40, 39, 76, -24, -115, -106, 113, -124, -19, 80, 78, -67, 10, -16, -99, 60, 57, -43, -85, -106, -37, -2, -44, 87, 22, -57, 64, -85, -8, 67, -97, 53, -127, -98, 73, -85, -114, 117, 71, 63, 1, -55, 29, 68, 61, 127, 30, 122, -80, -118, -54, -11, -26, 113, -107, 74, -81, 92, 9, 107, 38, 25, -49, -121, 21, 5, 85, 39, 124, -6, 49, 91, -62, -83, -92, -37, -43, -31, -83, -52, -117, 127, -73, -55, 100, 53, 47, 49, 0, -8, 114, 80, -60, -73, -103, -23, -120, 104, -108, -42, -120, -79, 11, -92, 119, 42, 27, 69, 104, -38, -111, 61, 83, -73, 101, 16, 108, 100, -77, -93, 25, -48, -42, -5, -66, -9, 98, -108, -39, -67, -34, -23, -116, 10, -104, 89, 108, 93, -16, -87, 124, -33, 105, -61, 60, -1, 45, 11, -27, 12, 86, 38, 125, 118, 19, 73, 108, -26, 35, -65, -84, -9, -50, -38, -87, -125, -121, 107, 32, 36, -111, 25, 60, -23, 69, -95, 1, 60, 28, -22, -32, -12, -10, 7, 70, 110, -104, 41, -87, 37, 93, -112, 91, 127, -56, -28, -20, 115, 30, 124, -5, 31, -109, -36, -57, 29, -88, 95, 61, -52, -53, -86, -4, 28, 115, 106, 53, -35, -121, -93, -15, 33, 8, 40, 58, 33, -56, -41, -83, 59, -46, 66, -115, -67, -81, 112, -90, -108, 89, -57, 40, 88, -92, 49, -73, 125, 34, 90, -17, -14, 121, 20, 26, 57, -35, -18, -58, 20, 116, 56, -79, 127, 96, 105, -52, 81, -63, 78, -121, 40, -53, -35, 95, -63, 52, 99, -53, 36, 117, 108, 57, 73, 115, -110, 57, -23, -84, 116, 23, 114, -73, -27, 69, -58, 110, 101, 84, -117, -19, 85, 55, -53, -34, 30, -48, 10, 11, -13, -66, 39, 74, 50, 126, 67, -126, -4, 42, 18, -17, 15, 6, -10, -6, -122, 118, 4, 50, 110, 40, 126, -118, -90, -106, 81, -44, 23, 58, -123, 115, 13, 49, 9, -49, -119, -69, 66, 82, 53, -2, 66, -8, 51, -65, -60, 11, -108, 35, 9, -37, 11, -27, -2, 105, 55, -6, -86, -20, -87, -82, 21, -85, 14, -72, -112, 65, 47, 96, 56, 7, -62, -36, -68, -112, -75, -27, 92, 2, 42, -64, -67, -29, 37, 68, 78, 116, -70, 93, -29, 77, 12, 124, -98, 63, -39, 92, 55, 121, -1, 107, 89, -23, -76, -45, 85, -109, 67, -38, -88, 52, 69, -90, 1, -84, 70, -41, -21, 29, 96, -112, 76, 30, -92, 32, 12, -47, 109, 91, 2, 81, -16, 78, -126, -97, 102, 9, -117, -110, -120, -65, 97, 27, 56, -89, 38, -93, 72, -6, 21, 61, 96, -36, -89, -105, -57, 18, 25, 27, 8, -41, -106, 107, 118, 49, -127, -3, 78, -121, 59, 3, -34, -9, -77, -18, -124, 27, 58, 116, -54, 106, -46, 27, -44, 50, 117, -74, 69, -92, -14, -14, -77, -20, 35, 105, 60, -80, 53, 96, 63, -97, 9, 90, -9, 96, 62, 112, -2, 56, -34, 43, -11, 102, -105, -114, -64, 107, 25, 74, -17, 17, 106, -104, -47, 67, -12, -92, 67, 9, 35, -119, -95, -94, -124, -102, 91, 83, -106, 26, 112, -54, 70, -17, -71, -81, -97, -70, -19, -115, 121, -22, -35, -63, 121, 70, -12, -29, -110, 55, -49, 83, 73, -20, -8, -33, 22, -18, 61, 27, 56, -84, -42, -35, 66, 46, -44, -61, -15, 76, -83, -13, -80, -66, 12, -103, -56, -93, 71, 58, 16, -102, -35, -29, -30, -110, 73, -15, -117, 100, 83, 11, 37, -91, 23, -32, 88, -123, -123, 24, 93, -65, -90, 57, 4, -41, -64, 38, -5, 78, -5, 121, 21, 31, 25, 30, 34, 1, -32, -50, -104, -96, 59, -75, 59, -105, -13, 110, 127, -7, 68, -92, -53, 105, 126, 72, -103, 66, 19, -24, -43, -116, -70, 106, 51, 89, -75, 12, 101, 119, -1, 109, 51, -105, 123, -6, -10, -18, -80, 15, -29, -2, -79, 88, -62, 55, 41, -2, 46, 0, -13, 44, 6, 33, 97, -118, -113, -9, -124, 24, 116, 6, 94, 110, 66, 39, -50, -73, 39, -85, -102, 62, -57, 7, -50, -9, -103, -33, -121, 102, -23, 43, 117, -28, -87, -40, 95, 106, 0, -106, 107, -29, 95, 70, 89, 92, 106, 35, 103, -16, 98, 44, 12, -2, -10, -37, -98, -25, 36, 14, -54, -6, -69, -67, 59, -111, 76, 54, -75, -30, 55, 60, -117, -66, -86, -1, 13, -83, 68, -95, -13, -10, -104, -10, 44, 64, 25, -55, -10, 78, -26, 77, 126, 103, 116, -43, 107, -20, 66, 48, -27, 77, -64, 73, -16, -66, -64, 35, 23, -65, 52, -19, 93, -45, -49, 37, -57, 92, -55, -108, 45, -38, 115, -56, -107, -7, 21, 57, -14, -11, 0, -84, -70, 70, -108, 127, 9, -87, -8, -28, -66, 33, -20, -113, -26, -1, 45, -36, 87, -3, 47, 48, 37, -117, -94, -63, 10, -112, 93, 120, 41, -32, -114, 65, 80, -63, -80, 36, 50, -85, 65, -22, -93, -34, 46, 123, -22, -29, -79, 61, 17, -70, 62, 64, 39, -23, -34, -26, 110, -17, 111, -71, -53, -62, -123, -69, -20, 57, 77, 23, -12, -69, -11, -26, 113, 107, -102, -55, 14, -78, -85, -118, 107, -35, 40, 112, 23, -127, 14, 77, -42, -17, -106, -88, 32, -24, -125, -9, 114, 30, 127, 28, -115, -104, -20, 123, -37, 23, -86, -12, -77, -36, -15, 23, -66, -14, 57, 62, 122, -49, 46, -24, -127, -95, -110, 4, -95, -16, 45, 55, 119, -118, 83, 1, -62, -50, -7, -24, 31, 105, -27, -42, 9, 56, 111, 123, -95, 115, -34, 59, -4, 123, 86, -98, -16, -117, 20, -45, -109, -25, 99, 105, -115, -125, -61, -89, -57, -1, 21, 8, -83, -43, -110, 39, -90, 67, 30, 113, -5, -36, 126, 54, 108, -64, -21, -76, -69, -126, -21, 99, 38, -23, 12, 108, 35, -32, -14, 91, -124, 12, 110, -102, -122, 85, 30, -73, -59, 50, 124, -120, 102, -122, -23, 42, -29, 70, -98, -43, -2, -100, 24, 44, 99, 14, -4, 27, 106, 109, -48, 21, -111, -5, 24, -39, -107, 2, 95, 93, -105, -109, 41, 1, -53, -7, -45, -106, -98, 90, 87, 48, -4, -38, 66, 24, -87, 32, -30, 55, 116, 84, 32, 52, 86, -53, 33, -22, 125, -13, 89, -4, 57, 14, 86, -111, 19, 96, 51, 53, 94, -1, -19, 48, 71, -25, 107, 126, 28, 29, -73, 73, 41, -13, -94, -22, -55, 65, 60, 12, -128, 14, 83, 42, 114, -82, -73, 26, 117, -17, -14, -5, 69, -33, 84, 76, -7, 104, 82, -1, 33, -42, 87, -72, 29, -47, -62, -57, 112, 95, 57, -61, 39, -88, 90, -50, 14, 39, 97, -51, 94, 2, -112, -105, -40, -110, 6, -63, 35, -93, 32, -66, -34, 69, -70, 5, 33, -77, 124, 43, -127, -11, 58, 71, -6, -2, -68, -95, -105, -67, -3, 91, 7, -120, 21, 60, 101, 123, -87, 8, 112, 4, 88, -117, 12, -89, -57, -84, -44, -30, 62, 37, 59, 23, 2, 16, -35, -36, 27, -68, -19, 35, -122, -46, 62, -53, 89, 7, 127, 106, 100, 37, 31, -34, -48, 75, -13, -27, 96, -59, 15, -73, 63, -10, 58, -62, -85, 86, 15, 8, -99, -50, 105, 20, -79, -102, -57, -63, -66, 32, 39, -94, 24, 39, -77, 124, 91, -47, 8, 19, 100, 74, -121, -95, -122, -101, 82, 17, 58, 116, -43, -49, -72, -28, 77, -55, -103, -22, -61, -29, -26, 60, 45, -52, 93, 4, 103, 6, -118, 53, 75, -62, -66, -45, -91, -112, 26, 62, 46, 71, -36, -124, -127, -24, 44, -108, -58, 98, 14, 37, 27, -72, 9, -50, -118, -117, -14, 100, 64, -44, 18, 110, -92, -54, -78, 17, -44, -104, 114, -78, -42, 65, -105, -54, 43, 123, 77, -94, 85, 55, -101, 107, -127, 123, -80, 116, -79, -103, -18, -82, -22, -46, 43, -1, 33, 22, 75, -104, 3, 78, 76, -126, -103, -60, 119, -89, 97, 17, -108, 86, 52, 40, 33, -69, -69, 60, -53, 58, -119, -43, -97, -123, 25, 12, 47, 87, -60, 53, -81, 111, 39, -38, 123, 44, 18, -123, 28, -2, 115, 89, 80, 20, 122, -7, -67, -75, -1, 5, 32, -48, 103, 106, 101, -24, 28, 67, 42, 30, 108, 34, 96, 122, 20, 24, -70, -14, 2, 58, -46, 7, 88, -56, -43, -56, -32, -94, -93, 91, 20, 27, 101, -72, -93, -59, 27, -60, 100, 65, -24, -116, 19, -45, -63, 70, 88, -21, 5, 12, -61, 93, 83, -103, 21, -71, -76, 7, -54, -39, -47, -112, 41, 95, 93, -40, -51, -45, 124, 26, 74, 46, -84, -62, -116, -80, 14, 118, 46, 90, -32, 51, 119, 6, -14, 55, 51, -126, -75, -87, -86, -29, 87, 0, -7, 85, -104, 12, -20, 107, -4, 58, 113, -6, -43, -98, 91, 116, -125, 0, -3, 47, -47, -88, 81, -103, 90, 14, -45, -86, 114, 38, 69, 62, 71, 60, 86, 103, 30, -81, -44, -83, -107, -119, -68, 92, 74, 16, -48, -17, 34, -42, -84, -44, -24, -33, 122, 35, -22, -48, -101, 23, 72, 68, -65, -126, -54, -20, -90, -113, 70, -104, 120, 76, -93, 81, 58, -15, 122, -16, 29, 126, -6, 92, -67, 88, -7, 68, 126, 45, -60, 33, -105, -36, 107, 27, -38, 50, 106, 27, -37, 18, 118, -86, 59, -65, 20, 101, -67, 18, -91, -35, -109, 31, -55, -57, 66, 109, -9, -85, 17, 90, 58, 43, 106, -94, -45, -7, 37, -3, -83, -26, -112, -8, 72, 55, -3, -106, 8, -114, -28, -88, 45, -24, 18, -19, -59, -14, 53, -37, 13, -36, 118, -108, 14, -92, -23, 32, -115, 90, -13, -104, -117, 23, -56, 75, -48, 11, -2, -48, 96, 59, 76, 32, 72, -48, -46, -24, -100, 41, 84, -9, 54, -74, 41, 111, 112, -128, 60, 28, -90, -59, -71, 58, -9, -113, 91, 88, 58, 72, -123, 50, -122, -124, -45, -51, -41, 82, -85, -23, 80, -16, 8, -80, 88, -74, 120, -61, 91, -7, -112, -6, 14, -86, -8, 108, 122, 84, -123, 1, -24, 70, 42, -1, -104, 116, 77, -113, 3, 36, 123, 69, -36, -96, -55, 104, -34, 89, -93, -2, -10, -93, -34, -125, -11, -13, 93, -119, 49, 0, 16, 101, 74, 79, -82, 71, 107, -66, -100, -3, -22, -63, -14, 88, -120, 94, 60, -10, 82, 61, 106, -49, 32, 6, -111, 66, -32, -108, -88, -11, -119, -101, 89, 52, -110, -128, -118, 0, 92, 7, -20, -13, 32, -122, 86, -101, -128, 32, 83, -126, -32, -109, -47, 12, 86, -63, 106, 120, 89, 113, 66, -90, 35, -75, 95, 115, 48, -41, 105, 123, 20, 38, -110, -40, 89, -75, -111, -122, 105, -60, 103, -102, 100, -77, -48, 119, 5, -89, -120, -14, -26, -45, 45, -107, -83, 88, 69, -2, -79, -64, 40, -77, 58, 125, -127, -80, -34, 26, 95, 93, 50, -102, 31, 86, -122, -12, -105, -118, 104, -124, 31, 61, 8, 0, -73, -42, -44, -91, 87, 115, 59, 59, -127, 61, 80, -6, -119, 11, 104, 40, 78, 89, -9, -112, -27, 57, 103, -54, 88, 45, 103, 18, -73, 113, -93, 14, 41, 45, -55, 97, 3, -1, 106, 76, 20, 40, -128, -97, -46, 94, -123, -25, -69, -33, 83, -95, 40, -117, 18, -35, 67, -98, -9, -12, -52, 39, 114, -27, 11, 45, -70, 30, -25, 106, -50, -119, 23, -85, 118, 61, 80, -35, 33, -98, -16, 89, 0, -107, 119, 58, 24, 71, -21, 25, 82, 87, -72, 14, 67, -109, -31, 103, 92, -59, 25, 56, 92, -81, -38, 71, -90, -38, -35, 57, -66, -24, 77, -76, -111, -95, -88, -119, 36, -69, 37, 100, 38, 29, -45, 38, -49, -82, 40, 63, -20, 89, 93, 39, -124, -71, -62, -118, 44, -8, -11, -89, -54, 8, -24, 118, -4, -101, 121, 29, -82, -100, -119, -76, -26, 30, 124, 55, 76, -53, 28, 60, 51, -100, 75, 80, -48, -86, 90, -45, 41, 0, -30, -1, 21, 15, 51, 93, -16, 85, -107, -1, 83, -9, 67, 70, -89, -93, 86, 78, -92, 105, -38, -76, -87, 124, -42, 67, -103, -51, 88, 47, 34, 19, 9, -66, 115, -94, 106, 42, -18, -6, -53, -27, 69, -125, -111, -12, 12, 15, 2, -115, 59, 55, -96, 13, 97, 32, 90, -115, 18, -43, -77, 80, 76, 45, -50, 116, -100, 45, 88, 68, 24, 83, 72, -27, -56, -49, -1, -44, 77, -99, -108, -102, 7, 4, -98, -18, -57, 65, -124, 5, 54, 120, -5, 34, 122, -2, -1, 125, -57, 41, -23, 102, 46, -93, -21, 86, -22, -94, 4, 9, 125, 0, -7, 62, -110, -82, -3, -112, -33, 94, -96, 71, 80, -119, 48, -91, 92, -10, 111, 68, -35, 119, -71, -10, -119, -15, 117, -100, -58, 123, -50, -57, -88, 109, -56, -94, -11, -50, 122, 77, 118, 96, -58, -30, -48, -80, 71, 25, 36, 80, 9, -112, 47, 30, 97, -113, 80, 21, -24, 83, -90, 60, 33, 6, 102, 117, 103, -120, -9, 113, -91, 118, 76, 103, 11, 63, 18, 97, -85, -109, -91, 4, 47, 58, 107, 83, 105, -63, -19, -22, -90, 8, -43, -35, -56, 64, -104, -91, -87, 91, -66, -5, 71, -23, -102, 45, 8, -32, -44, 123, -101, 83, -120, 16, -25, 44, 69, 125, -90, 79, -93, -44, -37, -18, -116, 123, -33, -43, 109, -33, -38, -91, 40, 1, -33, -100, -81, -63, -53, 96, 29, 122, 122, -125, 49, -34, -111, 123, -39, 120, 8, 42, 65, -67, -83, -34, 76, 109, -41, 2, -92, -120, 120, -121, 6, -38, -124, -29, -59, 115, 66, -87, 11, -110, -121, 109, 20, -45, -33, -74, 84, -77, 3, -15, -82, -45, 112, -122, 87, -38, 50, -21, 87, 44, 54, -118, -15, 104, 66, 16, 91, 22, -39, 12, -111, -83, -24, -82, 89, 49, -112, -28, 71, -12, -113, -82, 15, 7, 104, 107, 29, 90, 30, -17, -30, 33, 43, -79, -128, -34, -27, -87, -13, 24, -93, -19, -44, 69, 89, 76, -32, 61, 94, -37, -47, 24, 11, 124, -102, -44, -48, 110, 61, 5, -82, 20, -126, 77, 122, -37, -103, -118, 52, -78, 115, -40, -127, -75, 98, 89, -111, -64, 120, 63, 10, 29, -31, 48, 78, 123, 111, -27, -72, 18, -14, 54, 119, -114, -5, -43, 63, -125, -46, -39, 7, 16, -5, 36, 121, 96, -67, 17, -88, -107, -106, -106, -125, -47, -65, 12, -107, 96, -101, 126, -97, 77, 74, 67, 73, -101, -97, 112, -118, -89, -17, 102, 100, 68, 91, -24, 94, 67, 44, -125, 55, -96, -63, -51, -118, -82, -4, 41, -28, -95, -8, -92, -46, -100, -90, 109, 54, 121, -48, -123, 18, 97, -104, 81, -89, -92, 59, -100, 81, -13, 89, 126, 67, -23, 62, 15, -23, 112, 14, 3, -16, 84, -127, 85, 89, -28, -72, 99, 101, 105, -88, 103, -110, 60, 52, 61, -85, 11, -22, 89, 49, -89, 66, -12, -100, 75, -88, -124, 115, -2, 107, -2, 100, 97, 91, 92, -43, -87, 81, -17, 118, -88, -114, -22, 51, 44, 104, 43, 39, 100, -84, -80, 112, 62, -106, -64, -102, -86, 70, 58, 92, -66, -69, -78, -26, 46, 87, 82, 112, 63, -51, -39, 16, 83, -92, -78, 118, -120, 78, -35, -28, 27, -1, -44, -117, 92, 40, 121, -30, 117, -86, 8, 28, -127, 42, -101, 124, 113, -86, 92, 40, 16, 88, -57, -7, 77, 77, -104, 42, -91, 43, 103, -11, 39, -127, 16, 11, 84, -60, 35, 42, -24, 2, -10, -98, 122, 102, -94, 108, -53, -74, 31, 15, 118, 50, 56, -18, -2, 109, 75, -62, -49, -49, 104, 64, 59, 21, 98, -107, 105, 21, -104, -31, 47, 23, 106, -47, 124, 93, -89, 53, 5, 92, 95, -97, -68, 67, 34, -89, 127, -23, 59, -128, 98, -63, -71, -74, -125, 28, -63, 65, 71, 40, 80, -5, -113, -96, -10, -22, -30, -40, 105, 100, -10, -80, 95, 80, 111, 96, -48, 25, 4, 112, -117, 6, 4, 6, -91, -109, 22, -1, 92, -60, -71, 84, -32, -24, -61, 17, 113, -35, -35, 52, 63, -87, -74, -103, 122, -89, 68, -37, 61, 8, 0, -102, 96, 4, -35, 23, -47, -92, 72, -29, -47, -33, 104, -82, 97, 91, -109, -26, 3, 55, 17, -12, -25, -4, -108, 10, -83, -87, 22, 69, -63, -5, 37, 77, -82, -103, 44, -80, -24, -8, 21, -66, 120, 40, -50, 25, -87, 12, -114, -1, -41, 32, -106, -96, -95, 19, 90, -103, 100, -124, 126, 18, -67, 68, -88, 29, -8, 0, 16, -79, 69, -97, -90, -117, -128, -35, 42, -99, 68, 8, 124, -105, 15, 29, 104, -106, 116, -48, 24, 51, -73, -118, 14, 27, -13, -95, 116, 39, 42, 78, -96, -41, 36, 81, 104, 95, 112, -2, -20, 102, -34, -80, 126, -78, 30, -70, -80, -63, 45, 49, -102, 13, -34, -81, -79, -85, -27, 88, -86, 112, -108, -115, -46, -29, 10, 87, -31, -46, -39, -92, -64, 28, 39, 8, -31, 112, -91, 116, -118, -48, 64, -81, 37, -10, 39, -77, 90, 112, -60, -63, 107, -8, -125, 3, 116, 90, -13, 70, -62, -7, -59, 91, -36, -52, -15, -29, -124, -19, -54, -85, 111, 89, 24, 11, 10, -19, -101, -22, 102, -8, 118, -79, -105, -37, 22, 64, 36, 118, 111, 66, 108, -36, 47, 16, 39, 26, -43, 112, 65, -18, 102, -29, -116, -108, 120, 109, -112, -82, -74, 99, -69, -64, -46, -93, 31, 50, -25, 76, -115, 5, -58, 110, 72, 61, -63, 98, 55, 106, 10, 44, 30, -92, 5, -12, 63, 37, -41, 107, -52, 79, -107, 115, 30, -71, -121, -101, 46, 15, 32, 41, 64, 5, -57, 116, 81, 19, 85, 106, 120, 1, 69, -23, -37, -76, -49, 92, 5, 117, -82, -68, 32, 57, -4, -37, 73, 125, 20, 116, 52, -123, -26, -70, 52, -39, -106, -18, -72, -74, 43, -109, 8, 67, 69, 56, 42, 104, 47, 63, -27, -21, 93, -98, 83, 112, 27, -2, -21, 26, -57, -72, -8, 92, 70, 71, 49, 111, -46, 31, -38, 101, 12, 38, -12, -26, 97, -102, -58, 115, 123, -18, 78, 0, 98, -77, 108, 59, 118, 67, 64, 123, -52, -1, 15, -8, -61, -89, -67, -56, -90, -83, 109, -115, 111, -83, 87, -67, 2, -5, -27, 1, -60, 67, 93, -80, 112, 91, 4, -82, -80, 58, -115, 103, 127, 123, 52, -116, 93, 9, 40, -39, -58, -19, 108, 39, -64, -49, 88, 31, -63, 110, 28, 104, 113, -55, 84, 76, 49, -7, -17, 5, -45, 5, -86, -99, -15, 63, 3, -128, -7, -5, 79, -38, 59, 58, 68, 58, -68, -69, 8, 61, -7, -39, -1, 74, 76, 39, 100, 94, -90, -85, -85, -80, -29, -97, 103, 105, -21, 7, -105, -42, 108, -5, 71, -49, 11, 2, -121, -88, 113, 23, -89, -45, -49, -80, -44, -89, 118, -114, -97, 19, -123, 88, 60, -105, 71, -92, 120, 101, 43, -40, 70, -38, 40, 77, -61, -57, -105, 90, -39, 64, -86, -3, 46, -22, -76, 106, 89, 113, 60, -128, -16, -30, 83, -97, -28, 55, 9, 124, -28, 101, 110, -67, -13, -76, -1, -73, 22, -51, 107, -100, -68, 52, 42, -33, 58, 65, -33, -61, -79, 71, -75, -116, -16, 33, 51, -5, 76, -74, 10, -125, -111, 22, 58, 9, -24, 78, -74, -3, -106, -80, -90, -67, 71, -97, -90, -93, -72, 117, 95, 113, -41, 32, 53, 100, -70, -19, -91, -65, -125, 38, -1, -66, -55, 16, 101, -27, 16, -108, -37, -55, -127, 74, 110, 108, -19, 27, -32, 2, -71, 19, -26, -26, 50, 12, -76, 100, -6, 0, -104, -13, -115, 50, 57, 114, 14, 117, -93, 117, 83, 39, -5, 78, -26, -29, 95, -80, -96, -30, -99, 98, 59, -60, 11, -112, 118, -84, -128, -5, -114, -52, -114, -105, -112, -71, 122, -115, -86, -46, 69, -47, -23, 90, -93, 80, -43, -39, -64, 30, 55, -107, -32, -78, -37, 124, -16, -39, -58, 33, -122, -78, 3, 34, -32, -75, -3, 39, 115, 6, -109, -109, 122, 121, -104, -77, -16, -42, -109, -66, 125, 113, -116, -103, -98, -16, 10, 9, 110, 19, -34, -69, -57, -124, 91, 80, 27, 100, 48, -109, -125, -49, -11, -2, 37, -45, 78, 43, 81, 10, -110, -14, 59, -58, 13, -113, 65, -32, 27, 105, 46, -36, -108, -5, -13, 32, 1, -85, 82, -116, 80, -90, -8, 83, -74, 29, 91, -86, -101, 49, -100, 17, 21, 61, -24, 91, -59, -14, 84, -57, -26, 113, 94, 80, -72, -96, -18, -59, -119, -11, -6, 27, 14, -76, 15, -15, 15, 102, -41, -10, -77, -10, 108, 6, -35, -83, -38, 24, -5, 18, 24, 32, -8, 124, 25, -37, 69, 5, -76, 30, -52, 5, 93, -63, -29, 69, 82, 100, -22, 98, 109, 96, -89, 38, -41, 93, -113, 45, -12, 125, 84, -72, -100, 49, 67, -54, 8, -26, 113, -19, -51, -124, 20, -72, -55, 5, -49, -46, 79, -62, -80, 39, -88, 82, 42, -64, -101, 93, -11, 98, -18, 122, 122, 105, -106, -21, -21, -97, 121, -20, -15, -62, -57, 4, -105, -87, 9, -47, -5, 102, 59, -110, -46, 83, -107, 27, -2, -67, 44, 7, 82, -113, -115, -71, 25, 33, 110, 109, -82, -3, 7, 104, -96, -27, 68, 23, -117, 83, -125, 61, -90, 12, 21, -125, 92, 19, -45, 76, 67, 56, -55, 57, 12, -70, 5, -43, -96, -62, -107, -11, -105, -23, 43, -9, -99, -111, -26, 9, 58, 55, 50, 48, 33, 76, -120, -124, 69, -109, 69, 101, 88, 33, 72, -116, 4, 121, -126, -86, -101, -19, -118, 118, 12, -118, 77, 56, 98, 8, 29, -86, 3, 126, 89, 64, 116, -89, 33, 84, -25, -4, 40, 61, -70, 94, 105, 101, 58, 36, -124, 115, 88, -81, 124, 13, -23, -40, -119, 106, -90, 63, -3, -20, -31, -69, -107, 44, 4, 76, -15, -73, 125, -19, 120, 79, 123, 31, -110, 102, -87, 38, 94, -34, 36, 48, -73, 9, 56, -94, 99, 97, -125, -106, -105, -17, -118, -44, 116, -127, 112, 43, -25, -81, -109, -84, 86, -2, -69, -65, 63, -43, -95, 127, -75, 118, 70, 57, -94, 64, 36, 7, -105, -102, -15, -62, -83, -70, 84, -37, 27, 88, -68, -95, -63, -68, 59, 76, 35, -60, -89, 87, 17, -83, 10, 115, -25, 1, 33, -3, 2, -50, -46, 4, 34, -123, 65, -59, -49, -37, -120, 40, -10, -68, 9, 44, -122, -93, 57, -63, -9, -48, -43, -99, 11, 79, -64, 58, 77, -50, -3, -127, 45, 67, 66, 61, 45, 12, 122, 60, -78, 37, 96, -76, 115, -7, -1, -49, 69, 104, -100, 105, 5, 61, -125, -110, -116, -106, -46, -91, -126, 118, -69, -78, 54, -100, 28, -104, 48, -77, 101, -95, -33, 69, -26, -105, 42, -56, -22, 37, 114, -49, 119, -14, 36, 107, 62, -78, 78, -58, -42, -46, -42, -128, -114, -128, -80, 50, -68, -94, 18, 65, -75, 35, 46, 40, 27, -61, 35, 127, 122, -101, 27, -121, 95, -47, 122, -53, -112, -88, 81, 100, 98, 40, 46, 60, 58, 73, 69, -31, 11, 109, -4, 54, 78, 117, 19, -81, 18, -119, -8, 99, -79, -39, 11, 40, 39, -84, 36, 9, -3, 27, -51, -8, 22, 116, -123, 4, 97, -98, -117, 20, -78, -82, -82, 100, -100, -94, -40, -121, -114, 26, -70, -77, 113, -60, -23, -7, 114, 63, 70, 74, 112, -112, 9, 5, -48, -30, 32, 2, -79, -23, -101, 118, -35, -31, 31, 97, 23, 78, 10, -33, -84, 48, -20, -23, -108, 88, -29, 126, 19, 113, -66, -123, -10, 30, 110, 22, -60, -44, 107, 56, 115, -23, -107, -32, -76, 23, 38, -104, -72, -6, 106, -10, 84, -37, -5, -22, 124, -83, -16, -7, -43, -4, 81, 22, 68, 44, 30, 48, 41, -122, -31, -104, -10, -126, 41, 113, 41, -25, 54, 87, -118, -73, 25, 64, -127, -75, -63, -107, 34, -17, -82, -113, 53, 15, -3, -35, -31, -22, -111, 113, 23, 26, 46, 74, 43, -46, -33, 7, 56, 81, 66, -4, -5, 90, -106, 120, -59, 33, -90, -26, -34, 42, -21, -84, -10, 114, 69, 118, -74, -71, -73, 114, 39, -108, -7, -67, 101, -84, -67, -80, 30, -76, 82, -15, 123, -82, 17, -120, 87, -108, -49, 32, 48, 113, 106, -69, 79, 59, -21, 53, 9, 110, 28, 21, -68, 100, 89, -24, 37, 21, -97, 19, 88, -128, -10, 92, -112, 1, 120, -60, 123, 58, -104, 95, -121, -44, 47, 55, -4, -83, 19, -18, 18, -104, 55, -56, 60, -46, 122, -79, 17, -74, 20, 120, 50, -118, -60, -85, 54, 30, -4, -54, -113, 12, 94, 15, 124, 83, 116, 110, -67, 113, -83, -92, -112, -106, -127, 85, -17, -11, 5, -92, -79, 36, -106, -58, 29, 97, 101, -77, 21, 89, -74, -107, 45, 26, -54, -40, 106, 118, 79, 60, -121, -59, 118, -98, 18, -119, -83, 21, -89, -95, 69, 116, 80, 42, 64, -38, 6, 1, 125, 33, 119, -38, -94, -104, 37, -50, 92, 41, -80, 121, -82, 49, 83, 127, -68, 38, -83, -54, 97, 93, -112, -3, -122, 47, -101, 100, 127, 70, 104, 19, 54, -50, -80, -28, 45, 126, -104, -14, 101, -91, -1, -98, 112, -110, -25, -47, -37, 60, -33, 73, 103, 38, -8, 83, -62, -96, 41, 78, -13, -92, -43, -56, -16, 31, -80, 72, 31, 42, -6, -12, 63, 18, -4, 104, 123, 26, 56, 63, -35, 44, 118, -80, 45, 58, 90, -75, 82, 112, -102, -67, -69, 60, 117, 33, 12, -28, -36, -121, 46, -62, -117, -89, 10, 120, -123, 41, 9, -23, 9, -27, -32, 36, -86, -102, 50, 17, -66, -89, 74, -70, -36, 78, -22, -16, 108, 65, -74, 24, 117, 101, 116, 21, -16, -43, 5, -57, -114, 102, -90, 61, 90, 20, 68, 21, -111, 88, -107, -8, 6, -37, -97, -125, 67, -75, -35, -105, -122, 120, -9, 119, 8, -74, -110, -91, 46, 73, -18, -128, 84, -120, 79, 16, 75, -22, -91, -13, -12, -47, -4, -106, 83, 25, 77, 35, -15, -23, -19, -16, -78, 107, -20, -67, -23, 15, 64, -116, 84, 107, -25, -3, -81, 85, -3, 79, -65, 56, 124, 100, 113, -124, -104, -6, -70, -110, 71, -120, 42, -89, 82, -6, 55, 73, 8, 28, 119, 43, 64, 71, -77, -53, 15, -102, 64, 61, 117, 52, 25, -33, -29, 58, 63, 62, 115, 75, -24, -127, 2, -37, 93, 65, 55, 125, 108, -79, 71, -116, -106, 48, -14, -123, -15, 40, 71, -114, 109, 39, 105, -65, 72, 11, -24, 99, 49, -104, -109, 65, -80, 68, -104, -70, 80, 30, -97, -51, 100, 65, -25, -51, 19, -53, -33, 109, 47, -82, 108, 26, 17, -110, 97, -74, 19, 34, 93, 59, 5, 115, 72, 89, -67, 19, 33, 74, -116, 75, -60, 114, -92, -13, -90, -27, -52, 8, 53, -105, 97, -57, -6, 100, -102, 82, 122, -109, -112, -60, -26, 90, 105, -110, 118, 127, 110, -126, -45, 48, -106, 45, 121, -61, 60, 32, 65, 30, -26, 85, 122, 52, 25, -23, 37, -90, -44, 107, 78, -26, 66, 72, -116, 20, 118, -71, -2, 105, 79, 27, -128, 39, 48, -72, 118, 119, 47, 117, -98, 87, 105, -69, 107, -46, 75, 72, -21, 123, -91, -63, 104, 19, 68, -103, -43, 31, 66, -115, 120, -87, -49, -85, 9, 59, 17, -74, -105, -83, -114, 74, -98, -99, -53, 50, 100, 84, -116, -89, 121, -45, -33, -78, 78, -99, -122, 73, 25, 114, 63, -106, 58, 32, -116, -101, 105, 23, 31, -96, -15, 89, -55, -35, -53, -122, 8, -69, 17, -64, 53, 45, 91, 52, -49, 49, -82, -39, 84, 121, 67, 45, -69, -90, 70, -80, -36, -15, -74, -43, 24, -111, 79, -120, -65, -47, 80, -17, 32, 125, -82, 109, -80, -10, 56, 11, 35, 66, 3, 51, 76, -82, 95, 20, 39, -66, 17, 123, -115, -115, 44, -28, -126, -7, -122, -110, 56, 88, 39, -38, 54, 104, 65, 56, -82, 47, -15, -57, -126, 17, -123, 6, 86, -44, -46, 78, 57, -51, -8, -21, 116, 12, -65, -98, 106, 30, -39, 53, 50, -44, -96, -108, 22, 78, -27, 92, 97, -71, 84, 32, 122, -68, -35, -112, -78, -112, -36, -74, -101, -52, 66, 120, 57, -42, 40, 77, 25, 90, 41, -70, -15, -67, 10, 41, -114, -103, -110, -54, 23, 26, 35, 114, 47, -42, -102, -85, 95, -56, 106, -49, 125, -13, 91, -105, 46, 65, 120, 98, -43, -67, -73, -43, -79, 70, -106, -2, -63, -39, 119, -13, -104, -70, -21, -117, 60, 77, 65, -22, 20, 96, 17, 45, 91, -59, 45, 44, -100, -48, -58, 34, -49, -43, 91, -97, 44, 106, 115, -19, -80, 80, 35, -96, 45, -89, 73, 41, -86, -87, -76, -95, 100, 22, 64, 97, -73, 22, 58, -62, 45, 57, -51, -63, 12, -8, 6, -8, -124, -80, -44, -118, 27, 33, -36, 28, -99, -58, 33, -26, 73, 15, 0, 99, -21, -61, -101, -8, -34, -119, 26, 75, 52, 80, 75, -33, 91, 108, -91, 78, -74, 38, 4, 12, -125, -36, -118, -24, 14, 123, -76, -94, 103, 48, 93, 12, 115, 25, -63, 64, 110, 85, 26, 112, 2, 124, 93, -79, 15, -70, 111, -77, -109, 125, 11, -80, 19, 6, -77, 39, 79, 20, 118, 122, -83, -102, 85, 119, -115, -126, 58, 34, -113, -18, 27, 76, -5, 77, 84, 73, -54, 9, 2, 82, 61, 98, 114, -59, 49, -22, 64, 2, -31, 11, -2, -23, -71, 123, 10, 107, 45, -98, 50, 25, -127, -114, 78, -26, 78, 28, 57, -45, 56, -110, -47, 24, -122, 44, -22, 11, 109, 70, 90, -122, 47, -122, 72, 57, 37, 125, -97, 55, 89, -95, -23, 62, -80, -58, 100, 93, -6, -35, 75, 51, -90, -48, -112, 40, -75, 60, 2, 1, -69, 66, -101, 49, 52, 67, -45, 81, -105, 111, 75, -99, 3, -53, -38, 127, 48, -34, 28, 126, 123, -116, 100, -69, 54, -86, 11, -13, -9, 73, -54, 103, -48, 78, -83, 31, 81, -24, 77, 68, 56, -60, -33, -16, 1, 126, -26, -119, -18, -16, -36, -74, -84, 57, -42, 64, 45, -16, -85, -88, 19, -90, -16, -10, -5, 88, 3, 79, 73, -113, -92, -114, 67, 36, 35, -7, -14, -57, 51, -78, 20, -86, -62, 73, 119, 44, 113, -80, -15, -124, -83, -66, -113, -59, -110, -29, 100, 93, -110, -47, 61, 89, -3, -31, -74, 3, 62, 118, -72, -21, 118, -64, -113, -118, 83, 5, -1, 52, -37, -57, -42, -68, -47, -101, 34, -72, -56, -84, -33, -97, -16, 21, -73, -72, -119, 69, -112, 127, -44, -119, -94, -19, 93, 32, -68, -22, 126, -35, 121, 91, -45, -48, -9, -128, -63, 55, 14, -62, -46, 23, 120, 122, 103, 4, -66, 47, -24, -120, 74, -116, -21, 38, 70, -69, -128, -54, -66, 98, -94, 58, -12, -30, 71, 28, 17, 29, 24, -45, 83, 84, 114, 69, 84, 49, 37, -71, 11, -76, -59, -119, 59, -25, -99, 64, 31, -64, -67, 110, -38, 2, 50, 74, -93, 48, 30, -106, -89, -8, -62, 71, 109, -106, -127, 118, 21, -112, 65, 45, -58, -55, -124, -62, -99, -52, -84, 111, -107, 36, 112, 1, 57, 14, -93, 27, -26, 8, -11, -26, -103, -83, 22, 52, -79, -14, -95, -124, -36, -57, 77, -89, 57, -106, -28, 126, -14, -9, 0, -16, -58, 54, -73, 87, 95, -23, 104, -33, -90, -100, 44, -73, -14, -51, -128, 47, 68, 112, 8, -117, -105, -70, -113, -32, 126, -76, 22, 28, -28, -26, -52, -23, -9, -122, 8, 49, -85, 91, 109, -50, 28, 62, 78, -70, 20, -115, -33, -74, 75, 120, 125, -32, 85, -103, 49, -55, -91, 14, -31, -19, -96, -37, 41, -97, 78, -83, -84, 74, -51, 122, 3, -70, -28, -115, -43, 4, 78, 125, -21, 42, -121, 123, -11, 61, 74, 13, -93, 19, -68, 26, -53, -106, 5, -77, -43, -24, -19, -12, 124, 26, 76, 20, 33, -65, 67, 59, -87, 29, -86, 97, -45, -51, 10, -8, -73, -83, -122, -7, -84, -69, -6, 49, -121, 53, 77, 31, -36, 24, 32, 55, 68, 126, -76, -125, 60, -37, -1, -46, 110, -91, 4, -17, 119, -16, 44, -67, 106, -59, 63, 89, -47, 100, -20, 107, -114, -37, 88, 103, -41, -76, -71, -117, -122, -108, 25, -121, -54, 123, -71, 101, -21, 13, -76, 108, 16, -71, 120, -32, -53, 6, -87, -95, 47, 58, -16, -27, 106, 122, -38, 102, 41, 87, -70, -65, 16, 28, -32, 0, -83, 86, -90, -128, 65, 55, 25, -55, 79, -27, 43, -4, 117, -54, 94, -48, 25, 43, 97, -45, -43, -120, -118, -14, -126, 103, -57, -114, -103, -87, 86, -54, -50, -32, -77, -27, -27, -109, 16, 97, -109, 2, 107, -29, -71, 121, 79, 91, 72, -66, -6, 24, 58, -24, -82, 65, -50, 97, 99, 109, -37, 108, -3, -114, -2, 63, 98, 24, -60, -50, -38, -16, 89, -100, -1, -72, -67, 73, -112, -73, -58, -40, -39, -28, -60, 114, -90, -104, -101, -52, -21, 54, -81, 71, -30, -84, 122, -86, 28, 43, 28, -45, -17, 93, -16, 36, -7, 60, 42, -101, 36, 95, 72, -60, -35, -41, 119, -123, -101, -24, 107, 31, -77, 4, 98, -78, 104, -75, 6, -50, -2, 97, 119, -78, 53, -104, -113, -9, -79, 51, -123, 96, 19, 95, 106, -45, -64, -115, -15, -97, 42, -63, -66, 100, 83, 106, 82, -65, -15, 42, -107, 105, -82, -76, 34, 87, 19, -93, 124, 75, 68, 4, 37, 72, 117, -66, -31, 15, -119, 33, -38, 123, -27, -84, 77, -61, 123, -56, 64, -61, -96, 88, -56, -20, 14, 53, -31, 67, -37, -53, -2, 42, -94, -12, -6, -62, -97, 29, 4, 48, -23, 97, -49, 84, -21, 86, -66, -74, 120, -67, 96, 98, 18, -9, -66, 15, -74, 1, 83, -107, -48, -48, 117, 120, -50, 65, -94, 108, 43, 65, 110, 108, 100, 8, 19, 35, 94, -77, -39, 124, -4, 6, -31, -58, 78, -88, 37, -104, -94, -87, -2, -82, -126, 43, -40, -90, 68, -62, -116, -73, -40, 107, -21, -89, -51, 47, 26, -58, -5, -12, -117, 5, 55, -91, -89, -77, 21, 109, -33, 122, 96, -37, 126, 14, 11, -12, -94, -60, -128, -83, 55, -22, 1, 43, -5, 110, -77, -63, 126, 54, -30, -121, 106, 114, -52, 47, -128, -66, -117, -79, 68, 4, -27, -93, -34, 45, -47, -18, -117, -17, -69, -91, 11, 127, 18, -100, 104, -77, -9, -12, -93, -94, -47, 116, -113, 41, -11, 67, -100, 114, 21, 101, -78, -128, -72, 96, -11, -31, -120, 127, 113, -91, 62, -26, -81, -109, -82, -12, -18, -122, 37, 66, -119, 73, 0, -108, -27, 41, 104, 0, 125, 54, -114, -37, 65, -102, -53, 34, 90, 116, -60, -33, -110, 77, 82, 17, 60, -105, 122, -6, 58, -121, 90, -59, -105, 127, 126, 83, -93, -22, -23, 104, 87, -60, 87, 52, 127, 120, 47, -73, 33, 87, 55, -103, 123, 89, -30, -18, -89, 65, -64, 11, 6, -87, -45, 81, -124, 31, -16, 90, -26, 77, 90, -9, -28, 36, -65, -12, -108, 26, -128, 36, -29, -12, 58, 107, -123, -59, 53, -92, 72, -57, -27, 99, -80, -81, 7, -6, 84, 21, -107, -67, 81, 45, 70, 15, 18, -21, 43, 46, -108, -15, -10, -116, -15, 57, 1, 72, -50, -108, 25, -8, -120, 60, 41, 68, 125, -83, -73, -121, -75, -47, 124, -46, -3, 65, 118, 55, -55, -51, 120, 55, 65, -79, 83, 96, -97, 18, 10, 77, -59, 105, -31, 108, -106, -49, 2, -120, 65, -58, 19, 117, -104, 31, -111, 17, 19, 113, -65, 59, -91, 109, -77, -65, 79, -63, -54, -119, -96, 64, -45, -78, 5, 102, 13, 54, -21, 78, -118, -34, 51, 20, 57, -10, 72, -39, -70, -34, 87, -66, -13, -44, -123, -1, -76, -40, -54, 27, 46, 116, -99, -97, 106, 125, 104, 10, -18, 26, 68, 1, -51, 40, 92, 27, 63, 99, 59, -50, 13, -37, -67, 15, -83, 111, 113, -14, -41, 10, -51, -115, -102, 103, 92, 112, -118, -59, -19, 0, -47, -121, -84, -48, 18, -42, -86, 109, 16, 71, -46, -71, -41, -118, -87, 114, 14, 31, -97, -24, 67, -89, 54, -97, -126, 33, 25, -92, -120, -83, -61, 72, -114, 5, -74, -108, -45, -15, 57, 4, 22, 81, 123, -21, -103, 50, 90, -45, 80, 66, -35, 125, -110, 73, 38, -31, -74, -101, 28, -43, 12, 104, -125, -65, -77, 123, 57, 46, 87, 101, 49, 57, 99, 7, 53, 95, -112, 10, -107, -125, 117, 15, -83, -104, 25, 121, 78, -121, -105, 125, 77, -86, 10, 59, 32, 123, -101, 104, -56, -4, 114, -5, -97, 104, -43, 77, -40, -33, 110, -22, -79, 47, 3, 51, 86, -88, -1, -105, -75, -18, -8, 54, 119, -49, -77, 122, 67, 53, 57, -3, 1, 84, 119, 111, 33, 80, 44, 45, -15, 91, 36, -117, 103, 101, -15, 38, 89, -114, -56, 126, 111, 39, -7, -123, -21, 42, 1, 91, 85, 62, -92, 70, -89, -78, -44, -94, -106, -87, 23, -116, 1, 17, 47, 54, -48, -14, -20, -6, -53, 8, -3, -66, 88, 13, 13, -33, -77, -55, 22, -95, 74, -82, 35, 122, -57, -13, -105, -127, -6, -115, -54, -121, 78, -94, 36, 112, 1, 75, 58, 15, -121, 6, -60, -121, -50, 30, 101, -13, -113, 6, 88, -120, -16, -42, 37, 21, -69, 98, -44, -91, 61, 111, -48, 99, 25, 111, 95, 70, 21, -23, 52, 16, -95, 72, -57, -121, -8, 17, -116, 91, -39, 111, 59, -42, 10, 113, 68, 74, 50, 108, 11, 63, -115, 116, 35, 21, 59, -6, 100, 77, 48, 46, -126, -48, -10, 72, 48, -8, -82, -10, 97, -98, 118, 66, -112, -32, 74, -103, -78, -14, 65, -45, 91, -63, -13, -122, -77, 86, -110, -67, -120, 36, -57, 95, 115, 111, 11, 93, -106, 123, -115, -102, -69, 84, 108, -39, -125, -50, -108, 93, 29, 53, 19, 120, 112, 87, -32, 100, 125, 101, -11, 84, -49, 84, 86, 108, 84, 3, -90, 21, 122, -57, -123, -13, 21, 31, -4, 38, 77, -103, 56, 61, 105, -37, 12, -32, -34, -62, 69, 7, -85, -87, 82, 56, 39, -3, -46, 1, -95, -61, -24, -19, 82, 108, 112, 102, -11, 63, -74, -58, 122, 27, 50, -106, -91, 23, 86, 113, 13, 11, 89, 41, 67, 66, -63, -92, -28, 43, 70, -80, 94, -114, -60, 117, 119, -120, 105, -107, 69, -14, -70, -33, 22, -64, -75, 113, -87, 112, -125, 53, 103, 30, 68, 28, 13, 109, -111, 67, 82, -50, 16, -55, -128, 67, 35, 72, 47, 41, -5, -84, -115, -38, 105, 79, -84, -37, 51, -5, -45, -2, 104, 12, 9, 34, -64, 91, 99, -15, 4, 127, 92, -32, -105, 69, 70, -7, -98, 127, 5, -124, 81, -35, 124, 14, 74, 28, -110, -17, -79, 116, -53, -80, -99, -79, -7, 12, -95, -6, -119, 56, 80, -120, -84, 36, 114, -109, -128, 61, 61, -29, 22, -58, 15, 49, 19, 13, -72, 80, -20, 99, 2, 19, 107, -105, 51, -96, -62, 66, 38, 101, 112, -51, 66, -71, -47, -19, -67, 8, 26, -33, -103, 59, -55, 34, 126, 60, -78, 121, 52, -11, -116, -88, 57, -116, 91, -13, 63, -112, -14, -54, -31, -75, 35, -47, 95, -98, -115, 46, -30, -80, 59, 64, -11, -54, -71, -31, 125, 73, 16, 37, -7, 117, -56, -118, -69, -109, -44, 74, -116, 22, -49, -11, -55, 22, -9, -21, 54, 52, -98, 78, -38, 126, 101, 95, -2, -77, 78, -128, 57, 13, -25, 106, -104, 37, 84, 84, 33, -61, 103, 37, 79, -77, -51, 34, 103, 112, -17, 51, -105, -64, 71, 2, 28, -37, -112, 98, 127, -124, -62, 10, 123, 0, 71, -28, -58, 17, -113, 7, 11, -110, -67, 59, 38, 103, -61, 104, 24, -43, 5, -21, 11, -117, -128, 5, 59, -72, 40, 40, -3, -81, -66, 51, 19, -115, -46, 70, -117, 38, 73, -6, 64, -98, 65, -34, 104, 98, -8, 80, 67, -84, 12, 101, 101, -91, 44, -74, -92, -48, 45, -103, -92, -71, -52, -87, 126, -73, 41, -71, 22, -92, 48, -48, -102, 64, 21, -47, -85, -67, 45, -97, 85, 29, 86, -1, 96, -21, -83, 115, -48, 23, 72, -119, -110, 117, -57, -2, -109, -55, 50, -43, 123, 120, -18, 93, -121, -22, -51, 31, 119, 21, -60, -120, -80, 70, -87, -56, -127, -77, -91, 100, 88, 101, -31, 77, 10, -73, -39, -15, 80, 112, 39, 31, 22, 84, -123, -64, 61, 76, 47, 36, -47, 29, 82, -113, -86, -8, -36, -110, 8, 111, -29, 2, -16, 52, -91, 27, -30, -98, 17, 39, -50, 63, -11, -106, 66, 121, -34, -82, 127, -1, -54, 80, 117, 95, -1, -72, 124, -92, 80, 1, -79, -58, -109, -20, -102, -117, -95, -82, -108, -7, 119, -9, -122, -84, -39, -76, -124, -64, -51, 64, -84, 108, 30, 60, 78, 63, -114, 42, 41, -127, -71, 21, -117, -125, -59, 58, 23, -46, -119, 56, 103, 7, 55, 28, 30, 62, 53, 123, -67, 82, -29, 123, -46, 82, -68, 93, 90, 115, 127, 66, 1, -120, -77, -99, -84, 84, -37, 121, 43, -89, -94, 96, 88, -82, -43, 16, -35, -102, -35, 46, 97, 12, -40, -126, 0, -19, -41, 7, 21, -78, 115, 115, -106, 69, -118, -24, 105, 111, -79, 7, -27, 28, 117, -34, -46, 85, -29, 91, -4, -80, 101, -94, 101, 118, 113, 17, 68, -113, 70, -100, 66, -81, -126, -7, 61, 12, -99, 48, 48, -42, -116, -81, -125, 11, 4, 50, 62, 118, -63, -17, 63, 122, -38, 102, 95, 2, -41, 80, 14, -42, 57, 43, -31, 107, -21, 77, -16, -45, 10, -78, -48, -34, 62, 36, 12, -74, -13, -48, -58, 7, 48, -61, -4, -71, 36, 108, 104, -46, -90, -98, 18, -33, 111, 93, 74, -120, -23, 38, 96, 97, -123, -71, -108, -48, -104, -96, -67, 23, -116, -4, 82, -56, -73, -7, -114, -49, -17, -103, -20, -31, 91, 117, -102, 6, -39, 38, -117, -89, 3, 13, -75, -96, 50, 118, 51, -59, -93, -79, -56, -101, -97, -16, 75, 8, 83, 63, 122, 116, -109, -43, 37, 105, -128, 13, 16, 52, 97, 62, -28, -43, 103, -76, 43, -60, -9, 56, -61, 44, 53, -7, 17, 15, -11, 96, -94, 73, 77, 11, -17, 94, -30, 86, -27, 29, 124, 18, -34, 20, -4, 107, 66, 75, -84, -22, -58, -14, 57, -118, 118, 19, 10, -75, -124, 61, -95, 82, -114, -100, 13, -111, 50, 39, 54, 16, 83, 116, -71, -5, -120, -49, -110, -76, 68, 83, -77, 59, -55, -16, 109, 58, -101, -50, -45, -91, 51, 91, -59, 29, 85, 55, -126, 41, 105, -49, -23, 93, -36, 32, -112, 21, 77, -100, 37, -63, 110, 116, -104, -70, 94, 63, -58, -47, 93, 104, -30, 8, -29, -80, 35, -102, 15, 85, -102, 97, -37, 25, 127, 4, -63, 117, -125, 106, -75, -113, -107, 1, 53, 65, -100, 114, -28, 14, 25, -6, 104, 38, -77, -64, -34, -4, 107, -28, -14, -126, -89, -52, -106, -3, 8, 114, 119, -108, -109, 42, 14, 75, 91, -107, -27, 119, -87, -12, -91, 101, -48, -18, 56, -46, -80, -119, -61, 113, -92, -39, -38, -104, 60, 57, 39, -92, 104, -103, 21, -85, -61, -105, 80, -27, 26, -44, -19, 84, 53, -16, -50, 55, 85, -10, -122, 73, 125, 123, -119, -110, -76, -41, 109, -64, -81, -33, 106, 59, -119, 4, -6, -13, -69, 77, 117, 67, -46, -35, 81, 113, -49, -61, 127, -39, 52, 117, -45, 11, 62, 81, 6, -107, -10, 29, -49, -30, 57, -98, -95, 36, -72, 27, -25, 121, -111, 123, 66, 124, 19, 114, -16, -79, -108, -16, -44, -116, 86, -3, -108, -106, -65, 27, 45, -37, -55, 3, -57, -2, -109, -57, 11, 68, -56, -30, 44, 11, -99, -105, 97, 7, -72, 92, -22, 120, -78, -13, 126, 112, 30, -118, 93, -36, 29, -55, 33, 69, -84, -104, 9, -83, 106, 39, -60, 22, 48, -71, 127, 25, 83, 69, -106, 43, 2, -127, 0, -68, -46, 1, 17, 109, -109, 104, 124, -90, 98, 70, -75, -57, 93, -29, 91, -58, 38, 12, 91, -68, -76, 73, 23, 93, -12, -86, -18, 77, 42, 85, -34, -118, -77, -44, -128, 31, -38, 20, 58, -92, -113, 19, -120, -59, 44, 34, -89, 55, -34, 18, 3, 87, -4, 111, 106, 37, 81, 5, -116, -60, -9, 24, -54, -25, 88, 49, -81, 49, 95, -2, 23, 4, 125, -63, -3, -69, 43, -28, 78, 46, -98, 39, -3, -27, 35, 87, 0, 17, -108, -8, -35, 52, 102, 35, -34, 86, 16, -23, 19, -46, -26, 110, 124, -106, -95, 28, -14, -34, 65, 89, -45, -71, -111, -104, -59, -104, 42, -75, -91, -53, 93, -125, -30, -34, -19, -88, -108, -64, 53, -37, -111, -103, 56, 24, -50, 30, -13, -19, 1, 101, 29, -15, 43, -29, -70, -30, 87, -93, -53, 52, 20, -90, 122, 79, -21, 121, -55, 100, 103, 80, -96, -35, -89, 55, 14, 123, -91, -5, 89, 12, 101, 67, 85, -103, -32, -92, -18, -37, 111, -104, -52, -33, -72, -67, -121, -1, 103, -18, 71, -100, -49, -58, -103, 52, -64, 82, 19, 57, 107, -96, 10, 124, -84, -117, 45, 48, 62, 93, 111, 58, -47, -10, 67, -64, 108, 68, 58, 16, 57, -2, 93, 24, 60, -109, -103, 95, -11, -125, 70, 88, 58, -121, -27, 16, -126, -36, -118, 52, 91, -81, -30, 7, 26, 84, -108, 94, -50, 102, 99, 57, 15, -117, 105, 69, 21, -94, -120, 116, 50, 44, 61, -29, 119, -89, -109, -91, 110, -44, 115, -38, 23, 24, -113, 85, 75, -25, -58, -104, 51, -74, 67, -66, 96, 39, -28, 69, 37, -51, -12, 76, 14, 96, -17, 30, -113, -121, -93, -117, -6, -109, -50, 17, 7, 40, 48, -17, 124, 127, -71, 47, -44, -39, 109, -62, -66, 123, -35, -58, 71, 62, -37, 105, -71, -100, -5, 124, 60, -54, 107, -106, 40, 29, 83, 25, 2, 122, 123, -110, -21, -69, 51, 81, -114, -55, -118, 79, 35, -61, -11, 73, -119, -84, 6, -27, 87, -34, -52, 47, -75, 16, -72, 35, 27, 61, -24, 28, -4, 38, -6, -119, -109, -122, -121, -83, 118, 122, 10, 49, 7, 90, -50, 119, 26, -116, -59, 107, -96, 78, 125, 62, -22, -52, -60, 37, 16, -36, -49, -97, -74, 75, -65, -97, 12, -23, 60, 124, 116, -82, -117, 76, -128, 115, -98, 47, 58, -94, 100, 46, -95, -76, 44, -11, 16, -77, 15, -69, -116, 24, 68, 88, -97, -4, -48, 47, -67, 74, 49, 39, 103, -118, 1, 77, 108, 111, -126, -48, -41, -42, 14, 68, -109, 59, -89, 71, -114, -21, 2, -71, 2, -2, -27, 2, -68, -30, -18, -2, 127, -122, 86, -85, 94, -82, -79, 76, 22, 98, 59, 51, -71, 104, 29, -125, 22, -77, 92, -78, 124, -85, -99, 7, -94, 55, 70, 125, 22, -108, 16, 31, -99, 65, 58, 100, 97, -63, -21, 39, -33, -15, 49, -85, 92, 33, -123, 119, 16, -38, 118, -51, 109, -115, -13, 125, -108, -32, 64, 24, -40, 88, 95, 116, 108, -26, -14, 90, -47, -1, 64, 58, 38, 109, -56, 71, 50, 23, 76, 91, -71, 70, 11, 67, -27, -127, 81, 124, -1, -97, 117, 60, 6, 44, 85, 50, -56, -14, -57, 73, -110, -36, 67, 117, -118, 41, 27, 85, 51, -55, 36, -4, -87, 42, 47, 118, -45, 3, 103, 41, -90, 122, -14, -51, 55, -29, 52, 111, 23, 64, 68, -11, 65, 72, -23, -68, 51, -125, -107, 110, 87, -43, 76, -77, -85, -86, -58, 98, -25, 46, 67, 45, 77, -49, -117, 11, -59, 25, -127, 36, 58, 96, -30, 40, 108, -86, -57, 121, -63, -85, 125, -77, 117, 65, 126, -112, -112, -128, -80, 119, -91, -42, -81, 108, -88, -96, -100, -86, 124, 94, 113, -94, -51, 98, 81, -101, 108, -60, -41, -59, 98, -62, 59, 87, -46, -76, -116, -33, -98, 110, 18, -39, -39, 90, 7, 113, 14, -26, 89, 13, -4, 34, -101, -121, 112, -122, -37, 54, 87, -92, 68, -68, 46, 72, -101, 61, 48, -98, -47, -100, -6, -46, 92, 114, -35, 36, 121, 95, -72, -21, 94, 122, -12, 36, 64, -114, 76, 26, 126, 30, 75, -66, -126, 104, -90, -40, 34, 114, -100, 54, 91, 33, 91, -32, 35, -27, 32, 63, -28, -53, -35, 10, 46, 50, -23, 70, -25, 75, -116, -15, 55, 109, 65, -98, -118, -105, -93, 111, 49, -3, -115, -68, 54, 101, 101, -99, 16, 83, 114, -117, 106, -16, 109, -112, 104, -98, -103, 14, 5, -111, 84, 19, -35, 68, -123, -73, -63, 127, 99, -24, -23, -29, 25, 97, 121, -74, -17, -92, 34, 43, -31, -122, 99, -23, 25, 51, 72, -119, -30, 28, 75, -58, -55, -93, -3, 112, 108, 86, 51, -65, 63, -39, 19, 121, -110, 63, -128, 100, 55, 17, -102, -124, 62, -102, 122, 16, 36, 102, -119, 77, -16, -119, -41, 124, 12, 126, 40, 14, -30, -61, -7, 110, 77, -108, -12, -111, 125, 52, 99, -23, 67, -12, 11, 22, -127, -5, 43, 79, 64, 31, -4, 109, 54, 70, -99, 112, 80, -63, -69, -60, 88, 35, -119, -95, -110, 98, 106, 108, 126, -17, -30, -127, -62, 47, 32, 126, -50, -51, -58, 48, -122, 53, 85, -5, -100, 66, 41, -126, -72, -60, 59, -118, 35, -116, -126, -10, 116, 53, 42, -122, -109, -32, -104, -95, -21, -34, -62, -25, -8, 69, 98, -37, -118, -88, -27, 97, -124, -43, -37, 75, -48, 56, -27, -57, 55, -64, 14, -14, 75, 65, -69, 100, 106, -56, 115, -30, 111, 53, 43, 74, 34, 45, 84, -31, -86, 99, 63, 119, 7, -13, 1, 127, -55, -69, 35, -8, 4, 11, -101, -62, -12, -74, 81, -48, -24, -75, -61, 27, -17, -92, -96, -21, -34, -18, -81, -58, -70, 15, 61, 61, -108, -99, 15, 41, -77, -126, 59, -17, 20, 115, -10, -123, -120, 107, 15, -30, 39, 34, -100, -86, -103, -28, -99, 124, -91, 116, 61, -51, 75, -127, 95, -27, -62, -128, 89, 32, -110, -78, -111, 42, 61, 52, -119, 13, 60, -6, -107, -4, 118, -70, -111, -59, -37, -28, -53, 3, 103, -58, -118, -90, 118, 96, -126, 25, -110, 7, -57, -57, -11, -44, 125, 50, -116, -116, 40, 21, 106, 45, -35, 30, -26, -79, 61, 101, -97, 32, -105, -20, -124, -92, -53, 4, -32, 83, 53, 59, 126, 96, 61, -109, -112, 13, -24, -44, 87, 63, -65, -76, 13, 69, -114, -85, -109, -35, -98, -25, 65, 96, -50, 11, 61, -106, -81, 97, -32, 37, -85, 54, 43, 81, 31, -98, -58, 29, 101, 69, -86, 85, 61, 66, -102, -114, -86, -47, 107, 63, -68, 77, 21, -80, 15, -32, 23, -91, 0, 109, 12, 101, 3, -8, -16, -41, -36, 12, -119, -100, 127, -124, -51, 90, -17, -100, -110, 23, -91, -2, -118, 102, 84, -17, -127, 69, -72, 55, -67, -6, 55, -34, -11, -68, -12, 87, 88, 78, -67, -16, 106, -18, 31, -116, -99, -19, -101, 102, 37, -47, 22, 108, 45, -75, 58, -78, 66, 28, -111, -51, 27, -41, -30, -103, -41, 66, -110, -85, -83, 75, 13, 35, 39, 106, 32, 55, 119, -12, -93, -70, -62, 80, -92, -102, -62, -85, -38, 62, 86, -105, -1, -83, 30, -54, -44, -127, -20, -90, -46, -105, -22, -110, 8, -27, 97, -108, -82, 65, 75, 95, 3, 127, -21, 85, 35, -110, -122, 20, -74, 10, -8, -62, -96, -22, -15, -117, 10, -125, 26, -38, 110, -119, -77, 60, 25, 101, 53, -126, 92, -40, -84, 97, -11, 97, -83, -72, 46, 35, 51, 52, -47, 102, -72, 115, 42, -21, -121, -13, -57, -87, -99, 35, -115, -20, -73, -67, 6, -91, -22, -22, 108, -10, 77, -39, 62, 107, 78, -76, -27, -27, -27, 4, -67, -31, -69, 52, -120, -53, 52, 56, 66, 103, 26, -33, -14, 0, -108, -89, 76, -90, 119, -25, 36, 47, -89, 78, 102, 107, 106, 103, 66, 2, 54, -109, 63, 74, -22, 109, 97, -101, 49, -60, -126, -51, -87, 5, -123, -108, -80, -9, -100, 97, -124, 84, 36, -68, -99, 78, 124, -18, 111, -44, 98, -110, 45, -103, -1, 79, 37, 10, -93, 55, -124, -32, -79, -73, 85, -32, 58, 14, 52, -27, -88, -79, -60, 45, -117, -63, -11, -13, 33, -95, 90, -52, 56, 119, 27, -13, 68, -125, -53, -4, -35, 41, 33, 99, 5, -14, -65, 123, 66, 63, -38, -41, -45, 104, -24, -48, -73, 51, 33, 3, -79, -53, 106, -71, -43, 19, 81, 101, -97, 18, 68, -113, 80, -75, -128, -111, -8, -110, -22, 55, -2, -112, -46, -17, -50, -24, -54, 112, -95, 99, 23, 17, 80, 59, 59, -66, -44, -24, -77, 106, -37, 22, -88, -76, 101, 93, -43, -84, 44, 25, 55, -10, -112, -87, 34, 12, 100, -75, -89, 21, 126, 78, -66, 75, -8, 82, -12, -2, 41, -94, 92, -17, 82, -93, 64, 97, 90, -124, 106, 32, 18, 71, 20, -109, 61, -127, 16, 48, 16, 82, 54, 81, 93, -94, -100, 8, 36, 34, 51, 101, -98, -81, -124, -123, -78, 26, 32, 23, -20, 67, 92, -114, 110, 104, -108, 112, -40, -87, -88, 49, 70, 102, 8, 123, 49, 43, -91, -91, -112, 44, 5, -63, -117, 115, 85, -57, 40, -41, -28, -105, -96, -42, -127, 85, -110, 32, 15, -11, -8, 100, -99, 36, 100, 81, 105, -23, -10, -15, -30, 126, -101, 76, 57, 87, 47, -45, -57, -83, -17, 113, -9, -108, 103, 5, -22, 21, -69, 50, 92, 46, 77, -47, 25, -106, -49, 57, 49, -51, 1, -121, 73, 4, 1, -51, 99, 111, -98, 99, -93, -67, -120, 9, -68, 37, 71, -84, 0, -78, 37, -34, -54, -85, 16, 72, -64, -32, -43, 7, 105, 2, 61, -38, 9, -51, 57, -124, 36, -60, 69, 32, 3, -55, 84, 62, 47, 45, -30, -118, 48, -9, -76, 33, -84, -81, -27, 125, 23, 83, 79, -128, -35, -31, -17, -95, -1, 57, -22, 15, -65, 113, 17, -45, 121, -91, -22, 94, 73, 46, 56, -54, -60, 13, 79, 39, -10, 88, 2, 89, 67, -60, 118, 53, 107, 102, -68, 110, -15, -117, 82, 23, -67, -94, -114, 60, -82, -69, 87, 122, 47, 99, -124, 82, -35, -104, 101, -85, 91, -60, 68, 40, 8, 77, -12, -3, -78, -43, -7, 24, -9, -67, -90, -111, 87, 64, -83, 125, -13, -78, 84, -113, -99, 10, -87, -33, -43, 121, -17, -102, -7, 31, -20, -105, 30, 29, -38, 33, 60, 67, 85, 60, 34, 77, 104, 10, -87, 36, 84, -9, 31, 23, 107, 48, -33, 46, 99, -96, -72, 25, -16, 16, 33, 43, 36, 126, 4, 68, 8, 35, 75, 29, 66, 23, 3, -126, -83, -72, 51, 70, 107, -33, -23, -8, -109, -3, 111, -126, -107, -7, -104, 78, -105, 56, -92, 26, -9, -120, -116, 104, 116, -29, 28, -5, 113, 45, -63, -56, -82, 28, -9, -109, 117, 5, -82, 67, -64, -39, -92, -46, -15, 68, -43, 52, -8, -8, -120, 48, 96, 89, 33, -112, -70, -92, -127, 109, 116, -34, -95, 108, 87, 29, 37, -50, -38, -8, -123, -49, 113, -39, 105, -96, -14, -76, -47, 87, 77, 84, -76, 78, 111, 33, -117, 78, -57, -1, -6, 92, 52, 9, 84, 45, 109, 95, -89, 73, -78, 24, 39, 56, -127, -37, -26, -65, 105, -68, -121, -102, 38, 16, -46, 91, -62, -72, -43, -44, 45, -94, -3, -68, -75, -128, 61, -69, -118, -92, 10, 52, 67, 122, 53, 91, 1, 107, 78, 47, 14, -81, -68, 110, 88, 22, -119, 58, -127, -109, 86, -88, 22, 56, 60, 65, 56, 88, -3, -41, 77, 63, 125, -65, 126, -61, -124, -15, 9, 112, 26, 93, -35, -119, -87, 66, -13, -5, -92, -87, -69, 19, 74, 118, 50, -48, 77, -5, 83, -102, -5, 105, 6, -124, -74, 15, 62, -90, -47, -35, -7, 3, -110, -11, 64, 116, -46, -79, -117, 58, -32, 1, 101, -57, -40, 56, -2, 52, 91, -121, -126, 105, -62, -34, -91, -54, 98, 29, -78, 85, -118, -89, 44, -78, 46, 74, 26, -9, -79, -62, -115, -43, 82, -123, -47, 17, -44, -54, 25, -123, -88, 98, 37, 83, 108, -12, 47, -8, 0, -40, -90, -36, -17, -103, 9, -41, 51, 77, -92, -104, -18, 82, 0, -125, -124, -26, 126, -2, -123, 23, 18, -114, -44, 94, -34, -46, -41, 14, 122, -10, 104, 86, -26, -55, 53, 83, -27, 52, -38, -108, 40, 7, 33, 24, -11, -86, 66, -103, -4, 58, 102, -39, 116, 49, -37, 123, -117, -10, 88, -122, 57, -33, 70, 31, -15, -12, 1, 60, -120, 72, -27, -56, -36, -98, -78, -49, -81, 120, 88, -21, -44, -55, -64, -88, 85, -83, -114, 95, 61, 27, -63, -120, -127, -7, 114, -52, -20, -32, -94, 23, 62, -55, -110, -56, -103, -87, 98, -52, 82, 116, -65, 82, 108, 4, 125, 103, -68, -15, 12, 0, 71, 32, -11, -123, -61, 55, -29, 80, -68, 78, 69, -75, 80, 32, -73, -84, -119, 51, 24, 94, 124, 69, -44, -7, -119, 66, 31, 65, 101, 72, 111, -39, -78, 75, -45, -62, 103, 70, 70, -8, -58, -76, 44, 13, 109, -68, -84, -3, -96, 24, 27, 10, -128, 6, -41, -2, 22, -81, -44, 108, -57, 8, 17, 40, 116, 19, -89, 8, 46, -85, -77, 102, 25, -97, 70, -99, 44, -86, 88, -96, 8, -94, 56, -94, 91, -64, 106, 67, -52, -14, -92, 58, -55, -24, -31, 88, -20, -110, 126, 1, 64, -25, 20, 2, 94, -35, -40, -53, -13, -104, -109, -109, -18, 82, -118, 104, 96, 75, -91, -39, 39, -118, 12, -3, -76, 62, -54, -120, -30, 93, 78, -53, 77, -124, -5, -121, 109, 64, 13, 118, -68, 56, 127, 12, 60, -32, 7, -62, -65, 7, 52, -20, -107, 80, -60, 61, 17, 94, -25, -18, 12, 54, 21, -104, -84, 73, -42, 61, 60, -53, -35, -19, -103, -21, 118, -43, -42, -18, -48, 84, -2, 4, 13, -116, 7, -109, -52, -63, -60, 30, -112, 110, -115, 89, 71, -100, 52, -33, 124, 36, 36, 48, -113, -101, -50, 41, 69, -112, 117, 90, -112, -93, -75, 9, -10, -125, -115, 59, 6, -65, 80, 44, -100, 78, -116, 45, -103, -46, -24, 45, 14, 55, 32, 76, 82, -8, -99, 33, -26, -4, 42, 107, 57, -92, -99, -66, 40, 126, -102, 74, 124, -34, -67, 109, 112, 5, 57, -62, -47, -1, -40, -124, -20, 17, -61, -105, 87, -56, -1, -61, -94, 60, 115, -86, 106, 39, -36, -51, 26, -114, 41, 65, -108, 68, 49, -67, -11, 81, -52, 65, -46, -45, -74, -4, 99, 80, 88, 55, 90, -51, -49, 0, -12, 17, 33, -98, -20, -127, -127, 122, -6, 93, -45, 61, -30, -128, 102, 36, 73, 95, -10, 113, -98, -33, -109, 23, -12, 75, -33, -104, 9, 110, 93, -106, 33, -29, -114, 11, -55, -8, 120, -9, -10, -108, 114, -63, 83, -58, 24, 28, 9, -24, 85, -114, 76, 26, -9, 100, 74, 11, 103, -74, 19, 81, -59, -61, -59, -88, -83, -124, 30, -123, 122, 43, -16, -46, 95, 90, 124, 41, 51, -89, -114, 22, -127, 30, 109, -3, -55, 87, -91, 111, 89, 77, 90, -116, 17, -51, -97, -70, 91, -9, -123, -22, -109, -119, 74, 40, -100, 9, -45, 72, -34, 27, -56, 95, 125, -35, -93, -28, 100, 35, -12, 126, 83, 56, 43, -38, 111, -32, -89, 28, 87, 100, 17, 119, -22, -4, -20, -42, -27, -116, -63, 119, 27, 37, -125, 84, 50, -9, 64, -64, 10, -36, -40, 56, 6, 26, -44, 33, -59, 81, -127, 71, -119, 24, 119, 117, -66, 76, -98, 77, 77, 88, -78, -27, 87, -76, 41, -41, -128, 50, 110, 55, -94, 74, 89, -123, -74, -52, 96, 17, 72, -45, -11, -46, -20, 27, -34, -13, -4, 68, -108, 29, 52, 113, 94, -72, -115, 7, -104, -32, -17, 28, 84, -74, -108, 79, 111, -42, -32, -121, 49, 0, 68, -107, 8, 59, 4, -93, -43, 97, 41, 121, 125, 70, -70, -53, 124, 87, 19, -55, 109, -35, 107, 13, -89, -12, 18, 95, -15, -123, -70, -24, -90, 95, -117, 4, 60, 114, 108, -84, -93, -8, -27, 88, 73, -60, -100, 11, -62, 82, 110, 43, -41, 10, -62, -11, -122, 65, 117, 10, -81, -96, -4, -112, -88, 86, -83, 89, -51, -116, -97, -90, -41, 80, -106, -81, 43, -89, 41, 125, 70, -91, -102, -48, 6, 12, 31, -51, -71, 72, -103, -100, 68, 58, 127, -63, 31, -25, -24, 88, -124, 112, 38, 10, 88, 61, -75, -33, 67, -126, -19, -112, -106, 122, -88, 18, 106, 6, -32, -32, -50, -128, 126, 118, -16, 79, -69, -73, -118, 72, 20, 105, -35, -102, -86, 119, 13, 66, 53, -70, 117, -109, -37, 40, -54, 51, -20, 66, 8, -93, -112, 5, -54, 36, 16, -87, 73, 105, -54, -69, 68, -58, 73, 65, 20, -10, -37, 127, -55, -90, 68, -80, 80, -86, -120, 95, 1, -45, -6, 51, -56, 110, 37, -59, -98, 15, -93, -33, -119, 8, 63, 79, 111, -49, -118, 57, 36, 58, 85, 37, 93, 18, -23, -120, -55, 7, 3, 84, 111, -127, 16, 80, -90, -55, -93, -121, 7, -128, -127, -84, -16, 117, 7, 59, 91, -103, -15, -10, 123, 24, -95, -31, -6, 18, -98, 120, 127, -13, 14, -117, 60, 62, 118, 125, -54, -16, 109, 0, 125, 20, -49, -82, 35, 66, 29, -126, -21, -63, -65, -87, 45, -81, 124, 77, 36, 57, -24, 99, 12, 37, -30, -56, 98, -40, 81, 42, 54, 34, 104, 14, -48, 42, -30, -7, -96, -120, -55, -114, -51, -41, -33, -20, -45, -92, 107, -58, 31, -82, -104, -24, -30, -25, -42, 118, -77, -97, -81, 88, 72, -68, 76, 87, -15, -40, 84, 12, -98, -113, 16, 2, -20, -115, 43, -6, -104, -101, 20, 127, 49, -21, -57, -116, -27, 35, 72, 57, 67, 2, -115, -78, -66, -38, -76, 108, -99, -89, -88, -105, -98, -120, 25, 40, -23, 15, 14, 119, 44, 8, -93, 0, 105, 20, -5, -102, -31, -75, -57, 23, 99, -82, -21, -15, -108, -41, 36, 57, 70, -81, -26, -98, 36, -57, 61, -16, 110, 17, 91, 0, -56, -55, 48, -26, 109, -110, 66, -71, 98, -41, -105, 86, 34, 53, -50, -61, 107, -8, -118, -22, -68, 46, 86, -31, -17, -53, 9, -68, -99, -20, -3, 22, 7, -122, 102, 68, -30, -128, 98, -17, -41, 14, -25, 102, 12, -56, 75, 52, -115, -100, 64, 105, -42, 113, 27, 123, 115, 72, 104, -32, -116, -6, -84, -106, -58, 126, 119, 98, 14, 83, 107, -82, 37, 123, -42, -51, 84, -28, 88, -85, 49, 68, -2, 126, 43, -58, 15, -122, -98, 28, -61, 56, 95, 46, -84, -103, 47, 60, -80, -111, 90, 127, -103, 63, 66, 34, -79, -71, 1, 4, 122, -68, -62, 48, 68, -56, 104, 79, -103, 96, 78, 25, -64, 56, -127, 90, 98, 82, -66, -117, 91, 82, 94, 24, 68, -60, -20, -4, -71, -57, 11, 46, 66, -86, 105, 23, 127, 52, -112, -42, -53, 101, -122, -54, -114, -22, 47, -38, -72, -7, -96, 116, -27, 47, -104, -84, 94, 19, -117, 16, -38, 68, 121, 34, 1, -75, 117, 93, -69, -42, -46, -6, -67, -69, 123, 125, 81, -103, 55, 95, 54, 112, -8, 105, 98, 113, -4, -84, -102, 17, 107, 91, 44, 52, 26, -120, -112, -90, -118, -66, 4, 88, -33, 13, -85, 46, 68, -126, -7, -53, -27, -2, -90, -68, -41, 22, 39, 86, -27, -56, 117, 102, 79, 84, 50, 52, 36, 78, -102, 24, -104, -38, -92, 2, 5, -54, -73, 127, -31, -118, -89, -38, 19, 111, 126, 124, 71, 112, 64, -73, 111, 23, 114, 122, -15, -102, 62, 41, -94, 63, 65, 37, 47, -90, -109, 6, -42, 36, 11, -30, -22, 72, 41, 100, 8, -124, 117, 97, 70, -43, -66, -125, -74, -50, -106, -116, -108, 41, 103, 28, 111, 12, -11, 84, -68, 75, -81, 70, -41, 106, 118, 93, -41, 10, -17, -124, 95, 63, -35, -9, -95, -113, 42, -61, 60, -87, 51, -87, -49, 45, -127, -74, 93, -94, -106, -45, -69, 8, 33, -115, 76, 66, -80, 111, 58, 116, 28, -53, -55, 54, 101, 80, -38, -26, 9, -44, -102, -68, 18, 105, 25, -117, -126, -17, -72, -59, -58, 114, 108, 31, 16, 126, -32, -81, 56, 105, -81, 78, 34, -63, 54, -88, -90, 121, 110, -95, -100, 51, -9, 37, 114, -91, 124, 103, 16, -111, 45, 48, 24, 3, 0, 56, 89, 73, 58, -55, 46, -95, -117, 100, -3, -6, 110, 70, -59, 62, -121, -38, -111, 112, 93, -117, 12, 4, 66, -56, -50, -99, 57, -112, 4, -58, -84, 116, -73, -51, -48, 14, -111, 18, 99, -4, -61, 112, 10, -40, 84, 87, 113, 75, -127, -52, 46, 71, 83, -66, -45, -25, 30, 120, -117, 109, -73, -77, -101, -47, -99, -82, 34, 18, 122, -52, -107, 4, -115, 60, 46, 18, -75, -103, -71, -98, -78, -46, -70, -62, 3, 72, 115, 94, -104, 118, 24, -14, 65, 127, 32, 29, 117, 84, 123, 14, 25, -37, -41, -12, 3, -24, -47, 30, 33, 98, 99, -50, -102, 64, 3, -48, -46, 19, -89, 83, 78, 0, -85, 121, 41, 6, -120, 111, 26, -26, -17, -104, -80, -124, -3, 53, -19, 82, -59, -8, -113, -23, 53, 5, 103, 2, -15, -49, 21, -111, 121, 12, -10, 52, -69, -75, -60, 83, 21, -103, -109, 3, 100, 126, 43, -16, 29, 120, -94, -99, -89, 12, 75, -114, 115, 85, 1, -68, -74, -51, 69, 71, -71, 46, -60, -88, 74, 60, 117, 112, -122, -97, -75, -88, 57, 81, -72, -66, -99, 84, 74, -122, 21, -93, -41, -36, -46, 39, -109, -49, 26, 15, 35, 34, 6, -3, 88, -105, -32, 102, -31, -88, 64, 100, -117, 4, -52, -24, 68, 92, 47, -94, -17, -89, 81, 59, -1, -64, 57, -50, -37, -54, 112, 34, 57, 3, -55, -10, -99, 83, 26, -105, 117, 29, 81, -87, 95, 63, -35, -25, -119, -76, -98, -53, 70, 111, 7, -28, 81, 116, -83, -10, -19, -68, -54, 115, -54, -88, -106, 64, -36, 120, -5, 81, -101, -58, 54, 122, 24, -63, -45, 42, -72, 10, -4, -7, -29, 31, 45, 83, -90, 28, 18, 114, 101, -9, 90, -48, 103, 76, -106, 58, -102, -121, 118, 96, -63, -45, 54, -68, -48, -28, 99, -70, 106, -110, 105, 109, 5, -29, -110, 91, 30, -86, 64, -57, -68, 64, 99, 7, -31, -4, 73, 63, -50, -2, 7, 2, -64, -78, -8, -39, -64, 102, -126, -98, -68, -75, 30, -58, 86, 15, -70, -53, -50, -4, 35, -57, -117, 28, -99, -36, -106, 116, 98, -25, -15, 29, 4, 82, -26, -58, -19, 28, 109, 43, 17, -127, -113, 59, 90, -91, -103, -43, 61, 25, 30, -78, 2, -72, -34, -79, 46, -50, 75, 88, -80, -65, 78, 11, 4, 115, -26, -97, 100, -128, 83, -117, 11, -82, -63, 53, -116, -28, 109, 72, -9, -65, 73, 127, 89, 73, 69, 27, 115, 81, 83, 38, -29, -21, 81, -68, -110, -107, 35, 27, -50, 28, -16, -3, 9, 68, -29, 16, -63, -58, -39, -55, -124, 101, 32, 75, 49, -117, 46, -45, -124, 107, 71, 24, 3, -121, -106, -47, 90, -105, -104, -24, 106, -25, 33, 0, 92, 62, -108, -115, 124, -82, -119, -76, 91, 55, 4, 63, -91, 80, -106, 91, 124, 91, 100, 55, 107, -47, 24, -95, 57, -53, -68, -5, 109, 72, 76, -103, -118, -65, -104, 93, 127, -63, 1, -69, -78, 36, -115, -5, -68, 51, -50, 26, 86, -85, 97, -63, 89, 18, 106, 21, 90, -93, -78, -61, 76, 47 );
    signal scenario_output : scenario_type :=( -128, 127, -128, -16, 127, 127, 127, -39, -128, -128, -128, -128, -128, -128, 127, 127, 33, -128, -128, 66, -128, -128, 127, 127, 127, -128, 127, 127, -128, -48, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 65, 127, 127, 127, 127, 127, 127, 127, 127, 127, 23, 127, 127, 127, 127, 127, 127, 127, 127, -11, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 24, 127, 127, 127, -114, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -17, 127, 127, -128, -128, 127, 127, -128, 58, 127, 127, -128, 127, -128, -128, -128, 127, -47, -128, -2, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 117, -128, -128, -128, -128, 127, 127, -128, -128, 127, -76, 127, -128, 127, 127, 119, -128, 127, -128, -128, -128, -128, -118, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -127, 127, 127, 127, 127, 127, 127, 127, 0, 127, 127, 127, 127, 127, 127, 127, -128, -128, 28, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 123, 127, 127, 127, 127, 127, -128, -128, -128, -63, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 102, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -3, 98, 49, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -50, 127, 127, -128, -128, -95, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -16, -128, -128, -128, 111, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 63, 127, -17, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 29, 127, -128, -128, 113, -118, -128, 38, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 7, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 53, 127, 60, 127, -12, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, 88, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 81, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -8, -128, -128, 127, 127, 127, 127, 127, -17, -11, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 10, -128, 127, -128, -43, 127, 108, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -88, 127, -128, -128, -123, -128, -128, -128, 127, -128, -128, -128, -12, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 37, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -64, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 74, 127, 127, -128, 127, 127, 127, 127, 127, 42, 127, -128, -128, -128, 7, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -3, -128, -12, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 123, 127, 127, 88, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -119, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 102, 127, -128, 127, -128, -128, -128, 26, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 80, 127, -49, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 8, -128, -128, -128, 127, 127, 127, 127, -128, 52, -47, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -74, 127, -128, -128, 87, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 74, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -96, 127, 127, 127, 127, 127, 127, -128, -128, -128, 2, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -43, -128, -128, 127, -128, -128, -128, -128, -128, -63, 127, 127, 127, 127, 127, 127, 127, 26, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 15, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -71, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 76, -128, 54, -128, -128, 127, 127, -128, 50, 127, -128, -128, 127, 127, 127, 127, 127, -128, 44, -128, 127, 127, -24, -128, 127, -128, -128, -128, -128, 127, 127, -52, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 45, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 101, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -76, 0, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 12, 127, 127, 127, 127, -128, 127, 127, 36, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 103, 127, 127, 127, 21, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 15, -128, -47, 127, 127, 127, 127, 127, 127, 127, 65, 127, 127, 127, 127, 127, 127, 127, 127, -8, -128, -128, 92, -128, -128, -128, -102, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -13, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 17, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 55, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 57, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -7, -128, -128, -70, 127, -128, -128, 127, 127, -76, -128, 127, 127, -23, 127, 127, 127, -128, -128, -74, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 50, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 17, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -26, -128, 127, 78, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -79, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 95, 127, -11, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -98, -128, -128, 127, 127, 127, 127, 127, 127, -66, 127, 127, 127, 69, -128, -127, -128, -71, 127, 127, 127, 127, 127, -128, -29, -128, -128, -128, -128, -128, -128, 112, 44, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -109, -128, -128, -63, -128, -128, -7, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -91, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 18, -34, 48, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 12, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 59, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 2, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 68, -128, 127, -128, 127, 79, 127, -128, -128, -111, -128, 127, 127, 127, 50, 127, 127, -102, 127, 127, 127, 127, 127, 127, -128, 73, 127, 127, 127, 127, 127, 127, 127, -128, 127, 101, 127, 127, 127, 127, 127, 109, -64, -128, 127, 127, -69, -128, 127, 127, 127, 127, 127, 0, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -106, -128, -128, 127, 127, 127, 127, 127, 127, 127, 113, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -73, 127, -128, -128, -128, -128, -128, -128, 127, -119, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 26, 26, -128, -128, 127, 127, 127, -79, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 60, -55, -128, -128, 127, 127, 127, -128, 78, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -73, 109, 127, 127, 127, -128, 116, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -11, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 8, -128, -128, 127, 127, 53, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 70, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -111, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -59, -128, -128, 127, -128, -128, -128, -128, 127, 127, 65, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 44, 127, 127, 127, 121, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -5, -128, -128, -128, -128, -128, 28, 127, 127, -86, 65, -128, -128, 127, 127, 127, 127, -50, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 71, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 116, 127, -128, 127, -112, -128, -128, 127, -32, 127, 127, 127, 127, 127, -128, -128, -128, -17, -128, -128, -128, 127, -128, 127, 7, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -88, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -96, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -96, 127, -128, -128, -128, -128, -47, -128, 111, -128, 127, 81, -128, -128, -128, -128, -128, 49, -128, -74, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 54, 127, -128, -128, 127, 127, -128, 102, -128, -75, -128, 127, 127, 127, 127, -128, -128, -128, 39, -128, -128, 127, -128, -128, 127, -43, -128, 127, 127, -92, 127, -2, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, -101, -128, -128, -128, -128, 127, -65, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 38, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -55, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 17, -128, -128, -128, -128, -128, -128, 71, -128, -128, -128, -128, -128, -128, 127, 74, -128, 127, 127, -128, 127, 127, 127, -128, 127, -12, 10, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -58, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -36, 127, 127, 127, -23, 127, 127, 127, 127, 127, 127, 127, 127, -122, -128, -128, -128, -128, -128, -128, 52, 127, -114, -10, 127, -128, 127, -128, 127, -128, 127, -128, 87, -128, -128, -128, -128, -128, -128, 68, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 57, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 24, -128, -128, 127, -24, -128, -128, -128, -128, 127, -128, -128, -63, -128, 127, 127, 127, 127, 127, 127, 127, -11, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 95, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 119, 127, -128, -128, 127, 127, -128, 127, 127, 127, -101, 127, -128, 127, 70, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -107, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 121, 127, 127, 127, 127, 119, 127, -128, -128, 127, 127, -22, -128, -128, -128, 127, -93, 63, -128, -128, -128, -128, -2, -128, -128, -114, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -39, -128, -50, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -78, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -54, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -122, -128, -128, -128, -128, -128, 127, -128, 37, 127, 127, 10, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -7, -39, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 6, 71, -128, -128, -128, -128, -118, -128, 127, 127, 127, -128, 127, 127, 127, 127, -78, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 42, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 3, -128, 112, 127, 127, 127, 127, 26, -128, -128, 23, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 118, 127, 127, 127, 127, 127, 127, 127, -128, -128, 21, -128, -128, -128, 127, 127, 127, 127, 127, 127, 108, 127, -128, -57, -36, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 16, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 90, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -60, -128, -128, 127, -128, -128, -128, -128, -128, 71, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 116, 127, 127, -128, -128, 127, 0, -98, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 7, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -75, 127, 26, -128, -128, -128, -128, -128, -128, 31, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -59, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 45, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -76, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 49, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 71, 127, -128, -128, -128, -128, -128, -128, -128, 127, 36, 127, 127, 127, 0, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 53, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 111, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 17, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 65, -128, -42, -128, -128, -128, -128, 127, 127, 47, -12, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -45, -128, -21, -128, 127, -31, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -32, -128, -128, -128, -128, -128, -128, 127, 127, 127, 109, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -68, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 79, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -69, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 38, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 11, 127, 127, -128, -128, -74, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 43, 127, 127, 54, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 34, -11, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 36, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 117, 75, -128, -128, -128, -5, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 59, -128, -128, -128, -128, -128, -128, -128, -128, -91, -128, -128, -128, -128, -128, -128, 127, 81, 127, 127, 127, 127, 37, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 24, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, -10, -128, -128, -128, -128, -128, -128, -128, 127, 95, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -117, -128, -128, -128, -128, -128, -100, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 122, 127, 127, -128, 127, -91, 86, 49, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -42, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -22, 127, 127, -128, -128, -128, -128, -128, -128, -128, -33, -2, -128, 34, -128, -128, -128, -128, -128, 58, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 70, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 117, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -17, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -57, -128, -128, -128, -128, 127, 127, 127, -128, 64, -128, -128, 93, 127, -112, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 97, 127, 127, -128, -128, 127, -128, -128, -55, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -75, 127, -86, -128, -128, 71, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -96, -58, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -34, -128, -118, 127, 127, 127, 127, 127, 127, 127, -128, -121, 127, 127, 127, 127, 127, 127, -128, -22, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 12, -47, -128, 127, 127, -128, -128, 127, -70, 127, 127, 127, 127, -128, 127, 127, -128, -100, 127, -128, -128, -128, -128, -128, -128, 127, -128, -37, -128, -128, -128, -128, -128, -128, -128, -101, -128, -128, -128, 127, -128, -128, -128, -128, -93, 127, 127, 127, 127, 127, -128, -8, 127, 127, -128, 127, 127, 127, 127, 118, 127, 127, 127, 127, 127, 127, 127, 127, 127, -68, 93, 127, 127, 127, 127, 127, 127, 117, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 64, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -16, 127, 127, -128, 86, 127, -128, -55, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -95, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 65, 95, 127, -81, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 36, 127, -128, 127, 127, -32, -15, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 118, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 42, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 88, -128, 127, 127, -128, -128, 127, -48, -128, -73, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -101, -75, -128, -128, 127, 127, 47, -123, 127, 127, -68, 127, 127, -118, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 73, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -65, 127, 127, 127, 127, 127, 127, 127, 127, 127, 112, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -69, -128, -128, -128, 0, -122, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 74, -128, -128, 127, 127, -128, 63, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -76, -128, 127, -128, 127, -38, 127, -128, 127, -128, -128, -128, 53, -128, 29, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 22, -65, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -127, -128, 11, -128, 70, -128, -69, -128, -128, -128, -128, -128, -128, 80, 127, -128, -128, -128, -128, -128, -128, -128, -128, -112, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -54, -128, -128, -31, 127, 127, -112, 127, 36, -128, -116, 127, 127, 127, -128, -11, -128, -128, -128, -128, 127, 127, 127, 124, -128, -128, 118, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 111, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -58, -128, -128, -44, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -22, -128, -128, -128, -128, -128, 127, 13, -128, -128, 127, -128, -128, -128, 127, -3, -128, -128, -128, -128, -128, 127, -128, -128, -55, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -22, -128, 127, 65, -128, -128, -7, -128, -79, -128, 127, -128, 127, -45, -128, -128, 117, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 21, 127, -128, 127, -128, 127, 127, 127, 122, -128, 127, -128, -128, -79, -128, -128, 127, -108, -47, -128, 127, 127, 127, 127, 127, -101, -128, -128, 127, 127, 127, 127, 127, 81, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 50, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 114, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -76, -8, -128, -128, -128, -128, -128, -128, -128, -128, 27, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -28, -128, 127, 127, -10, 127, 127, -128, -128, 127, -86, 127, 127, 127, 127, 127, -10, 127, 127, 127, 127, 127, 97, 127, -128, -128, 127, 127, 53, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -49, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -74, 127, 127, 127, 127, 127, 127, 127, 127, 7, -128, -128, -128, -128, -128, 8, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -27, 8, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 31, 127, 127, -128, -128, -38, 127, -58, 127, 127, 127, 39, 127, 127, 127, 127, 127, -128, -128, -128, 70, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -32, 117, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 21, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -33, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 34, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 53, 127, 127, 127, 127, 127, 127, 127, 111, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -24, -128, 127, -128, 116, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -50, -128, -128, -128, 127, -128, 39, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 101, 127, 127, 127, 127, -128, 127, -128, -128, -128, -71, -128, -128, 16, 127, 127, -128, 127, -128, -128, -128, 113, -128, 8, -128, 127, 127, -80, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -71, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -111, 127, 5, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -47, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 50, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -66, 127, 127, 127, 127, 127, 127, 127, 127, 127, 102, 86, 74, -128, -128, -128, -128, -128, -128, -128, -128, -128, 0, 127, 127, 127, 127, 127, 127, -33, 127, -128, -128, -59, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -45, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -26, 127, 127, 127, 119, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -107, 127, 127, 127, 127, 127, 127, 2, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -119, -106, -128, -128, -128, -128, -128, 127, 127, -128, -21, 127, -63, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 18, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 88, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -58, -128, -112, 127, 127, -24, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -86, -128, -128, 127, -128, -128, 127, 118, 18, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -23, 127, -103, -21, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -92, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -111, -128, -128, -128, -128, -128, 127, -100, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 63, 127, 48, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 112, -128, -128, -95, -37, 127, 127, 127, 127, 127, -128, 127, 127, 18, -128, 127, 127, 127, 127, 127, 127, 127, 69, 127, 127, -74, -128, 127, -106, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 26, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -76, 127, -78, -128, -128, -128, -128, -128, -128, 28, 127, 127, 127, 127, 127, 127, 96, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -79, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 0, -128, -17, 127, -95, -128, -128, 127, -1, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 100, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -24, -128, -128, -128, -128, -128, -128, -116, -128, -128, -128, -33, 127, -128, -128, -128, 127, 127, 127, 111, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 75, 127, 48, -128, -128, -79, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 5, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -98, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -28, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 95, -128, 127, 127, 127, 127, 127, -43, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -16, 106, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 114, -128, -128, 127, 127, 127, 127, 127, 127, -128, -93, -128, -128, 127, -2, -128, 113, 127, 74, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 24, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 100, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -100, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -31, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -15, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 91, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -101, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 69, 127, 112, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -52, 127, -128, -128, -128, -128, -128, -64, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -107, -128, -128, -128, -128, -128, 127, 127, 127, -128, 88, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -97, 127, -128, 127, -36, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 23, 127, -128, 127, 127, 127, 86, 127, 127, 127, 127, 127, -23, -128, -119, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 78, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, 98, 127, 127, 127, -128, 127, 127, -128, -91, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -106, -70, -5, 127, 127, 124, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -50, -128, 81, -128, 127, 127, 127, 127, 127, 127, 127, -11, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 112, -128, -26, 73, 127, -128, 127, -128, 24, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -86, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 10, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -123, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -29, 127, 127, 48, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 70, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 5, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -27, 32, 49, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -37, -128, -128, -128, -39, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -11, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 74, 127, -73, 127, -128, 127, 127, -128, -87, 127, 127, -128, 127, -128, -128, 2, -128, -128, 127, 23, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -86, 127, 127, 127, -128, -128, -128, -128, 44, 127, 127, -6, -128, 127, 127, -128, -128, 127, -128, -128, 127, -12, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -60, -128, 85, -128, 127, -85, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 106, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 8, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 90, -128, -128, -128, -128, -128, -128, -128, -128, 117, 127, 127, 127, 127, 127, 127, 127, 127, 7, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -36, 127, 127, 127, 127, 127, 127, 127, 59, 127, -128, 127, 127, 127, 127, 127, 127, 127, 93, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -3, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 108, -128, -128, -21, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 124, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -108, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -87, 127, 127, -128, -128, -128, -128, 127, 127, -118, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 1, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -21, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -76, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 88, 70, -128, -128, -128, 127, 127, -102, 0, 127, 95, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -68, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 0, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -101, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -96, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -54, 127, -75, 127, 106, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 63, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -80, 127, 127, 127, 90, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 122, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -71, 127, -128, -128, -128, 127, -128, -128, 109, 127, -128, 127, 127, 127, -128, 127, 127, -128, 63, -128, -128, -128, 127, -128, -128, -128, -128, 26, 127, 127, 127, 127, 127, -45, -128, -128, -128, -128, -85, 127, 127, 127, 127, 127, -128, 127, 127, 23, 127, 127, 127, 127, 127, 127, 127, -128, 49, 127, 127, 127, 127, 127, 7, -121, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 28, -128, -128, -71, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -47, 127, -128, 127, 127, -128, 127, 127, 15, 66, 127, 127, 49, -16, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 116, 127, 127, -128, -128, -128, -128, 127, 91, 127, 127, 127, -128, 127, 127, 127, 107, 127, 127, 127, 127, 127, -128, 118, 127, -128, -128, -128, -128, -128, -128, -73, -128, -128, -128, -128, -128, -128, -128, 127, 2, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -78, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -86, 73, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 101, 127, 127, 127, 127, -128, 15, -27, 127, 103, -114, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -38, -128, 112, -81, -128, -128, -128, -128, 127, 127, 114, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -117, 117, 127, 93, 127, -128, -92, -128, -112, -128, -128, -128, 127, -128, -128, -128, 127, -119, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 106, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -32, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -43, -128, -128, -128, -128, -103, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -28, -102, 127, -128, -128, -128, -128, 34, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 108, -128, -128, 127, -5, -128, 127, 127, -128, -128, -128, 127, -128, 127, 74, -11, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -69, 127, -128, -128, 127, -128, 127, 127, -66, 127, -128, -73, -128, -128, -128, -91, 127, 127, 127, 127, 127, 127, 127, -128, -15, 127, 127, -39, 127, 127, 127, 127, 127, 127, -128, 29, -128, -38, 127, 127, 127, 127, 127, -128, 127, 43, 127, 127, 127, -128, -128, 127, -128, -128, -79, 127, 127, 127, 127, 127, 127, 127, 32, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -36, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -85, 127, 127, -98, 29, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -17, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 122, -119, -128, -128, 127, 127, -60, -128, 52, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -8, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -107, 127, 127, -58, 127, 127, 127, 10, 127, 127, -119, 127, 127, 127, 127, 127, 127, 127, 127, 127, -107, 127, 45, 127, 127, 127, 127, -44, -128, 127, 127, 127, 127, -17, 127, 80, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -22, 52, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 63, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -86, -128, -128, -128, -128, -78, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 93, 127, 127, -128, 127, 127, 127, -116, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 80, 127, 127, -28, 127, 127, -128, -128, 127, -128, -128, 127, 127, 95, 127, 127, -128, 34, -63, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -73, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -45, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 3, -128, -128, -128, 124, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -28, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 58, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 58, -128, -128, -128, -128, -128, 81, -128, -128, 127, -42, -128, 18, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -5, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 70, -128, -128, -128, -128, -128, -128, -128, 0, -128, -128, -128, -28, -128, -128, -128, -128, -128, -43, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 81, -128, -128, -128, 127, -128, 127, 127, 127, 87, 127, 127, 127, 60, -128, -22, -128, -128, -128, -58, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -109, -128, -128, 127, 127, 127, 127, 127, 127, 127, -53, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -3, 87, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -32, -128, 58, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -21, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 64, 64, 80, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 87, -128, 127, 127, 127, -101, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -44, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -43, -128, -128, -128, -128, -128, -128, -128, -24, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -100, 111, -5, 81, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -16, 127, 127, 127, 127, 127, 127, 127, -112, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 57, -128, -128, -128, 127, 55, -128, -128, 127, 127, -128, 127, 127, 45, -128, -128, -128, -128, -128, -128, 17, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -47, -47, 127, 127, -63, -128, -128, -128, 6, -128, 127, -128, -128, -128, -128, -128, -76, 36, -128, -128, -128, -128, -128, -128, -128, -128, -128, -76, 127, 127, -15, -52, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 21, -124, -128, 117, 127, 127, -128, 127, -128, -128, -128, 127, 127, 48, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 80, -32, 127, 127, 127, 90, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -53, -128, 127, 127, -128, 127, 36, -128, -128, -128, -128, -128, 127, 69, 127, 127, 34, -128, 127, 127, 127, -128, -128, 17, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 69, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 96, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -92, 127, -128, -128, 36, -128, -128, -128, -128, 127, -128, 16, 127, 127, 127, 127, 117, -128, 127, 127, 127, 29, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -39, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -98, 127, 127, -128, 26, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -90, -128, 127, -85, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 50, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 10, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 59, 127, -128, -128, -128, -128, -128, 127, -53, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -97, -128, -128, 127, 127, 127, 127, 127, 127, -78, 127, 127, -128, 127, -128, 69, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 7, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 44, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -127, -128, -128, -128, 127, 10, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 96, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -58, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -15, -128, -128, -128, 92, -128, -128, 127, 127, 100, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, 38, -128, 11, 127, -128, 2, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 5, -128, -128, 127, -128, -128, -128, -128, -128, -128, -71, 127, 127, 127, 127, 127, -106, 127, -128, -128, -86, 127, 127, 127, 127, 127, 127, 127, 127, -21, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 11, -128, 31, 127, 127, 127, 127, 127, 127, 127, -128, 114, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -63, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 7, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 24, -128, -128, 127, -1, -128, 127, -128, -128, -128, -128, -128, -128, 58, 127, 127, -128, 127, 127, -128, -128, 48, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -38, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -2, -128, 57, -128, -128, -128, 127, -11, -128, 95, 127, 6, 127, 127, 127, -128, 127, 127, 127, -45, 127, 127, 127, -128, -128, 127, 127, -128, 16, 127, 127, 127, 127, 127, 11, -128, 127, 127, -92, 127, 127, 127, -66, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -124, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -28, 22, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -70, -111, -128, -128, -128, -128, -48, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -59, -128, -128, -128, -128, -128, -128, -128, -128, 32, -128, 127, 88, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -73, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 85, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -44, 127, 127, -128, -128, -128, -128, -73, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -42, 127, 127, 127, 127, 127, 127, 127, 127, 127, -60, -128, 1, -128, 127, 127, 127, 127, 127, 127, 127, -42, -128, 127, 127, 127, 127, 127, 127, -49, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -69, 127, -128, 127, 127, 79, -106, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 2, -70, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -79, -128, -128, -128, -128, -128, -128, 127, 117, -128, -128, 127, -128, -128, -58, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 102, -128, -128, -128, 127, 127, 127, -116, 16, 127, 127, -128, -128, -128, 32, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -106, -128, 127, 10, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 42, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, -31, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 11, 21, 127, 127, 127, 127, 127, 26, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -119, -128, -54, -97, -128, -128, 127, 127, -128, 127, -128, -128, -75, 127, 127, 127, 127, 127, 127, 121, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -60, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 55, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 87, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -101, 127, 127, -128, -128, 108, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 109, -128, -128, 127, 116, -128, 127, -128, 88, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 103, -128, -128, -128, -37, -128, 127, 127, -128, -128, -44, 58, -128, -128, -128, -128, -128, -92, -128, 127, 127, 127, 127, 127, -45, -85, 0, -128, -128, -128, -128, -128, -128, -127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 119, -128, 127, -128, -128, -128, 127, 127, -128, 127, -39, -128, -128, -128, -128, -128, -128, -128, -11, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -116, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 26, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -26, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -12, -128, -128, 23, 127, -60, 127, -128, -128, 127, -128, 127, -10, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 68, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -27, 90, -128, -128, -128, -63, 127, 127, 127, -128, 127, 117, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -8, -128, -128, 33, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 79, -128, -128, -44, 127, 127, 127, 127, 127, -119, 127, -128, -128, 127, 127, -128, -8, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 37, -128, 127, -128, -128, 54, 127, -128, 127, 127, -128, -128, 69, -128, -128, -128, -128, -128, -128, -128, -124, -128, 127, 79, -128, 127, -128, -128, -128, -128, -128, -128, -128, 22, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 90, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 103, -128, -128, -128, 127, 127, 127, 127, 127, -16, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -5, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 54, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -38, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -31, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 124, 2, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -86, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -92, 93, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 27, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -91, -128, -128, 127, -128, -128, 127, -60, 127, 127, 127, -87, 127, 127, 127, 127, 127, 127, 127, 127, 127, -13, 78, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 16, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -116, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 13, -58, -128, 127, -128, -47, 127, 127, 127, 127, 127, -128, -70, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 112, 59, -48, -128, -128, -128, -128, -128, -22, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -10, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 17, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -109, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 52, 127, 127, 127, 127, 10, -128, -128, -128, -128, -39, 127, -128, 127, 127, 57, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 60, -128, 127, 127, 127, -69, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, 93, 127, 127, 127, 127, 127, -128, 127, 127, -86, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 52, -128, -128, 127, 127, 127, -11, -124, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 114, -96, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -24, 127, -128, -27, -128, -128, -114, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -68, -128, -128, 127, -128, -50, -49, 127, 127, 127, 127, 127, 127, 127, 127, 36, -128, -128, -128, -128, -128, -128, -128, 127, 127, -98, 127, 127, 127, 127, 127, 127, 127, 127, 127, -90, -128, -128, -128, -128, -128, -116, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 66, -21, 127, -128, -128, -128, -128, 127, -128, 50, 127, 127, 127, 127, 127, 127, 127, 127, 127, -122, -128, 90, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -8, 127, 127, -34, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 119, -128, -128, -128, -128, -128, -26, -128, -128, -128, -128, -128, 33, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 7, -128, -128, 100, -128, -128, -128, -128, 16, 60, -128, -128, 127, 127, -128, -128, -128, -128, -128, -112, -128, -68, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -122, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -2, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -31, 127, 127, 127, -128, 121, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, 43, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -103, 127, 127, -108, -128, 127, -128, -128, 127, -27, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -38, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -119, -128, -128, 127, 127, -128, 127, 118, -6, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 7, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 98, -128, -128, 116, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -5, 127, 127, 127, 127, 127, 127, 127, 127, 127, -23, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 74, 127, 127, 127, 127, 127, 127, 127, 3, -128, 127, -128, -128, -128, -42, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 70, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -112, 127, 127, 127, 127, 127, -128, 15, 127, 127, -128, 127, 127, -70, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -34, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -109, 93, -128, -128, -128, -128, -128, -113, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 124, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -43, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -108, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -73, -128, -128, 127, -128, -128, -128, 127, -114, 3, 127, 127, -128, 127, -114, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -78, 127, 127, -128, 127, 127, 127, -128, -123, -128, -128, -128, -128, 127, -123, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 122, 127, 127, 127, 127, 127, 121, 127, 127, 127, -1, 127, -66, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -18, 12, -128, 127, 127, -97, -128, -70, -128, -128, -128, -128, -128, -128, 127, 127, -50, -44, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 98, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -90, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 54, 127, -7, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -76, -128, 127, -85, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -107, 75, 127, 127, -128, -128, -128, -128, -69, 28, -128, -128, -128, -128, -128, -128, 95, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 24, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -27, -128, -128, -128, -128, -128, -128, 127, -128, -65, 127, 127, 23, 127, 127, 127, 127, 127, 122, -128, -128, -128, -128, -128, -128, -128, -128, -50, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 76, -128, -128, -119, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -54, -128, -128, -128, 59, -55, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -79, -128, -128, 127, -128, 127, -128, 127, 127, -6, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -71, -128, 127, -96, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 75, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -47, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 36, -128, -128, -128, 127, -128, -118, 127, 127, -128, -128, 101, -128, -128, -128, -128, -128, -49, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 13, -128, -128, -128, 1, 127, 127, 127, 127, 127, -107, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -29, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -101, -128, -121, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -13, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 123, 127, -128, -128, 127, 127, 71, 127, 127, 127, 127, 127, 119, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -8, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -98, 127, 127, 127, 127, 24, -128, -128, 101, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 118, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -58, 127, -114, 127, -78, 127, 127, 127, 127, 127, 127, 127, -60, 78, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 42, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 18, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 124, -128, -128, 127, -3, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -78, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -101, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 32, 127, 127, -128, -128, 127, 114, 101, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 23, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 27, 127, 127, 127, -128, 127, 127, 113, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 34, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -113, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 45, -128, -128, 127, -128, 127, -128, 127, -128, 34, -128, 127, 127, 127, 127, 44, -128, -128, -128, -78, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -79, -128, 127, 127, 127, 127, 127, -114, 32, 63, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 97, -128, -128, -128, -128, -128, 127, -128, -95, -123, 127, -128, 127, 127, 127, -26, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 95, 127, -128, 17, 127, 127, -128, -128, 66, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 109, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 43, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 29, -78, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 69, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -63, -128, 127, 127, -128, 112, -128, -128, -37, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 18, 127, -128, -55, -98, -16, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -95, 127, 75, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 22, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 112, 74, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 111, 65, 2, -6, 127, 127, 127, -128, 48, -128, 127, 127, 127, -24, 127, -128, 127, 127, -128, 127, 127, -128, -79, 127, 118, 127, 127, 127, 127, 127, 127, 103, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 71, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 68, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 12, -128, -128, -128, -128, -128, -128, -106, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 111, -128, -128, -128, 127, -108, 127, -128, 127, -128, -128, 96, 127, -128, 0, -128, -128, -128, 127, -128, 127, 127, 13, 109, 127, 127, -128, 48, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -65, 127, 127, -114, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -85, 127, 127, -75, -128, -64, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 33, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -55, 7, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 18, 21, -128, -128, -128, 127, -128, 127, 127, -48, 29, 127, 127, -128, 26, 127, -43, -128, 127, 127, 127, -128, 127, -128, -128, -128, -117, -128, -128, -128, -128, -128, -10, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -75, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 124, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 50, -23, -128, 32, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 71, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 58, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 100, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 92, -128, 127, 127, 127, 127, 127, 127, 127, 71, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -86, -128, -128, 122, 127, -128, 127, 127, 127, 108, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -112, 127, -128, -128, 127, 127, 22, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -107, -128, -128, -128, -128, -128, -128, -128, 10, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 64, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 75, 117, -128, -80, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 124, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -79, -128, -128, 127, -63, 127, 127, 127, 127, 127, 127, 127, 39, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -33, 31, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 33, 44, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -86, 127, 116, -128, -128, -128, -128, -128, -128, -64, 23, -128, 127, 1, 71, -128, -128, -128, -128, 57, 127, 127, 127, 127, -128, -85, -128, -128, -128, 37, -128, 127, 127, -43, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 97, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 12, -128, -128, 127, -128, 127, -37, -80, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 79, 127, -128, -128, -128, -128, -128, -128, -90, -71, 127, -64, 22, 123, 127, -106, -128, -128, 127, -128, -128, -128, -128, -128, -128, -65, 127, -128, -128, -128, 48, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -16, -100, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 48, -128, -128, -75, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, -65, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 21, 127, 114, 127, 42, -128, -128, 86, 127, -128, -128, -128, 118, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -109, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -42, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 70, -128, -128, -128, -128, -128, 127, -128, -121, 33, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 98, -128, -128, -128, -128, -128, -128, -52, 127, -128, 127, 127, -128, -128, -128, -128, -128, 36, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 86, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -118, 39, -128, 127, 127, 127, 127, 127, 127, -128, -58, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 31, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -114, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 65, -92, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -80, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 23, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -55, 127, 127, -128, -128, -50, 127, -128, -55, 127, 127, -15, -128, -128, -128, -128, -128, 26, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 21, -128, -128, -128, -128, -128, -128, -128, -128, -3, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -90, 127, 127, -128, 127, 127, 127, -128, -39, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -71, -128, -128, 127, 127, 127, 127, 127, 127, 127, -31, 127, 127, 127, -128, 127, -128, -60, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -122, 8, -18, 100, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -107, 127, 119, 127, 127, 127, 127, 127, 127, -128, -128, 45, -128, -128, -128, -128, -86, -128, -128, 127, 127, 74, 127, 127, 127, 119, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -58, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -91, -128, 127, 127, 127, 127, 127, -128, 53, 127, -128, -128, 127, -33, 127, 127, 127, 127, 127, -27, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -73, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -43, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 21, 127, -128, 127, -128, -128, -128, -128, -128, 127, -48, 127, 127, 127, 127, 127, -128, -128, 127, 127, 10, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 24, -65, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -24, 114, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 108, -128, -128, 127, -114, -128, -128, 127, -128, -114, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -79, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -74, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -26, -103, -75, 127, 127, -80, -128, 127, -119, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 73, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -38, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -26, 127, 127, -18, -15, 127, -128, 127, -15, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -103, -109, -68, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -63, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 119, 127, 127, 127, -128, 127, 127, -1, -128, 127, 1, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -23, 127, -13, -128, 96, -128, -44, -128, -128, -128, -128, -128, -128, 127, -128, -128, 79, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -86, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 69, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -79, -128, -128, 127, 127, 127, -44, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -27, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 8, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 32, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -123, -128, 127, 127, -128, 127, 127, 3, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -124, -128, 127, 127, 91, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -24, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -117, 127, -128, -128, 127, 127, -32, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 81, 127, -79, -128, -128, -128, -128, -128, -128, -128, -128, -118, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 42, -128, -128, -128, 127, 127, 127, -16, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -49, -128, -128, -128, -102, -44, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 58, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -63, 92, 127, -79, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 0, 127, 127, 127, 76, -128, -36, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 17, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -13, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -73, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 15, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 45, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -50, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -31, -128, -128, -128, -128, -128, 15, -128, 127, -128, -116, 37, 127, -128, 127, 122, 127, 127, -128, 127, 127, -128, -121, 127, -128, 127, 127, 127, 2, 127, 127, 127, -128, 127, -128, -128, -101, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 6, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 29, 127, 127, 127, 0, -128, -128, -128, -128, -128, 127, 45, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 47, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 8, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 23, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -18, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -37, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 90, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 45, 127, 127, 127, -128, 127, -90, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 43, 127, 127, -128, -128, -128, -128, -33, 127, 127, 127, 127, -128, 127, 127, 127, 85, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -32, 127, -128, -128, -128, 109, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 123, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -48, -44, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -22, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 54, -128, -128, -128, 127, -128, -128, -128, -93, -128, -128, 127, 127, 127, 127, 127, 5, 127, 127, 127, 127, 127, -55, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -63, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 108, 127, 127, 127, 127, 127, 127, 127, 127, -16, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -31, -128, -128, -128, -128, -128, -128, -128, 36, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -116, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 90, -27, 127, -128, 127, 127, -128, -128, -128, -128, -128, -31, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 50, 127, -128, 127, -70, -102, 127, -128, -128, -128, 127, -128, 127, 127, -22, -42, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -101, 127, 127, -128, 60, 127, 127, 127, 127, 127, -128, -128, -112, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 37, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -88, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 31, 127, 127, 18, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -93, -128, -128, -128, -128, -128, -128, -128, -128, -122, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 36, 127, -128, 127, 127, 127, -102, 127, -128, 88, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -70, 127, -128, -128, 127, -86, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 106, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -57, -87, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 78, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 122, 127, -128, -128, -128, -128, 127, -128, -128, 33, -128, -128, -128, -128, -79, 127, -128, -128, 127, 127, 127, 127, 127, -128, 6, 54, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 17, -97, 127, 127, 127, -17, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -8, -128, -128, -128, -128, 127, -128, 127, -128, 64, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 58, 127, -128, -128, 127, 127, 127, 69, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 8, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -112, 127, 127, 127, 127, 127, -128, -128, -128, -128, -90, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -43, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -5, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 80, -128, -128, -128, 127, -128, -3, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -55, -128, -128, 127, 127, 49, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -3, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -2, 127, 127, 127, -121, 127, 127, -119, 127, 127, 127, -95, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 50, 16, 39, 127, -128, -128, -128, -128, -128, -128, 127, -37, -3, 124, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -8, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 32, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -92, -128, -128, -33, 80, 127, 127, -128, 127, 127, -128, -32, 127, -128, -128, -128, -128, -128, 127, -60, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -2, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 8, -128, -128, 127, 127, -128, 127, 127, 127, -59, 127, 127, 127, -128, 44, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 26, -31, 127, 27, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 111, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 117, 81, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -37, 127, -43, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -44, 127, 127, 127, 127, -128, -58, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 12, -128, -112, 127, 127, 96, 59, 69, 80, 127, -49, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -27, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 18, 127, 127, 127, -128, 127, -49, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -55, -128, -128, -29, -128, -128, -128, 127, -128, -128, 127, -128, 26, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 78, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -117, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -127, -128, -128, -64, 127, 127, 127, 127, 127, -113, -128, -128, -128, -128, -128, -128, 127, 127, -128, -123, 118, -128, -128, -128, 127, -128, -128, 127, -69, 127, 127, 127, -117, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -13, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 102, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 55, 29, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -74, 102, -127, 127, 127, 127, 127, 127, -85, 3, 127, 109, -128, 127, 127, 127, 127, -128, -128, 37, -128, -128, -128, -5, -128, -128, 127, 127, -128, 121, -128, -128, -128, -128, -128, -74, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -17, 127, 127, 0, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 32, 127, 127, 127, 127, 127, 127, 127, -128, -128, 3, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -36, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -76, 127, 103, -128, -79, 127, -128, -128, -128, -128, -128, -128, 127, 113, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -97, 127, -128, 127, 127, 127, 127, 21, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -80, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -48, 92, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 93, -111, 127, -124, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 112, -128, -128, -128, -128, -128, -128, -128, 48, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -114, 86, -128, -91, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 96, 127, 127, 127, 127, -128, 86, -128, 127, -128, -128, -85, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -55, 5, -128, -128, -128, -128, -128, -128, -128, -128, -21, 3, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 45, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 52, -128, 127, 91, -128, -128, -113, 127, 127, -128, 127, 127, 127, -128, 3, 127, 127, -128, 127, 127, -107, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 63, 127, 39, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 52, -128, -128, -128, -128, -128, -128, -128, 127, 80, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 103, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -36, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -68, 127, 127, 127, -116, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 63, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -73, -50, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 5, -128, 127, 127, 114, 127, 127, 127, -128, 127, -128, 57, -50, 127, 127, 127, -128, 69, 127, 127, 10, 127, 127, 127, 127, -128, 127, 127, 127, -79, -128, -128, -128, -128, -128, -128, -128, -128, 16, -128, -128, -128, -128, -128, 127, 58, -128, -128, 127, 103, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 29, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 24, -63, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -44, -128, 127, 127, 85, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -118, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 75, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 123, 127, -128, -128, 127, 127, -60, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -117, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 43, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -29, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -6, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 76, -128, 127, 127, -128, 127, 127, -128, -103, 127, -128, -128, 127, 127, 127, 127, 127, 64, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -85, -128, 127, -128, 127, 127, 127, 78, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 47, -75, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 29, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -33, 127, -128, -128, 85, 54, -75, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -13, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -2, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 36, -112, 127, 127, -128, -128, 127, 127, -3, 127, 127, 127, 127, 127, 127, 127, -128, -128, 32, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -63, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 88, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -54, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -11, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -78, 127, 127, 127, 127, 127, 127, 127, 79, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 93, 70, 127, 127, 127, 127, 127, 127, 127, -33, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -13, -128, -128, -10, 127, 127, 127, -128, 127, 127, 127, 53, 127, 127, -128, -128, -128, -128, -128, -128, 127, 31, -128, -122, -107, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -28, -128, 127, -128, -128, -128, 1, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 121, -128, -128, -128, -128, -128, -49, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 64, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 60, 127, 127, -128, 127, 39, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -44, -128, -109, 127, 127, 127, 127, 127, 127, 127, 127, 17, -128, 127, 127, -128, -128, -128, -128, -128, -128, -11, 127, 127, 127, 127, -128, -128, -128, -128, 0, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -13, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 57, -47, 127, -128, -128, -128, -128, -128, 31, -128, 52, 17, -49, 127, -128, -128, -128, 127, 127, 0, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 42, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -101, -24, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 117, 127, -128, 127, 75, -128, -128, -128, -128, -128, -128, -128, 107, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -103, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 118, 127, 127, 127, 127, 127, 33, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 109, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -44, -128, -128, 127, -128, -128, -128, -48, -128, -128, -128, -86, -128, -128, -128, 127, -128, -128, -128, 1, -32, -128, -128, -128, -128, -42, 127, 127, 127, 127, 127, 127, 74, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -113, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 1, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -43, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 111, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -7, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -73, -109, -128, -128, 127, 127, -128, 127, 127, 127, -66, 127, -128, -128, -128, 13, -128, 118, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 63, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 53, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 57, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 86, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 47, 90, -128, -95, 127, 127, -128, -113, -96, -128, -128, -128, -128, -128, -44, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -106, 127, -39, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -59, 127, -128, -128, -128, -128, 70, 127, 127, 127, 127, 127, 127, -128, -128, -45, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -80, -128, 127, 127, 73, -128, -128, -128, -128, -128, -128, -128, -128, -123, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 31, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -18, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -109, -128, -47, -128, -128, -128, -128, -128, -128, -128, -34, -128, -128, -128, 127, 127, 127, -59, 127, -128, -116, -128, 1, -128, 127, -128, 127, 127, 127, 127, 127, 85, 127, -128, -128, -128, -128, -128, -128, 92, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 66, -128, 127, 127, -49, 127, 127, 127, 127, 127, 127, 127, 127, -128, 58, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -73, 127, 127, 127, 127, -128, 43, -128, -128, -128, 127, 127, 127, 127, 127, 127, 3, -63, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 49, -128, -128, 127, 127, -128, -128, 54, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -116, -128, -128, -128, -128, 55, 127, 127, 127, -128, -128, 86, -128, -128, -97, -128, -128, -128, -128, -128, -5, -128, -128, -128, 44, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -45, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -38, 127, 127, 127, 121, -128, -128, -128, -128, -76, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -49, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 109, -128, -86, 127, -128, -128, -128, -128, -128, -96, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -69, -128, -103, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -16, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -76, 127, -128, -128, -128, -128, -128, -128, -128, -128, -109, 127, -128, 127, 81, 127, -128, -128, 127, 18, -128, 127, 127, -92, 127, -31, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -96, -128, -128, -128, -128, -18, 127, 127, 127, 45, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -71, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -68, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 50, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -85, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 34, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -34, 127, 127, -128, -53, -128, -128, -128, -128, 127, 127, 57, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -102, 127, 127, 127, 127, 127, 127, 7, -128, 127, 127, 127, 127, 127, 127, 127, -128, 45, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -80, -128, -128, 127, -128, -118, -128, 127, -128, 45, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 91, 127, 127, 127, 127, -49, 127, 85, 6, -128, -128, -128, -128, -128, -128, -91, 127, 127, -123, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 109, -128, -128, 127, 127, 127, -128, 113, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -50, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 29, -128, -128, 127, -128, -128, 127, 127, 49, 127, -128, -128, -69, -128, -128, 127, -66, -128, -128, -92, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 98, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 70, 127, -128, 127, -128, -37, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -34, -128, -128, 127, 127, 127, 127, 57, -128, -128, -128, 127, 127, 127, -128, 127, 127, 76, 127, 127, 127, 63, -128, -128, -128, -128, -128, -128, 88, -128, -128, -128, -128, -128, 103, -128, 127, 127, 127, -123, 127, -128, -128, -128, -128, 12, 127, -128, -128, 127, -128, 127, 127, 58, -128, -128, -128, -79, 127, 127, 127, 127, 127, 127, -52, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -100, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -29, -128, 127, 127, -128, -128, -128, -128, -128, -128, 0, -11, 127, -128, 106, -128, 127, 127, 127, -128, 127, -128, 127, 127, 123, 127, 127, 127, 127, 127, 127, 127, 52, -128, -124, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 73, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 78, -6, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -113, -112, 127, -128, 127, -128, 127, -128, -128, -5, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -102, -128, -128, 127, -128, -128, 127, 127, -128, -128, 86, -55, -128, 97, 127, 127, 108, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -15, 127, 127, -128, -128, -128, 127, 127, -116, -128, -28, 127, -128, 127, 127, 127, 127, 127, 127, 127, 24, 127, 127, 127, 127, 127, 127, 127, 127, 124, -128, -128, -47, -128, -128, -128, -128, -128, -31, 127, 127, 127, 127, 127, -128, -128, -122, -128, -88, 127, -128, -128, 93, 127, 127, 127, 127, -128, -128, -128, -90, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -80, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -103, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -114, -24, -128, 127, 127, 127, -128, -57, -128, -128, -128, 127, -124, 127, -128, -128, 127, 127, 127, 53, -128, 80, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 24, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 2, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 85, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -36, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -49, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 95, -128, -128, -128, 76, -128, -128, -128, -128, -128, -128, -29, 127, 127, -128, -128, -128, -128, 127, 127, 127, 79, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -75, -128, -128, -128, -128, -128, -128, 55, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 38, 3, 127, 127, -128, -128, 127, -26, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 60, 127, -95, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -24, 127, 127, -128, 127, 127, -6, 127, 127, 127, -79, 127, -128, 127, 127, 127, -78, 127, 127, 127, -53, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -59, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 44, -128, -21, 127, -128, -128, 13, 52, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 45, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -32, -57, 127, 90, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 29, 74, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -63, -23, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -53, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 100, 78, -128, -50, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -122, -128, -128, -128, -128, -128, -128, -128, -18, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -32, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 23, -128, 127, 127, -128, -128, 127, -128, -128, 127, 103, 127, 127, 127, -24, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -55, -128, -128, 127, 127, 127, 127, 127, -128, -128, -108, -128, -128, 127, 127, 127, -128, -96, -128, -2, -128, -128, -128, -128, -128, -128, -128, -128, 43, -128, -128, 15, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -21, -128, 23, 127, 127, 60, 22, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 37, 127, -128, -128, -128, -128, -128, -87, -128, -128, -128, -128, -128, -128, -128, -128, 69, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -80, -128, -128, -128, -81, -68, 127, 127, 127, 127, 127, 57, -128, -128, 127, -128, -128, 127, 50, -128, 127, 127, 73, -128, 127, 127, -128, -118, 88, -128, -128, -128, -128, -128, -128, 70, 127, -128, -128, -128, -128, 21, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -34, -128, -128, -128, 38, -128, -128, 127, 127, 127, 127, -73, -128, -128, -128, -128, -128, 127, 127, 127, -71, 127, -128, -128, -128, -128, 127, 127, -128, -128, 113, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 124, -128, -128, 123, -28, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -76, 127, -128, -128, 127, 127, -128, 50, 127, -128, -128, 127, 127, 127, 127, -123, -86, -128, -128, -128, 127, -114, -128, -128, 127, -128, 127, 127, 127, 127, -128, -90, -128, -128, 127, 127, 127, -128, 127, 127, 127, 122, 78, -128, -128, -128, -128, -128, -128, 127, 127, 127, -121, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 95, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 102, -128, -34, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -121, 127, -128, 127, 127, 127, 127, -128, 127, 127, 118, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -97, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 55, 3, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -71, -74, 127, 10, -128, 127, 127, -128, 127, -128, -128, -128, -75, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 24, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 112, -128, -128, 127, 127, 127, 31, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -3, -128, -128, 127 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
