-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            -13, -13, -3, -2, 2, -3, -9, 17, -1, 14, 2, -20, -20, 14     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( 41, 36, 66, -33, 119, -21, -55, -6, 75, 76, 14, 84, -90, 54, 17, -24, 105, -34, -79, 42, -90, -19, -32, 101, 9, 81, -20, 51, -124, 84, 18, -52, 98, 28, 57, 110, -19, -99, -84, -119, 33, 5, 119, 17, -44, -3, -16, -119, -61, -56, 124, 19, 71, -52, 110, 26, 105, 67, 124, -18, 42, 22, 51, -99, 79, 114, -62, -56, 25, -80, -88, 75, 68, -36, 49, 31, 60, 67, -12, 118, 9, 75, 111, 65, 15, -2, 37, -27, 15, 36, -99, 77, -88, 91, 13, -32, 2, 56, -45, 44, -100, -52, -109, 38, -114, 6, 0, -127, -117, -99, -26, 88, 110, -83, -110, 104, 70, 15, 114, 80, -6, -123, -87, -49, -77, 16, -74, 19, 95, 59, -74, 78, -61, 100, -117, -110, -115, -16, -90, -106, 80, -43, -36, 35, -81, -51, 31, 52, -18, 17, 111, 121, 107, 62, -123, -100, 111, 92, 45, 56, 105, 84, -52, -26, -74, 68, -69, 31, 60, -4, 55, 49, 107, 85, -51, 16, 54, 99, 92, 99, -40, 124, 19, -14, 19, -25, -101, 107, -4, 41, 88, -109, 7, 112, -13, -40, 103, -37, 127, -119, -76, -56, -75, -77, -127, 57, -36, -20, -23, 95, 91, 90, 47, -107, -117, -101, -52, -2, -77, 85, 7, -113, 43, 31, -82, 119, 105, 35, -104, -119, -19, 86, 55, -57, 76, 57, 33, 70, -22, 48, -29, -126, 91, 76, 29, -61, 14, 27, -25, 29, 119, 60, 112, 79, 80, -94, 90, -92, 48, -113, -88, 117, -21, -41, 74, -18, 101, 1, -79, 9, -36, 6, -73, 38, -113, 8, 37, -121, -24, 28, -39, 29, 64, -44, -65, -17, 72, 36, -55, -25, -95, 115, -54, 108, 21, 43, -87, -74, 10, -58, -62, 95, 28, 65, -116, 59, 53, 6, 47, -17, 48, -2, 3, -50, 9, 15, 74, 122, 107, -74, -85, -60, 103, 121, -61, 105, -42, -49, -115, -38, 109, -88, 28, -53, -116, -103, 81, 49, 98, 120, 71, 46, 88, -92, 28, -92, -83, 62, 108, 42, 99, -85, -92, 6, 80, -13, -12, -76, -14, 54, 103, -87, -72, 124, 61, -62, 33, 22, 67, 27, -36, 59, -10, -38, -21, 6, 89, 1, 40, 71, 79, -68, 1, -72, 9, -100, 89, -128, 9, 113, 20, 95, -4, -1, -61, -61, 35, 44, 95, 0, 51, -1, -23, 65, 67, -25, 2, -90, -6, 53, -61, 66, 81, -121, 3, 43, -94, 69, -95, 29, -109, 123, -4, 106, 44, 2, -76, 56, 97, -3, -5, -52, 110, 103, -121, -91, -59, 91, 9, 120, -69, -97, -42, -108, -69, -33, -87, 53, -3, -112, 87, -101, -50, -22, -95, 73, 97, 35, 74, 124, -39, 88, -16, -96, -125, -81, 49, 88, -56, 111, 59, 10, 64, -70, 46, -39, 60, 104, -24, -125, 70, -28, -122, 66, 125, -109, 104, 104, 62, 61, -125, 18, -121, 78, -77, -124, 114, -72, -69, -96, -110, -23, 2, 11, 75, -50, -63, 103, 111, 93, 45, 26, 45, 118, -4, -1, -115, 45, 112, 66, -90, -18, -86, -2, 26, 7, -43, 25, 63, 67, -122, 13, 113, 95, 126, -9, 85, -108, -52, -59, 59, 91, 127, 28, 40, -48, -99, 63, 46, -122, 10, 113, 61, 57, -109, -92, 13, 103, 76, -52, -35, -67, 93, -14, 2, -22, -43, 8, 4, 37, 37, -88, 94, 70, -77, -87, 127, 39, -45, 115, -78, 110, -105, -46, 51, 2, -29, -63, -122, 22, 40, 84, 127, -16, 9, 49, 25, -96, -89, -50, 29, -106, -8, 126, -13, 125, 88, 48, 56, -30, 104, -13, 118, -95, 125, -81, 69, -128, -100, -48, 85, -21, 75, -60, 63, 112, 79, 37, 105, 105, -79, 75, -128, 102, -35, -98, 19, -97, -121, 72, -32, 77, 95, -74, -26, 77, -83, 111, 36, 5, -75, 110, 118, 51, -44, -86, -122, 39, 88, 78, 55, 102, 32, -64, -97, 120, -89, -16, 58, -15, -22, -81, -10, 85, 121, 70, -14, 57, 21, -112, -43, 101, 58, -86, 88, -121, 55, -9, 12, 68, 25, 116, 55, -104, 121, 70, 19, 43, -103, 60, 95, -111, 93, 111, 32, 127, 8, -14, 16, 83, -48, -125, 111, 105, 95, -107, 48, 57, 17, 100, 32, 5, -119, -65, -98, -75, 56, -106, -43, 68, -93, 5, 88, -62, 22, -48, -96, 106, -14, -67, 126, 52, -103, -3, -61, 87, -70, 89, 102, 67, 127, -15, -36, 37, -106, 76, -6, -30, 68, -113, -60, -58, -79, -2, -6, 38, -64, -77, 98, 103, -108, -56, 53, -78, 58, 107, 79, -53, -30, -90, -20, 56, 79, -77, -75, -17, 5, 116, -12, 92, 63, -12, -17, 8, -109, -40, 56, -32, -31, 33, -86, 67, 57, -50, 60, 41, 75, 93, 61, 117, 38, 104, 36, 44, 11, 19, -21, -123, 17, 3, 12, 4, -61, -62, 65, -8, 37, 36, -20, -12, -80, 115, 103, -111, 103, 43, 123, -65, -95, -31, -63, 11, 7, 125, 62, 110, 101, 74, 109, 120, 94, -117, 26, 12, 40, 70, -1, -89, -27, -112, -82, 110, -101, -27, -126, -35, 67, 69, 32, -22, 70, -114, -107, 56, 19, 12, -57, -28, -48, 99, -48, 65, -77, 5, 102, 50, -116, 77, -4, 107, -87, 62, -87, 83, -66, -67, 118, -14, -40, 78, 94, 33, -7, 8, -127, 102, 30, 113, 17, 29, -21, -120, 43, -114, -36, -99, -83, 59, 94, -95, -122, 46, -82, 50, -61, 58, -54, -111, -49, -117, -4, -56, -30, 71, 113, 93, -20, 112, -51, 57, 26, 121, -113, 122, 91, 36, 65, -27, -46, 28, -60, 31, -105, 23, 19, -12, -1, 52, 37, -69, 11, -106, -81, -93, 19, -85, 6, 11, 55, -20, -68, 6, 53, 119, -106, -116, -13, 37, 44, -106, -36, 41, 113, 126, -73, 22, -86, 23, 46, -108, 27, -8, 54, -48, 82, -22, 15, 85, -3, -99, 77, -103, 51, -46, -85, 66, -11, 107, -116, 13, 57, -53, -93, 121, -128, -19, -20, 68, -88, -35, -87, 104, 19, 5, -94, 52, 4, 68, 81, 10, -24, 112, -45, 35, 76, 9, -90, 18, -34, -58, 85, -43, 81, -33, -120, -112, 49, -6, 81, -64, -81, 96, -37, 97, 41, 96, -22, 40, -85, 0, 20, -60, 101, -49, -99, 33, -68, -10, 33, -59, -112, 86, 86, -17, -4, 116, 83, 10, 111, 96, 77, -54, -67, -19, 83, 44, -53, -128, 39, -17, 64, -58, -63, 127, 101, -29, -64, -98, -33, -57, -127, 122, -8, -113, 112, -41, 48, -76, -85, 4, 58, -20, 26, -12, -120, 60, 115, 87, -24, 125, 108, -118, 9, -6, -103, 85, -111, 117, 10, 90, 31, -69, -66, 80, 117, 112, 57, 103, -57, -67, -126, -60, -17, 111, 40, -101, 90, 99, -12, -112, -34, -87, -48, -67, -127, 25, -121, 67, 23, 114, 62, 113, 104, 102, 126, -101, -106, 60, -108, 54, -116, 114, 93, -50, -110, 20, -105, -45, -84, 60, -57, 41, 126, 110, -110, -5, 72, -42, -8, -126, -50, 110, 106, 64, 44, -53, -16, 106, -15, -111, 64, 94, -25, 32, -104, -63, 20, 65, -23, -69, -117, 101, -20, -70, -17, 97, 43, -84, 101, 10, -2, 56, 61, 126, -25, -72, -77, -55, 102, -66, 15, -106, 123, 107, 34, -47, 15, 17, 84, -116, 48, -48, 94, 20, 69, -51, -125, -51, -120, -95, -4, -115, -46, -115, 64, 30, -105, -79, -9, -93, 45, 95, -106, -54, -5, -96, 41, 44, -88, 84, -100, -83, 123, 28, -105, 4, -111, -123, 42, -15, 28, 22, -91, -38, -74, 35, 2, 1, -109, 41, 12, -79, -105, 57, 74, -122, 8, -118, -90, 104, 57, -48, 51, 52, -68, 10, 122, -70, 79, -24, 113, 55, 120, -109, -70, 81, 80, 12, -4, 76, -99, -106, -82, 68, -105, -3, 5, 4, 121, 52, -30, -88, -118, -121, -88, -20, 1, -59, -103, 108, 42, 111, -23, -118, -15, -65, -18, 75, -63, -63, -64, -117, 47, 31, -111, -85, -117, 99, 47, 37, -37, -6, 102, -98, 127, 67, -105, -90, -95, -40, -64, 101, 39, 127, 124, -26, 41, 36, -75, -9, 99, -54, 2, -115, 45, 15, -60, -70, -39, -32, 121, -40, 79, 105, -39, 26, 106, -121, -56, -82, 92, 48, 17, -105, 12, -83, -73, 85, -8, -74, 34, -43, -13, -86, 16, -17, -96, 49, -110, 78, -57, -89, -28, 57, 19, -115, 72, 74, 111, 84, -51, -37, -83, 101, -77, 45, -42, 61, -56, -86, -65, 80, 107, -41, 16, -105, -103, 16, -77, -75, 43, 118, -85, -71, -28, 36, -52, -76, 116, 81, -102, -105, 96, -126, -126, 94, -101, 38, -1, -12, 66, -107, -117, -87, -101, 10, -122, 57, -52, -25, -70, 70, 26, -72, 59, 32, 56, 114, -58, 101, 63, -116, -92, -95, -66, -69, 99, 27, 80, 73, 84, 76, -85, -39, 40, 51, -98, 17, 111, -78, -38, -23, 61, -102, 28, -101, -69, -40, -14, -103, -98, -12, -112, 55, 103, 50, 44, 24, 4, -25, -28, 26, -104, 109, -6, -50, -62, -72, -37, 69, -3, -84, 32, -88, -29, -40, -105, -15, 115, 52, 5, 34, -41, 122, 61, 60, -29, -114, -89, -85, -17, 59, 74, -67, -29, 40, 19, -44, 62, -72, 63, 3, -44, -117, -73, -58, 64, 24, -56, -10, 115, -105, 91, 42, 5, -121, -84, -64, 6, 49, 20, 65, 69, -11, -57, 115, 91, -93, 91, 89, 116, 64, -62, -2, -89, -100, -118, -92, 79, -81, -34, 91, -77, 106, -61, -60, -110, -45, 75, -23, 52, 11, 105, 104, -75, -27, -18, 110, -1, 87, 76, -39, 70, 119, 70, 32, -66, -64, 103, -12, 40, 81, -22, 46, 76, 80, -59, 47, -36, -98, -100, 28, 104, -32, 98, 110, 123, -100, 37, 41, -50, 92, 22, -20, 65, -99, 94, 49, 72, 0, 54, -42, -74, -32, -39, 125, 66, 112, -44, 118, -112, 61, -60, 68, 73, 112, -99, -99, 89, -38, -17, 108, 10, 26, -76, -75, 78, -10, 64, 91, -1, 39, -24, 53, -124, 45, 113, 13, 77, 46, 60, -19, 72, 78, 25, 40, 0, 45, -119, 16, 16, -128, 75, -115, 11, -15, -45, -81, -122, 61, 18, 100, 47, 95, -1, -100, 78, 20, -101, -50, 86, 63, -122, 103, 35, 70, -11, 101, -41, -67, 62, 36, 32, 122, -35, 55, 78, 59, -48, 118, -103, -66, -112, -13, -47, -12, 108, -76, 57, -42, 125, -37, 36, 60, -112, -115, -41, 125, -109, -65, 96, -85, -29, 43, -87, 32, 35, 76, -102, 46, 124, 26, 111, 70, 47, -51, -91, 20, -65, 99, -23, 76, -123, 43, 77, -63, -40, -56, 87, 43, -81, -126, -124, 104, -127, 124, -104, 94, 48, -20, -32, -1, 8, 73, 114, 22, 88, -78, -85, 71, 85, 71, 75, -73, -107, -21, 124, -13, 24, -31, 98, 8, -50, -27, -102, 123, 117, 87, 80, 64, 74, 59, -73, -1, -69, 34, 23, -112, -81, -109, 95, -33, -50, -109, 22, 120, 19, 47, -123, -108, -63, 32, 10, 12, -26, 74, -99, -23, -11, 118, -66, -34, -46, -68, 119, -46, -3, 118, 90, 95, -61, -2, -63, 121, -10, 55, -27, -113, 87, 71, 16, 44, 82, 99, -64, -22, 117, -5, -39, -114, 7, 79, -122, -122, 104, -74, -15, 9, -113, 53, 30, 61, 114, 59, -23, -7, -10, -97, -97, -55, 118, -7, 3, 85, -87, 92, 127, 110, -14, -37, 83, -45, 16, -29, 34, -81, -64, -89, 44, -70, -54, 29, 12, -89, 98, -27, 15, -31, -25, -16, -101, -52, -90, -71, -47, 18, -62, 47, -18, -13, -102, 54, -65, 62, 32, -62, -41, 50, -77, -81, -32, -54, 38, -59, -91, 113, 87, -12, -72, -14, -47, -128, 63, 50, 99, 14, 40, -68, -103, 91, -19, 81, 88, 115, 28, -71, -21, 32, -52, 116, 11, 40, -115, -24, -127, 86, -60, 120, -82, 127, 35, -31, -110, 29, 124, -66, 28, 118, 17, -3, -12, -47, -36, -102, -31, 68, 27, -111, 48, -93, 29, -76, -15, -40, 111, -82, -119, 97, 61, 51, -47, -51, 106, -40, -76, 87, 112, -62, 32, -46, -16, -109, -119, 31, -103, 25, -19, -126, -68, -58, -88, -75, 28, 106, -108, -107, 71, 5, 58, 36, 16, 35, -70, 24, 66, -60, -26, 78, 41, 36, -87, 124, 31, 68, -9, -125, 42, 62, -95, -57, -96, 13, 114, -46, -22, -111, -50, -115, -51, -55, 110, 78, -122, -97, -6, 46, -21, -80, 89, 53, 35, -82, 126, -113, -109, -33, 91, 64, 38, -18, 98, -92, -69, -78, 17, 124, -30, 120, -61, -91, -89, -63, 43, -103, 3, 36, 49, -32, 96, 121, 44, 27, -7, -10, -47, -22, -123, -67, -65, -58, -121, -118, 42, 94, 32, 122, 111, -107, -41, 121, 1, 46, 126, 45, -77, -94, -17, 87, 53, 61, 8, -50, -82, -26, 121, 19, 9, -54, -51, -96, -70, -41, 44, 88, 70, -20, -1, -120, 3, -88, 19, 17, -100, -54, -60, -119, -17, -5, 76, -79, -28, -53, 48, 85, -93, 10, -115, -64, -125, -120, 110, 57, 21, -83, -51, 91, -3, 14, 26, -66, -12, -29, 121, -9, 115, 7, -65, 35, 117, -57, 91, -36, 40, -117, 49, -65, 120, 20, -39, -15, 83, -68, 7, -46, 111, 115, -95, 112, -67, 127, -58, -92, 32, 101, 16, -115, -125, 28, -110, 96, 99, -47, -36, 61, 60, 31, 90, -83, -113, 2, 46, 6, 83, 17, -58, 99, 82, 93, 36, -78, 108, 58, 110, -60, 79, 5, 59, 92, 41, 83, 103, -95, 41, -21, -47, 31, -67, -126, 40, 54, -17, 50, 39, 8, 106, -56, -13, -41, 77, -78, 124, 97, -113, 47, 101, 71, -9, -42, 29, -76, 103, 95, -91, -75, 102, -128, 62, 30, -80, 72, 6, 104, 113, 23, 47, 55, 122, -18, -84, 62, 21, -31, 116, -54, -111, 36, 20, 4, -69, 120, 118, -88, -41, 29, 59, 53, 89, -67, 3, -9, -29, 24, -31, -111, -88, 18, -100, 33, -60, -32, -117, 98, -42, 123, -73, 112, -87, -93, 72, -83, 109, -87, -40, -27, 21, 34, -110, 23, 87, 62, 88, -68, -36, 26, 82, -2, 102, 25, 41, -11, 7, -112, -53, 34, -17, -66, -47, 4, 18, -53, 122, -87, 19, -118, 73, 108, 3, 55, -96, -112, 56, -66, -30, 102, 112, 62, 35, 80, -56, -27, 109, 52, -111, -13, 36, -117, 50, -122, 76, -114, 21, -49, 5, 79, -113, -91, -30, -72, -56, -117, -87, -116, -108, -26, 22, -48, 1, 43, 58, 92, 31, -124, 57, -67, 102, -29, -28, 30, 17, 96, -53, -87, -1, 98, -80, -5, -109, 30, 122, 127, 124, -33, -38, -91, 13, 101, 56, -111, -75, 85, -117, -58, -100, 20, -56, -21, 90, 99, 118, -60, 72, -91, -86, -48, -123, 55, 111, -26, -45, 29, 17, 45, -12, -44, -6, -63, 94, -51, 94, 27, -109, -79, -81, 44, 6, 49, 125, -112, 4, -31, -37, 9, -35, -47, 101, -90, 105, -117, -127, -13, 116, 90, -25, 38, 73, -22, 54, 51, 37, -26, 108, 17, -119, -97, 87, 124, 5, -94, 8, 41, -109, -105, 126, 100, -76, 17, -27, 33, -7, -7, 46, -87, -57, -92, 14, 63, 109, -8, 64, -106, 115, -86, -82, -43, -91, 85, -117, -13, 77, 0, 10, 86, -37, -1, -107, -26, -27, 10, -27, 11, -38, -95, 44, -48, 52, -123, 9, 106, 73, 9, 78, 100, 51, 78, -58, 65, -21, -31, -99, -123, -46, 66, -122, -19, -117, -11, -7, 126, -33, -111, 44, 127, 42, -94, -59, -95, -105, -9, -114, 121, -3, 3, -56, 125, -120, 48, -74, -45, 36, -40, 38, 27, 0, -51, -38, 69, 78, -14, -88, 83, 97, -42, 65, -42, 106, 108, -126, -64, 49, -119, -49, 50, 93, 38, 66, -120, 84, 101, -101, -58, 0, 27, 98, -72, 55, 91, 108, 110, -119, -124, 76, -29, -112, -91, -120, -36, -124, -128, 93, 19, -89, -27, -33, 126, 85, 46, 54, 105, 73, -104, 122, -107, 71, -22, -27, -84, 39, -52, -84, -49, -27, 105, -87, 67, 114, -124, 47, 33, -14, -12, 126, -107, -121, 126, 71, -76, -80, 2, -96, -41, -63, 37, -117, 30, 18, 10, 60, -116, -72, 46, -42, 24, -92, 28, 4, 81, 70, 21, 69, -16, -71, -53, 111, 27, -31, -92, 35, 62, 95, -112, -106, 57, 8, -125, 21, 113, -128, -1, 53, 77, -1, -5, 103, 24, -63, 38, -52, -54, -118, 12, -111, 79, -24, -80, -6, 63, 6, -82, -70, 91, -67, -79, 39, 88, -49, -10, -71, -23, -47, -67, 22, 11, 21, 73, -112, -73, -50, -94, 93, -96, 97, -85, -25, -57, -128, 97, 104, -122, -74, 84, 118, -77, 39, 42, 95, 118, -5, 59, 126, 49, -107, 70, 22, 102, 17, -74, -7, 78, -87, 105, -32, -74, 103, -11, 95, -112, -46, -51, -2, 83, 65, -86, 48, -45, -36, 3, -87, 101, -64, -72, 76, 53, 39, 69, -7, -112, -60, 80, 78, 8, 60, -89, 2, 57, -84, 127, 107, -101, -70, -124, 114, -55, 118, -16, -29, 101, -16, 26, -12, -96, -89, 61, -75, -18, -23, -5, 100, -31, 119, 15, -99, 104, 59, -29, 5, 59, 4, -81, 89, 83, 39, -28, -98, 32, 25, 71, -52, 27, 40, 54, 49, 10, -97, -92, -103, 73, -118, -101, -100, 36, 5, -101, -24, -30, 61, 32, -87, -38, -95, 11, -69, -114, 21, 16, 56, -87, -107, -29, -17, 46, 118, 88, 19, 69, 92, 75, -107, 108, -12, -123, -89, -94, -16, 72, 111, -53, -77, -116, -48, 70, 5, 96, -17, -120, 20, -26, 91, 70, -39, 4, -121, 22, -82, -88, -102, -67, 118, -70, 98, -28, -37, -113, 16, 58, -119, -92, 121, -44, 57, 85, 126, 0, -67, 59, -1, 4, -123, 55, 65, 117, 90, -116, 113, 66, -96, -88, -23, -107, 49, -85, 54, -73, -33, -66, -18, -12, 0, 39, 4, 5, 109, 114, 73, -89, 101, 121, -112, -107, -116, 100, -12, 22, -93, -69, 92, 98, 21, 48, -4, 19, 110, 65, 73, 58, -86, -19, 66, 102, 99, 119, 76, -102, 65, 79, -116, -7, -120, -4, 111, 104, -73, 76, -110, 10, 93, 0, -106, 8, -61, -122, -51, 35, 12, 69, 102, -34, 46, -126, -92, -115, 89, -37, 20, -112, -57, -113, 57, -68, 34, -73, -124, -89, -32, -81, -30, 28, -91, 23, -119, 6, -73, 103, -70, 67, -115, 89, 53, 45, 33, -117, 30, 63, 14, -41, -114, 80, 47, -86, -49, -89, 41, -95, -71, 101, 110, -42, 119, -107, 118, -110, 107, 19, -25, 52, 88, -112, -47, -42, -94, -125, 110, 75, -79, -112, 25, 106, 20, -111, 35, 41, -101, 83, -115, 20, -126, -71, 42, 8, -5, -128, -92, -6, -104, -82, 45, 122, -12, 25, 82, 74, -10, 6, -60, 21, 105, 31, 115, 111, 57, 99, -1, 66, -16, -119, 19, 65, -78, 46, -79, 108, -77, 26, -83, -16, -25, -6, 33, 67, -115, -34, -118, 13, 21, 20, -47, -72, 123, -70, 32, -78, -22, 8, -29, 39, -1, 20, -2, 7, -67, 25, -69, 126, -5, -87, -75, 56, -87, -106, 31, 95, -117, 41, 110, -90, 81, -70, -56, 73, -119, -79, -126, -45, 111, 45, -79, 37, -59, -88, -80, 85, -112, 26, 79, -106, 71, 82, 115, -76, 104, 99, -41, -10, 56, 114, 33, -19, 70, -25, 47, -57, 109, -21, -32, -122, -61, -90, 56, -25, 12, 127, 75, 113, 17, 31, 26, -9, 107, 95, -16, 125, -16, -29, -10, 32, 7, -57, -36, 1, -44, -57, -82, -58, -96, -56, -73, -116, 98, -127, 122, -104, -12, -80, -112, -5, 51, -98, 80, -63, 107, 51, 67, 36, 89, -16, 23, 101, -79, -30, 56, 49, 38, -115, -121, 121, 85, -91, -86, 123, -96, -43, 53, 101, 46, -35, 85, 101, 7, 121, -12, 49, -66, 75, 5, 57, -124, 98, -86, -87, -47, -75, 93, 7, -18, 34, 60, -79, 78, 24, -66, -58, -54, 51, 21, 115, -54, 38, 113, -53, -107, 45, 22, -96, -128, 123, 45, 48, 45, 109, 92, -89, -74, 89, 91, -112, -96, 4, 105, -94, 126, -109, 82, -119, 36, 124, 126, 115, -16, -60, 1, 52, 83, -96, 61, 7, -106, 94, 91, -77, -75, 110, -51, 16, 38, -14, 55, -72, 75, -41, -16, 58, -37, 80, -61, 41, -42, -114, -116, -2, -32, 108, -99, -58, -12, -53, -44, -70, -45, -34, -111, -104, -47, 29, 15, -81, 44, -13, 118, -58, 78, -47, 77, -100, -18, 14, -83, 81, -52, 83, -91, 86, -19, -27, -64, 18, -12, -112, 93, 92, 110, -24, 93, -93, 5, -83, -75, -116, 105, 111, -120, 114, 44, -77, 91, -22, -98, 112, -73, 84, -39, -2, -10, 29, -53, 30, 10, 103, 20, -70, -89, 84, 58, -84, 17, 25, -12, -120, 106, -67, -125, 58, -25, 6, 36, -116, 80, 24, 22, -56, 48, 102, 50, 51, -23, -126, 75, -94, -88, 118, 36, 23, 69, -125, -121, -1, -99, 11, 59, -79, 96, 85, 105, -61, 110, -82, 6, -17, -77, -87, 10, 116, 7, 123, -70, -70, 55, -9, -81, 15, -23, 80, -19, 38, 6, -93, -79, -104, -82, -80, -74, 65, 108, -53, 82, 48, -78, -57, 17, 103, 77, 62, 99, 125, -4, 108, -14, 101, -78, -70, -110, -103, 89, 86, 108, -125, 98, -76, 110, -121, 108, -87, 36, 38, 0, -41, -126, 80, 85, -83, 29, 113, 118, -99, -114, 75, 41, 96, -59, -35, 7, -109, -121, 21, -55, -104, -58, 3, -116, -44, -78, 117, 77, -23, -22, -33, 0, 55, 124, 118, 93, -64, -41, 64, 53, -58, 40, 25, 51, -14, -12, 31, -121, -109, 17, 89, 73, 23, 9, -57, 66, 28, 116, -80, -101, -24, 87, 1, -109, -51, 19, -30, 75, -56, -89, -67, 14, -84, -53, -115, 12, 91, -112, 107, -14, -3, 112, 50, -51, -74, -119, -124, -95, 26, 38, -116, 65, 32, 6, -70, -128, 89, 94, 55, -84, -82, 23, 113, -25, 74, -86, -76, 45, 66, 88, 71, 78, -104, 33, -124, 22, 119, -89, -43, -4, 98, -6, 121, -122, -40, -25, 85, 99, -128, 34, 114, 88, -77, 105, 85, 36, -10, -72, -102, -10, -48, -57, -46, 125, 98, -59, -1, -86, 78, -19, 73, -4, -34, -26, -16, 124, 38, -4, 98, -102, 72, -52, 53, -88, -110, 4, -64, -9, -109, 62, 101, -75, 12, 13, 18, 112, 59, 80, -12, 124, 91, -46, -9, 51, 99, 108, -69, -20, -36, 121, 52, 21, -83, 12, 42, -77, 108, -22, 120, 59, 16, -13, 39, 91, -120, 85, -41, -78, -87, 2, 119, 77, 22, 103, 71, -51, -24, -86, 31, 63, 38, -98, 51, 1, -37, -7, -1, 105, -45, 51, 120, 87, 30, -23, 98, -48, -113, -124, -28, 92, -69, -107, -71, -88, -52, -32, -65, -78, -32, -127, -11, -103, -101, -11, 10, -15, -70, -9, -28, -87, -10, -90, 51, 5, 104, -101, -50, -42, -52, 110, -117, 60, 31, -112, -14, 102, 86, -18, 90, -97, -7, 61, 125, -54, -72, 35, -67, -103, 111, 35, 64, 21, 7, 6, -66, -29, -79, 18, 9, -3, 119, 99, -124, 83, -46, 15, -21, 55, 53, 31, 111, -87, 81, -53, 99, 115, -62, 115, -104, -72, 16, 79, -85, 83, -26, -11, 125, 51, 25, 126, 107, -90, -101, -65, 86, 121, -105, 94, 93, 125, -125, 104, 80, 91, -73, 73, -51, -25, 78, -77, -83, -33, -68, 2, -107, -97, -19, 84, 63, 4, -46, 86, -17, -128, -79, 96, 22, -74, -12, 121, 80, -33, -17, -45, -28, 120, -63, 1, -54, 41, 1, 95, -55, 54, -43, 66, 10, -109, -128, -122, 113, -83, 126, -31, 105, -9, -97, 54, -112, 108, 69, 38, -47, -90, 107, 89, -31, -43, -99, -105, -85, -16, 95, -38, 124, -28, -115, 57, 126, 110, -45, -5, 27, 107, -12, 74, -52, -108, 60, -14, 32, -69, -84, -84, 49, 33, -54, -59, 63, 86, 108, -23, -48, -72, 82, -26, 100, 114, 51, -5, 120, -79, 12, 44, -90, 31, 39, 105, -54, -126, -29, -40, 110, 98, 84, 28, 35, -29, -6, 12, 38, 21, 37, -72, 123, -125, 42, -109, 56, -44, -15, -37, -125, -18, -90, -77, -32, 74, -16, -27, -36, -51, 79, 67, -62, -68, 79, -123, 31, 55, 105, 12, 53, 34, -30, -36, 85, -61, -96, -95, 105, -2, 49, -87, 105, -50, -78, 127, 89, -80, -50, 31, 68, -7, 39, -21, 37, -87, 25, 92, 87, -3, 40, 88, -44, 66, 47, -9, 37, -36, 12, -118, 5, -119, 66, 79, 70, -40, -49, -82, 0, -6, -58, 112, -78, 29, 108, -94, -109, 39, 127, 79, 7, -42, 13, -77, 38, -107, 98, -103, -91, -60, 90, -39, 45, 124, -80, 90, -121, -99, -10, 31, 59, -18, -23, -32, -4, 64, 90, -27, 116, -83, -47, -119, -96, -44, -25, 21, 19, 56, -118, -54, -35, -58, -68, -12, -64, 14, -86, 17, -111, 26, -23, 14, -79, 45, -50, 22, 79, -125, -126, -104, -115, -77, -99, -128, -80, 0, -105, -30, -78, 92, 30, -62, 12, -26, 0, 57, -6, 54, 65, -128, -30, -126, -103, -14, 39, 21, -38, 87, -103, -115, -73, 54, -20, -61, 101, 106, -84, 10, -119, 116, -7, -37, -14, 105, 70, 52, -52, -9, -109, -47, 0, 124, 77, -27, 30, 74, -61, 19, -86, -113, -4, 97, 78, 5, 15, -31, 4, 73, 30, 60, 11, -115, -128, -14, 51, 113, 105, 88, -30, -63, 44, 73, 103, 119, -86, -60, 10, -54, 1, -92, -40, -39, 64, -3, -32, -87, -109, -63, 12, 30, -69, 100, 120, -14, 11, -42, 82, -38, -56, -38, 61, 17, -114, 38, 104, -50, -108, -46, 117, 76, -24, -3, 8, -9, -62, -107, -42, 82, -61, 116, 70, -103, -61, -21, -79, 36, 62, -44, 61, 77, -109, 13, -16, -44, -72, 81, -1, -75, 63, -82, -88, 18, -10, -108, -52, 9, 70, -82, -28, -35, 33, 47, -97, 122, 31, -79, 37, 28, -89, -61, 59, 123, 95, 68, 14, -64, 72, -122, -45, 60, 9, 82, 80, 75, -44, 93, -99, -111, -84, 35, -55, 14, -98, -93, 12, -61, 8, -40, 106, 125, -47, -25, -77, -89, -111, -47, 9, 116, 16, -64, 96, -92, 53, 120, -41, -39, 14, 25, 122, -43, -71, -53, 13, -94, -114, -24, 69, 77, -15, -52, -92, -88, 107, 3, 115, -46, 8, 41, -1, -27, -28, -115, -12, -106, 100, -24, 3, -43, -23, 92, 95, 3, 47, 30, 42, 18, 34, -122, -85, 83, -49, 81, 21, -100, 11, -43, -120, 121, -80, 82, -119, -95, 111, -100, -95, -126, 52, -82, 82, 117, 87, -3, 13, -127, 19, 57, -70, 98, -89, -20, -92, -85, -100, 23, 5, -107, -18, 121, -126, 123, -118, 52, 14, -58, 106, 15, 16, -2, 121, -87, 93, -16, 12, 101, 62, 92, 38, 30, -31, 44, -37, 107, -43, 26, -2, 101, -2, 40, -5, -33, -97, -50, -101, -11, -23, -48, -26, 109, 52, -84, -97, -107, 77, 99, 68, 105, -108, 88, 39, -1, 71, 85, 111, 50, -4, 20, 90, 95, -71, 77, 29, -125, 29, -81, -46, -26, -84, 48, -113, -34, -23, -21, -2, 45, -18, -106, -77, -39, -62, -79, 96, -23, -36, 28, -85, -19, -16, -86, -3, -95, -127, 123, 17, 47, 122, -88, 102, -83, 42, -44, -68, -31, -69, -109, -78, 70, 101, 88, -41, -119, 103, 26, -75, 42, -124, 68, 36, -37, -41, -59, 44, 85, -75, -70, 77, 106, 118, -128, -97, -121, 71, -23, 124, -71, 27, -5, -16, 99, 127, -23, 90, 38, -51, 42, -90, -57, -33, -6, 91, 1, 109, 11, -35, -40, 88, 26, 33, -14, -75, -22, -1, 59, 51, 114, -65, 89, -79, -15, -79, -55, 0, 26, 108, -49, 45, 23, 15, -22, -94, -27, -24, 76, 110, 79, 35, -82, 95, -102, -88, -16, 81, 103, -3, -113, 64, 71, 77, 36, 126, -9, 51, 85, 53, -87, -55, -34, 23, 46, -54, -87, -114, -36, -124, -42, 68, -45, 104, 113, 59, 75, -9, 15, -74, -122, 50, 112, -103, -1, -126, 55, -88, -114, 27, -70, -74, -36, -52, 107, -11, -29, 72, 17, 45, -117, 81, -48, -51, 39, -45, 43, -127, -87, -6, -39, -67, -8, -9, -99, -74, 53, 89, -71, 96, 22, -115, -3, 42, 94, -84, 32, -62, -100, -94, 95, 59, 127, -5, 10, 80, -61, -19, -75, -14, 115, 83, -8, 13, -7, 127, -104, 73, 5, 47, -9, -102, -44, -79, -49, -5, -10, -41, 20, -122, 124, -3, 112, -54, -125, 91, 51, -30, 30, 115, 32, 60, -57, 14, 64, 87, -103, 35, 104, -39, -2, 5, 91, -32, -21, 27, 12, -75, -87, -12, 62, -25, -114, 71, 11, 76, 0, -86, 2, 35, -80, -86, -56, -108, 124, 1, -84, 75, 69, -6, -110, 71, -76, 18, -15, -15, -87, 108, -106, 114, -72, -97, 68, 87, -128, 45, 74, -5, 57, -77, -77, 125, 54, 74, 108, -53, 40, -26, 10, -93, 2, -36, -72, -74, -80, 15, 75, 0, 83, -11, 43, 71, -12, -105, -100, 109, -4, 18, -34, -102, -104, 2, 71, -24, 62, -91, 16, 47, 101, 125, -67, -117, -11, -44, -114, -46, -80, -113, 34, 70, 64, 94, 21, -93, 69, -74, 33, 25, -119, 103, -95, -111, 62, -25, 28, 21, 11, -52, -22, -117, 23, -42, 33, -41, -11, 88, 59, -12, -13, -13, 23, -91, 48, 56, -21, -70, -107, 48, 65, 24, -97, -101, -63, -12, 100, -44, -70, 110, -127, -66, 102, -91, 117, -52, -118, 79, 29, -123, 93, -35, -109, 106, -4, -61, 58, 98, -49, 102, -128, -19, -8, -34, -38, -123, 39, -80, 66, -126, 0, -12, 60, -88, 35, -82, -27, -5, -54, 25, 45, -44, 87, -25, 2, 36, -109, 112, 22, -50, 11, -91, 84, -39, -78, -61, 26, -49, -27, 71, -67, -89, 87, -45, 34, 100, -38, 59, -24, -79, 57, 59, 12, 27, 9, -96, -120, 23, -126, 54, -115, 63, 51, 89, -80, -43, 66, -109, -109, 50, 70, -64, -31, -40, 100, 48, -74, 118, 110, 86, 90, 107, 67, 103, 9, -78, 92, 115, 19, -124, 84, 29, 16, 65, 2, 29, 6, 115, -47, 56, 105, 83, 98, -123, 4, 119, -21, 122, 120, -98, -114, -15, 70, 93, -64, -27, -85, -26, 92, -113, -24, 53, 37, -127, 17, 60, -114, 94, 58, -9, 19, -8, 66, -70, 82, 25, -55, 71, 90, -29, -122, 15, 10, -16, 108, -15, 26, -90, -81, 93, -10, -123, 106, 108, 68, -2, 120, 36, 92, -105, 21, -32, -1, -116, 40, -102, 80, 96, -99, -111, 71, -101, -89, -90, -49, -16, -55, -10, 121, -24, 29, -113, -13, 68, -83, 67, -61, 74, 39, -29, 84, -9, -17, -95, -16, 13, 104, 18, 98, 38, -15, 19, 26, -86, 99, 30, 107, -30, -98, 74, 34, -55, 54, 97, 2, 10, -33, 54, 101, 101, 55, -66, 88, -21, -35, -23, 119, -108, 20, -112, -24, 109, 24, 100, 30, -51, -20, 118, -74, -76, -94, -78, 117, 70, -100, 73, 82, -26, 22, -79, 32, -108, 126, 105, 106, -9, 68, 11, 68, 1, -116, -55, -116, 55, 53, -101, 81, -47, 111, 72, -120, -73, -23, 121, 30, -24, -95, -5, -89, 107, 37, 89, -124, -84, 93, -94, -101, -49, 70, -77, -38, -51, 26, -123, -8, 73, 42, 59, -79, -15, 0, -100, 19, 1, -104, -15, 54, -128, 81, 110, 98, 49, -128, -10, -79, 123, -92, 5, -2, 72, 93, -45, -13, -55, 126, 21, -56, 84, 4, -81, -124, -115, 125, 83, -88, 117, 11, 15, -96, -122, -25, 74, -60, 83, 111, 15, -26, 123, -10, 73, -51, 34, -97, -120, 23, 0, 106, 101, 1, -96, -49, -93, -17, -32, -102, -92, -120, 41, 118, -10, -74, -59, -87, -102, 75, 118, -99, 21, -67, 120, 92, -67, -32, -117, 59, -47, -41, 61, 123, -87, 47, -81, -87, 16, -124, 93, -11, -17, -42, -18, 98, 41, 38, 72, -61, 121, 35, -39, 55, -11, 73, 125, 104, 7, 0, 41, 13, 62, 18, 10, 47, 81, 46, -45, -11, -60, -125, 36, 7, -46, 58, -20, 14, -51, 25, 67, -74, -82, 122, 79, -72, -122, -44, -6, -110, 2, -52, 113, -128, -55, 40, -6, -82, 70, -44, 20, -43, -91, 22, -18, -78, 73, 29, 2, 27, -98, 72, -36, -84, 84, 12, -97, -105, 8, -74, -12, 99, -124, 89, -22, 9, -19, 50, -48, 121, 0, 88, 66, -67, 89, 122, -99, -59, 1, 31, -75, -40, -64, 31, -9, 41, 31, -43, -6, 50, -56, 79, 26, 42, -30, 95, -75, 29, -66, -124, -67, -121, 52, -2, -101, -40, 3, -20, -77, 88, 29, 116, -66, -50, 36, -50, -81, -9, 107, 31, 82, 72, -60, 46, -11, -69, 52, 26, 116, -49, -26, -94, 76, -12, -120, 33, 13, -91, 6, -32, 116, -29, -55, 105, -107, 42, -53, 26, -69, -28, -26, -97, 6, -87, 24, -107, -56, -30, -4, -63, 68, 77, 55, 68, -41, -80, 77, 37, -99, 88, 35, -69, 12, -22, 75, 82, -34, 112, 3, -78, 92, 30, 15, -115, 55, 84, 98, 109, 75, 31, 85, -59, -38, -22, 126, -60, -55, 24, -16, -84, 32, -19, 89, 38, -1, 19, -30, -67, -3, -74, 17, 85, 25, 24, -59, -65, -120, 114, -106, -34, -124, -98, 81, -127, -121, 11, -119, 76, -76, -109, 119, -11, -81, 53, 71, -30, 107, 123, 79, -85, 40, 106, 109, -120, -91, -105, 3, 39, 41, 105, -5, -81, -7, 30, -27, 0, 4, -35, -98, -116, 117, -109, -48, 22, -21, -67, 37, -12, 50, -117, 117, 42, -102, -126, -52, -12, -92, 59, -47, 124, 106, 63, -23, -1, 36, 98, -113, 27, -128, -104, 105, 76, -112, 127, 75, 35, 37, -42, -46, -80, 18, -123, 38, 113, -84, -39, -118, 26, 7, 55, 81, -113, 23, -53, -75, -120, 38, 120, 74, 25, -21, -2, 85, -11, 91, -101, 47, 101, -32, 36, 85, -74, 0, 49, 15, 51, -76, -61, -108, 106, 43, 22, -18, -41, 82, -106, -46, 96, 0, 121, -77, 27, 49, -128, 96, -86, 83, 65, 119, -87, -122, -100, -67, 81, -53, -114, 42, -2, 82, -3, 6, -47, 63, 83, 122, -124, -46, -81, -45, 116, -37, -117, -40, -87, -11, 11, -126, -118, -88, -59, 16, 125, 86, -99, -79, 119, -127, -37, 50, 116, -124, -46, -62, -94, -46, 124, 85, 110, 39, 29, -21, -38, 106, 37, -17, -103, 69, -43, -8, -15, 0, -92, -63, 26, -34, 50, -61, -125, -121, -128, 43, 63, -95, -78, -85, 109, 101, -62, -12, -117, -99, 94, -80, -52, 3, 55, 127, -18, 63, -101, 35, 27, 121, 95, 118, -25, -122, -2, -38, 71, 62, -58, -28, -9, 117, 65, 50, 69, 111, -41, 127, -40, -83, -45, -67, 117, 86, -60, -94, 108, 99, 18, -118, 60, 83, 119, 32, 1, -54, -55, 75, 7, -13, -90, -67, -4, 23, 34, -110, 121, -60, 62, 50, -11, 97, 76, -115, -50, 38, 108, -11, -125, -48, 35, 95, 45, -74, 39, 94, 29, -71, -117, -2, -75, 103, -90, -47, -29, -70, -73, -85, -89, -31, -40, 120, -122, -55, -79, 33, -39, 22, 77, 19, -89, 108, 66, -23, -128, -116, -68, -93, 68, 13, 99, 125, 39, -86, -123, 44, -120, 13, 75, 105, -26, 72, -77, -121, 101, -54, 80, 43, 69, 116, 68, -58, -58, -18, -120, 75, -91, -20, 121, -84, 94, 48, 74, 47, 65, -68, 16, -23, 82, 63, 110, -46, -123, -80, -23, 99, -120, 109, -32, 20, 65, -127, 59, 69, -110, -92, -102, -103, 115, -46, -45, -6, -19, 44, -61, 110, 21, -28, -22, -93, 7, -116, -87, -45, -70, -68, -76, -31, 62, 7, 65, 118, 93, -63, -87, 101, -127, 108, -26, -32, 47, 31, -88, -62, 42, 37, 15, -47, 99, -64, 121, 83, -59, -82, -127, -35, 35, -51, 85, -30, 12, 62, 80, 94, -52, 119, -106, -78, 117, -18, 39, 25, -24, -75, -42, 45, -77, 100, -29, 116, 74, 60, 112, 7, -47, 69, -88, -28, -27, -101, -76, 48, 64, 42, -119, -12, -42, -4, 121, 90, 14, 83, -89, -113, -44, -57, 17, 113, -88, 77, 42, -106, -111, -106, 74, -127, 119, 16, -34, 94, -52, 64, 102, 5, -83, -33, 100, -3, -60, -18, 55, -101, -96, -50, -8, -93, 17, -13, -41, 97, -48, 66, -126, 36, 110, 77, 101, 70, 79, -6, -81, -35, 88, 97, -56, 70, -82, 61, 5, -74, 56, 21, -58, -114, -22, 73, 104, -98, 4, -93, -68, 18, 15, -14, 15, -64, -52, 63, 67, -36, 76, 105, 127, -54, -41, 20, -8, -77, -41, -34, 51, -37, 100, 57, 74, 47, -123, -113, -10, -29, 86, -124, -109, 89, -44, -65, 22, -89, -55, -115, -12, -95, -114, -75, -126, -53, -119, -100, -13, 47, -75, -50, 127, 0, 82, -31, 73, -67, -18, -105, -108, -60, -51, 104, 56, -12, -37, 15, -113, -97, -70, -96, -48, -127, -47, -33, 78, 8, -54, -55, -125, -3, 90, -124, -91, 107, -57, -115, -97, 108, 95, 30, -123, -97, 35, -13, 114, -18, 90, -61, -117, -127, -73, 69, 84, 116, 25, 6, 83, -45, 118, 20, -114, 106, 41, -125, -50, 15, -41, -9, -81, 21, -125, 28, -100, -110, 42, 98, -94, 50, 126, -104, -4, 22, 65, -40, -100, -27, -91, 30, -39, -18, 23, -70, -13, -48, 57, 118, -49, 61, 101, 2, -19, 61, 3, 49, -49, -72, 29, -122, -124, -91, -39, 113, 38, 64, -96, 22, 2, 13, 64, 18, -92, -35, -60, -45, -107, -50, -105, 64, -73, 51, 76, -7, 93, -48, -126, -79, 53, -25, 8, -1, 69, 8, -8, -62, 56, -29, -81, -114, -88, 99, 29, -6, 64, -27, -105, -6, -110, -12, 109, 4, -95, 121, -83, 95, -25, 23, -58, 121, 59, -77, 116, 17, 55, -62, -83, -2, -69, -15, 107, 82, -62, -79, 43, -68, 90, -86, 121, -7, 119, 11, -43, -127, 105, -62, 76, 5, -36, -34, -80, -22, 80, 63, -86, -119, 30, -74, 20, -106, -110, 116, 77, 91, -108, 44, -55, 105, 26, 99, -48, -99, 28, 88, 99, 51, 70, -1, -117, 127, -30, 126, 110, -34, -64, 11, 74, -37, 50, -101, 56, -73, 89, 51, -36, -56, 79, 87, -110, 21, 43, -47, -88, -60, 14, 108, -82, -42, -29, -80, 25, 15, 114, -12, 15, -34, 117, 85, -13, -117, -86, -69, -121, -43, -80, 59, 46, -17, -42, 111, 67, -55, -125, -44, 55, 102, 20, -126, -118, -42, -57, -115, 49, 19, -67, 25, 1, 16, 76, -25, -103, -47, -102, -101, -36, -98, -103, 100, 39, -5, -118, 73, -69, -9, 37, 92, 78, 68, -128, 95, -23, -121, -89, 114, 113, 84, 10, 100, 30, 73, -104, -97, 126, -25, -15, 71, -71, -2, 84, 82, 27, -70, -33, 34, -26, -26, 44, 78, -1, 121, 60, 33, 113, 46, -70, -53, 19, 81, 120, 78, -112, 88, -7, 33, -24, -30, 71, 31, -115, 22, -106, -35, -39, -93, -54, 124, 90, -25, -70, -128, -65, 121, -64, -88, -92, -16, 105, 61, 84, -85, 8, -69, -120, -29, 100, -64, 5, -93, 77, -97, -113, -66, -16, 122, -16, 56, -80, 51, 17, -46, -104, 32, 37, -91, 76, -24, -3, 82, 41, 58, -102, 18, -104, -21, -39, -99, -103, -114, 127, 56, -42, -27, -107, -36, 29, 23, 54, -81, 104, 81, -84, -59, -32, -127, -55, -26, 93, 76, -78, -122, 17, -56, 31, 73, -13, -70, -41, -74, -67, 80, 93, -46, 100, -72, 124, 3, -126, 86, -80, -110, 45, 115, 1, -41, 1, 35, 80, -73, -127, -37, -35, 104, -89, 66, 125, 114, -38, 106, -124, -59, -52, -91, -45, 82, 61, 37, -57, 40, 11, -23, -8, -79, 112, -10, -20, -93, -104, 72, 92, 68, 26, -72, 11, 31, -40, -51, 71, -100, -9, -93, 42, -109, -31, -87, -30, 17, -63, 106, -1, -65, 93, 85, -59, -119, -109, -26, 51, -54, 39, -65, -102, 64, 4, 109, -81, 103, 60, -25, -32, 53, -7, -33, -60, -7, -17, 81, 62, -128, 94, -17, 45, 93, -30, -99, 103, 115, -112, 72, 84, -38, -28, 56, 23, -103, 50, -13, -102, 14, 42, 117, 19, 24, -62, -34, -105, -94, -116, -42, -91, 57, 60, 55, -79, -51, 47, -105, -28, -6, -7, -111, -32, 43, -21, 123, 124, -53, -89, 79, 61, 96, 70, -38, -74, -98, 24, -86, -50, -77, -81, 79, 77, -56, 81, -99, -115, 4, -5, 24, 52, 6, -100, 97, -128, -43, -63, 116, 49, 94, -48, -90, 29, -79, -16, 120, 116, 121, 42, 45, -109, -100, 54, 86, 91, -56, 70, 39, -46, -51, 83, -105, -88, 96, -92, -79, -36, 117, -76, -68, 19, -9, -68, 35, 3, 107, 67, -86, -58, -42, -9, -90, 84, -67, -18, -26, 1, 65, 80, -124, 77, -12, 75, -88, -8, -100, 58, -39, -14, -33, 43, -15, -110, 69, 77, 80, 97, 37, 121, -125, 67, -67, -4, 127, -70, -108, 97, 60, -44, 127, 110, 93, 58, 19, -32, 35, 68, 6, -47, -115, 107, 1, -89, -91, 94, -28, -15, 86, -128, 48, 29, -3, -74, -91, -72, -81, -67, -68, -26, 106, -96, 99, -73, -43, 61, 61, -93, 109, -119, -77, 95, -44, -68, -28, 23, 60, -119, -50, 77, -16, 114, 126, 43, -72, 68, -84, 2, -30, 45, -110, -25, 37, 63, 120, 77, 99, 81, 6, -24, -74, -68, -70, 122, 51, 20, -63, -46, -43, 31, -12, -42, -48, 62, 12, -104, 115, -104, 27, 50, 24, 78, -78, -61, 1, -117, -12, -70, -1, -66, -116, -14, 65, -37, -71, -101, 105, 59, -124, 54, -84, 79, -62, 39, 46, 3, -70, 36, -12, 126, 126, 105, 22, -74, 2, 30, 62, -122, 39, -41, -47, 107, 81, -48, -107, -49, -32, -95, 48, 95, -123, -91, 11, -106, -72, 10, 4, 85, -71, 82, -114, 20, 38, -66, 25, -92, 67, 106, -8, -18, -63, 74, -31, 46, -89, 54, -93, -64, -75, 67, -104, -38, 113, 47, -32, 18, 126, -65, -30, -37, 111, -44, -62, -124, -30, 3, 54, -127, 123, -122, -64, 40, -80, 101, 120, 1, 29, 63, -11, 52, 41, 7, 25, 59, 83, -36, 9, 15, -116, -45, -24, 35, 9, -1, -111, 98, 52, 72, -87, 21, -45, -52, 38, -82, 41, -37, -101, 123, 14, 4, 55, 19, -49, -3, 111, 48, -28, 13, 57, -12, -93, -107, 123, -96, 45, -36, 38, 105, 35, 46, -10, 107, 125, 19, 48, -125, -81, -95, -9, -52, 13, 10, 81, 118, -18, 104, -80, -76, -98, -59, 57, -96, 104, 117, -122, -29, -111, 62, 63, -89, -15, -102, 35, 7, 89, -106, 60, 43, 84, 61, 108, -76, 3, 21, -125, 62, 124, -87, 22, -20, -127, -36, -127, -43, 9, -26, 66, 48, 5, -89, -36, 94, 36, 86, -101, 60, 115, 18, 43, -71, -13, 91, 44, -32, 47, 2, -123, -19, 11, -42, -128, -57, -119, -125, 58, 93, 89, 78, -52, 111, -128, -102, 122, 5, -42, 91, 17, -24, 41, 114, 94, -92, -109, 56, 86, -29, -46, 13, 121, 13, 110, -67, 89, 76, 32, -7, 101, -24, 64, 26, -24, 73, -8, 98, 92, -110, -22, -9, -9, -96, 99, -54, 60, -33, 113, -55, -78, 60, 24, 65, 101, -83, -3, -94, -119, 69, -81, -123, 9, 10, 61, 53, -126, -21, -10, 105, -116, 107, -91, -48, 8, 60, -6, -62, 109, 89, -125, 78, 74, 28, -1, 4, -11, 57, -37, -64, -6, -106, 32, -10, -95, -13, 0, -10, 56, 24, -93, -31, 52, 69, 15, 45, 15, 93, -115, 22, 30, 88, 59, -113, 15, -98, 54, 77, -23, 105, -58, -20, -83, -12, -91, 59, 32, 97, 36, -104, -23, -96, 43, -26, 66, -81, 37, -63, -15, 60, -41, 101, -53, -119, -7, 104, 47, 125, -107, -126, 46, -84, -26, -103, 62, -15, 52, 44, -60, -39, 121, -48, 127, -51, 108, 70, 56, 17, 62, 57, 73, 88, -71, -2, -92, 121, -14, 116, -25, -39, 49, 39, -11, 118, 121, 66, -2, -27, 98, -9, -72, 124, 94, -34, 47, 44, 15, -30, -85, 57, 89, 15, -120, -76, -125, 72, 81, -74, 53, -43, 114, -126, 20, 79, -62, -112, 64, -83, 13, 51, 10, -82, 123, -97, -125, -33, 63, -12, 42, 43, 40, -119, 115, 102, 18, 60, 48, -70, 0, -70, -69, -125, 80, 48, 101, 127, -54, 69, -33, 86, -68, -7, 26, -118, -80, -72, -77, 2, 18, -93, -60, -24, -60, 104, 94, 110, 47, -85, 25, -115, -23, 126, -41, -106, -52, 121, 95, 86, -16, 86, -68, 5, -96, 126, -93, 62, -53, -106, -76, -16, 26, -23, -33, -74, 63, 49, 57, 1, 115, -4, -99, 19, 57, 105, -118, -41, -54, -43, -117, 117, -23, 103, -46, -128, -99, -13, -5, -35, 5, 90, 18, 57, 120, -42, -38, 123, -12, 95, -72, 46, -49, 117, -56, -104, 109, 30, 123, -63, 103, -16, 2, -52, 2, -128, -68, -22, -12, -109, 116, -29, -45, 12, 51, 87, 72, 123, 97, -101, -42, 71, 10, -90, 114, 33, 10, -89, 110, 82, -102, -111, -44, -117, -58, 92, -88, -76, 114, 89, -116, -59, 117, -6, 126, -67, 64, 90, -68, -78, 93, 121, -80, -11, 117, 85, -6, 102, -73, 63, -54, 33, 73, 70, -99, -82, 39, 50, -25, -97, 9, 1, -27, 58, -54, -122, -70, -128, -29, 107, -23, 21, 63, 92, -82, 115, 64, -82, 61, -64, -39, 60, 3, 54, -13, 15, 124, 78, 3, -104, 106, -11, 41, -26, -124, 111, 15, -64, -18, -120, 110, 33, -26, -30, 90, 15, 72, 1, -125, -56, -6, -50, -46, -20, -123, 74, 4, 70, 77, 76, 33, -74, -56, -87, -3, -102, 99, -26, 114, 117, -6, -63, -39, 79, 20, 97, -53, -95, 70, -111, 112, -63, 119, 105, -44, -4, -14, -77, 70, 42, -70, 37, -128, 103, 117, 44, -30, -51, -32, 28, 119, 108, -118, -127, 74, -78, 64, -42, -2, 89, -50, 40, -83, -29, 33, -117, -34, 3, 70, 9, 21, -5, -123, 49, 15, 65, 51, 55, 23, -128, 98, -27, -103, -19, 52, -32, -20, -14, -48, -63, -37, -70, 111, -64, 115, -6, 118, -101, -50, 71, 107, -91, -64, -125, 18, -39, 102, -71, -14, -6, -121, 108, -22, -75, 31, -121, 45, 77, -116, 23, -57, 39, 92, -109, 115, -13, 52, -93, 43, -84, -105, 51, -101, 5, 95, -22, 50, -14, -98, -95, 88, -77, 47, 47, -126, 19, 10, -56, 98, -11, -127, -121, 28, -53, 1, 59, -5, 56, 19, 28, -90, 108, -12, 127, -91, 125, -23, 83, 30, -113, -78, -42, -121, -91, -30, -37, -127, 66, 25, -124, -9, 17, -19, 74, 110, -25, 41, 63, -124, -37, -39, -38, 123, -114, 103, 69, 75, 91, -106, -128, -5, -62, 5, -56, -13, 32, -117, -83, -103, -60, -66, -101, -81, 74, 48, 6, -8, 2, 67, -85, -48, -68, 122, -35, 65, 49, 38, 48, -3, -32, -114, -23, 110, 109, -67, -94, 59, 122, 107, 91, -34, -51, 76, -99, 17, 42, 4, -23, -104, 76, 83, -28, -116, 56, 67, -3, 105, -81, 20, 31, 123, 106, -40, -108, 50, -112, 94, -37, -44, 121, 4, -79, 4, 27, 35, 31, 55, 115, 102, -58, 45, 127, 65, 110, 89, 19, 124, 57, -50, -107, 109, 71, -48, 9, 87, -69, -119, -16, -111, -104, 30, -2, -76, -106, 12, -41, 63, -89, -80, 84, -30, 125, -57, 121, 64, -73, 19, -6, 22, 8, -82, -1, -10, 53, -2, 1, -109, -34, -73, 54, -100, 25, 108, 73, -48, 69, 119, 0, 20, -54, -58, 94, -36, -5, -19, -118, 5, 103, -51, 38, -69, -81, 120, -117, 18, 23, 22, 11, -120, -36, -37, 73, -96, 104, -110, 18, 95, -20, -115, 43, 31, 94, -57, 8, -101, -67, 21, 123, -107, -97, -74, -77, 45, 95, 83, 5, 119, -54, -101, -78, -81, 63, 30, 97, 126, 0, 118, 20, -59, -110, -65, -47, 35, -60, -72, -64, 123, -90, -121, -84, -40, -70, 50, -103, 49, 121, 34, 73, 3, 42, -53, -87, -122, 48, -12, -79, -68, -1, -43, -62, -68, 60, -64, -120, -33, -73, 89, -11, 60, -46, 7, -31, -116, -47, 68, 0, 126, -3, -102, -1, -9, -63, 121, -102, -15, 51, 124, 79, 35, -7, -39, 10, -110, -3, 79, 62, -27, 78, 97, 56, -111, 116, 66, -115, 42, 43, 71, -90, -15, -62, 3, -36, -99, 112, 54, -17, -72, -77, -85, 74, -84, 12, 97, 72, -11, 74, 103, -35, -56, 34, -30, -17, 110, 16, 90, -121, -7, -65, 122, -113, 98, -75, -67, -27, 73, -47, -39, -54, -110, -33, -44, 16, -22, 117, 92, -4, 120, -62, 101, -42, -81, -45, 111, 81, -7, -46, -64, -67, 101, -54, 126, 11, -39, -116, 114, 13, 35, -67, -49, -128, 41, -17, 45, 119, -101, -55, 69, 68, -42, 66, 86, -8, -101, 83, 25, 6, 83, 87, -92, 53, -35, -17, -94, 8, -42, 97, -25, -105, -76, -15, 123, 38, -66, -44, -124, 76, -34, 3, -41, 23, -8, 108, -87, -86, 2, 101, 19, 7, -95, 45, -37, -13, -12, -114, -66, 85, -54, 109, 60, 20, 8, -67, 21, 59, -31, -112, 27, -93, -102, -36, 84, 82, 123, -21, 41, -13, -1, -128, 107, -118, -86, 43, 79, 98, 63, 47, -24, -65, -120, 0, -8, 39, -96, -1, -78, 1, -91, -22, 54, -117, -75, -38, -8, 62, -14, -100, -71, 40, -123, 127, 117, -82, -89, 122, 102, 86, -20, -11, 102, 106, -77, 15, 39, -18, 109, -107, 114, -121, 51, 103, -82, -14, -25, -33, 23, 29, 19, -52, -17, -47, -117, -123, 51, -100, -64, 42, 37, -42, 90, -1, -66, -99, 37, -60, 100, -100, 18, 28, -74, -69, 92, -1, 50, -82, 97, 4, 100, -111, -105, 28, 7, -80, 87, 126, 100, 110, -30, 117, -42, 30, 105, -73, 14, -46, -90, 89, -96, 86, -123, -82, 48, -93, 40, 77, -3, -7, -109, 103, 89, -7, 23, -81, -34, -7, 104, -106, -91, -40, -96, -81, 73, -58, -3, 115, -32, -94, -93, 106, 126, -67, -70, 72, -5, -64, -106, 88, -33, 105, -47, 23, 119, 36, -53, -37, 72, -1, -38, 97, 79, 91, -82, -94, -76, 29, -19, 93, 73, -86, 110, 29, -54, 65, 5, 112, -128, -8, -50, 117, -65, 100, -83, 37, 116, 50, -117, 74, -86, 92, -91, -85, -40, 59, -50, -76, -18, 39, -79, -36, 56, -24, 122, 66, -102, 53, 98, -21, -81, -54, -55, -76, 121, -109, 6, -81, -7, -88, 41, 103, 22, 51, -61, 77, 118, -70, 7, -127, 97, -52, 85, 23, 80, -83, 113, -63, -33, -80, -3, -25, -48, 115, -44, -93, 4, 10, 36, 57, 123, -79, 92, -86, 20, 65, 111, 56, -83, 21, -95, 63, -109, -49, 90, 93, -11, 44, 110, -36, -31, 50, -121, 15, -68, 101, 27, 124, -127, -81, 68, 14, 81, -83, 71, -109, 122, -62, -97, 4, 121, 84, 90, 73, -3, 77, -73, -123, 48, -122, 52, 114, -65, -23, 13, 98, -8, -111, -38, 58, -13, -90, 69, -121, 90, 82, 114, 39, -12, -51, 85, 86, -14, -28, 94, 65, 81, 72, -95, 66, -64, 33, -89, -77, -21, -78, 121, -91, -104, -43, -119, -13, -78, -78, -34, 59, 98, 115, 3, -4, 82, 7, 37, 66, -53, -110, -103, -112, -24, 14, -40, -25, -108, 56, -100, 22, -108, 52, -113, 126, -6, 122, 4, 0, -73, 111, -90, 18, -76, 73, 38, -58, -50, -40, 46, 110, 61, -59, 97, -22, -50, 35, 42, -61, -40, -29, -60, 50, 127, 88, 47, -51, 22, -108, -22, 53, -123, 101, 89, -95, -12, -86, -87, -53, 116, 3, 120, -50, -104, -19, 27, -126, 30, 21, -42, 52, 59, -127, -109, -9, -91, -77, -82, 124, 79, 48, -53, -22, -114, -127, -4, 86, -111, -59, 53, 48, -57, 78, 110, -40, 119, 105, -77, -70, 23, -95, -70, 32, -18, 8, -48, -63, 22, 88, 1, -18, -113, 55, -58, 24, -94, 6, -90, -18, 73, 75, 49, -120, -14, 114, 73, -3, -2, -109, -53, -51, 72, 41, -120, 88, -52, -43, 0, -108, -11, -28, 94, -115, 93, -7, -18, -75, 108, -8, 83, -28, 117, 55, 46, 40, 111, 64, -30, -68, -40, 37, -127, -110, 67, 38, 15, 95, 9, -74, 122, -72, 45, 22, 82, -110, -76, 9, 106, 69, 93, 7, 85, -81, -26, -112, -125, 50, -106, -88, -27, 58, 98, 15, -44, 8, -101, -2, -55, 56, -51, 44, -115, 111, 9, 34, -121, 23, 59, 38, 95, -49, -13, 98, -127, 27, 125, 79, 34, 9, 108, 75, -30, -106, -87, 25, -63, 5, 9, 63, 91, -17, -128, 83, -40, -114, 113, -72, 100, 79, 118, 68, -33, -38, 15, -101, 72, -46, -120, -62, -14, 25, -62, -105, 69, -48, 41, -25, -5, -60, -120, -3, 72, 0, 39, 54, -101, -28, -13, -13, 21, 16, -26, -77, -80, -14, 15, 37, 48, -63, -80, 33, -35, -53, 89, -127, -117, -26, -96, 48, -22, 80, 110, 46, 93, 6, 0, -105, 35, -119, -85, 4, -53, -128, -45, 1, 19, 45, 26, 94, 51, -35, -50, 6, -24, 99, 118, -71, -102, -68, 89, -6, -119, 122, 65, 46, 23, 24, -126, 49, 35, -34, 71, -117, -30, -22, -27, -18, 22, 28, 44, -15, 25, 57, -121, 109, 78, 27, -126, -115, -63, -48, 47, -78, -112, -46, -44, -82, -110, 81, 55, -40, -14, 5, -96, -86, 87, 2, 82, 83, 50, 89, -4, -25, -110, -8, -99, -106, -16, 32, 16, -102, 101, -70, 96, 40, -105, 90, -98, 7, 6, 67, 74, 28, 19, 99, -32, 32, 54, 8, -81, 46, 103, 24, 88, -112, 55, 110, 8, -12, 122, -82, -92, -68, -96, 109, -64, 49, 69, 75, 117, -75, 92, 68, -47, 33, 20, 19, -89, -18, 110, 43, 67, -91, -26, 9, -103, -92, 77, 22, 126, 0, 37, 31, 116, 6, 29, -90, -65, 103, 33, -60, -67, 38, 19, -43, -35, 91, 48, 70, -114, -22, -35, 6, -122, -65, -15, -111, -26, -27, 1, -118, -82, 108, 89, -84, -41, 122, 48, -30, -18, -110, 12, 34, 27, -24, 87, -78, -112, -78, -128, -53, 74, -127, 101, -12, 60, 3, 56, 127, -39, 96, -16, -74, 110, 44, -96, -51, -11, -39, -113, 98, -37, 97, 36, -119, -80, -88, 31, -4, 11, -19, 59, -84, -121, -70, -79, 97, -25, 22, -8, -79, -60, 39, -108, -79, -72, 46, 124, -9, -18, 121, -93, -128, 95, -98, -24, -17, -79, 62, 95, 64, -55, 85, 70, 116, 41, -8, 35, 18, 82, 15, -13, -106, -92, 96, 84, -17, 102, 75, -33, 6, 74, -108, 56, -46, -77, 60, -47, -31, 112, -23, -64, 27, -15, -126, -94, -72, -86, -48, -73, -49, 99, -23, 66, -108, 109, 8, -28, -105, 73, -7, 109, 85, 31, 66, -128, -4, 42, -61, -18, -61, -122, -4, 69, -80, -119, 93, -89, 119, -128, 113, -76, -98, 99, -115, -55, 105, 72, 25, -87, 40, -98, 79, -117, -87, 32, -77, -45, -37, 73, -105, 74, 113, -6, 38, -113, 66, -25, 45, 19, -77, 51, -29, -15, -79, 42, 50, 43, -25, 94, -92, -116, -28, 78, -96, -17, 42, -81, 68, -124, -43, 91, -25, 115, 5, 33, 40, 59, -33, -69, 18, 57, -39, 117, -45, -18, -90, -108, -67, 11, -116, 112, -99, -77, -67, -55, -127, -109, 48, 76, 15, -85, 65, -29, 79, -102, -74, -12, -42, 18, -73, -66, -122, -40, 61, -59, 63, 46, 121, 27, 104, 23, -3, 87, 112, 78, 87, -66, -26, -61, -42, 24, -52, 40, 90, -5, 18, -34, -47, 25, 9, 7, -79, 116, 102, 110, 95, 0, -68, -1, 56, 61, 11, -127, 60, 107, 117, 89, 10, -49, -115, 89, 62, -32, -14, -10, -110, -59, -51, -113, 75, -120, 48, -17, -97, -58, 106, -81, 22, -27, -46, -121, -75, 88, 29, -103, -3, 73, -38, 22, 96, -79, -47, 84, 72, -77, -73, -41, -75, -50, 81, -106, 79, 70, -45, 97, -121, 62, 70, 9, 71, 8, -116, -29, 67, -90, 69, -89, -16, 84, -12, -38, 64, 95, -34, 98, -45, 109, -52, 70, 28, -1, 25, -46, 120, -86, 86, 4, -21, 29, -42, 20, -42, 22, 11, 49, 76, 24, 113, -71, 35, -117, 7, 50, 64, 9, 105, -77, 108, 87, 93, 59, -124, 45, -82, -49, -38, 79, -88, -5, -41, 108, -15, 42, 29, -126, -97, 4, 42, 45, -106, 114, -50, -112, 122, 22, 31, -9, -56, -103, -98, 116, -127, 17, -14, 70, -10, 22, 123, 78, 114, -43, -10, 7, 57, -108, -5, 28, 118, -6, -12, 52, 25, -115, -112, 78, -109, 104, -24, -15, 29, 55, 6, 120, -2, -63, -74, -91, 115, 124, -127, -29, -119, -32, -23, 66, -11, -125, 104, -60, 106, 17, -69, -45, -67, -39, -8, 99, -10, 40, 72, -122, 126, 103, 10, 93, -30, -49, -105, -67, -41, 71, -43, -9, -124, -89, -66, -55, 11, 45, 79, 68, 48, -128, 40, 39, 3, 62, 40, 77, 51, 73, -90, -89, -23, -48, -37, -64, 56, -83, 119, 29, 57, 86, -111, 65, -21, -117, 59, 53, 22, -72, 117, -65, -22, 67, -86, -26, -93, -50, 103, -87, -65, 69, 80, -85, -67, -40, 106, 95, 10, 55, -98, 83, -35, 124, 110, -60, 61, -16, -92, 101, 29, 103, -106, 116, 114, 98, -23, -99, -19, -54, 60, -112, -56, 42, 87, 88, 123, -93, 0, -87, 15, -45, 81, -21, 51, 113, -91, -93, 107, 13, -1, -86, 62, 23, -8, 4, -58, 94, -65, 90, -37, -23, 109, -71, 124, -109, 99, -76, -45, -14, -76, 82, 42, -91, 62, 89, -80, -118, -105, 75, -77, 115, -54, -102, -101, -60, -18, -18, 33, -19, -19, -22, -12, 104, 97, 31, 46, 91, -128, -6, -41, -108, 80, -96, 57, -117, -36, 31, -109, 41, -123, 106, 5, -58, -88, -14, -102, -44, 60, 52, -22, -8, -116, -29, 38, -106, -22, -118, 83, 7, -23, 86, -69, -25, -76, -84, 41, 82, -20, 6, 124, 5, -113, -59, -56, -103, 30, -84, -60, 47, -109, -83, 0, -128, 58, 4, -41, -126, 18, -87, -78, 91, 57, -23, -81, -56, -83, 29, -19, 106, 75, 33, 75, 117, -49, -98, 41, 4, 8, 48, -61, -21, 92, 73, -51, -53, 23, 123, -25, 45, 59, 49, 40, -37, -56, -3, 122, 73, -123, -108, 127, 115, -46, 3, -104, 126, 72, -38, 69, 18, -99, -70, 59, 110, 2, -127, 3, 6, -102, -41, -43, 90, 47, -102, 3, -84, 27, -87, -121, 80, -43, -74, -26, -93, -70, -23, 39, 14, -23, -94, -78, 5, -32, -1, 73, -105, 90, 88, -47, -6, -83, 68, 36, 6, 72, -74, -106, -103, 27, 40, -3, -127, 92, -53, 107, -20, -127, -78, 83, 14, 62, 41, -117, 28, 61, 74, 105, -56, 88, 2, -65, 98, -33, -47, -66, 111, -100, -98, -119, -68, -103, -62, -17, 63, -103, -89, 1, 113, 49, 24, 27, -11, -18, 61, -111, -80, -10, 6, -85, -15, -74, -17, -26, -123, 104, -88, 49, 116, -110, -50, -93, 30, -27, -41, -81, 101, -88, -4, 32, -36, 50, -106, -3, 51, 5, 89, 31, -121, 44, -67, -84, -6, -25, 18, 55, -76, 98, -77, -81, 61, 67, -66, 85, 90, 105, -12, 126, -29, 45, 1, 18, -118, 103, 120, 50, -123, -105, 7, -70, 38, 46, 32, -123, 127, 65, 65, 13, 4, -27, -96, 32, 79, 4, -94, 78, 83, 36, -101, 5, 119, -86, 111, -96, -118, -3, -94, 38, 88, -47, 26, 56, 9, -98, 40, 86, 3, 96, -117, -25, -121, -1, -65, -55, -105, 78, 89, -2, 111, -29, 115, -103, -31, 1, -99, -116, 64, 121, -7, 107, 17, 96, -63, 18, -117, 55, -83, 52, -8, -10, 15, 25, 50, 17, 79, -87, 18, 60, 70, -119, -59, 33, 14, 55, 15, 99, 48, 28, 39, -105, 68, 22, -4, -63, 62, -45, 108, 112, -55, -95, 17, -14, -79, -117, -121, -3, -66, 124, 89, 18, -80, -102, -103, 105, 105, -82, -38, 34, -104, -73, -90, -123, 51, 75, -34, -114, 116, -81, -119, -5, 81, -9, 38, -111, 54, 71, -79, 66, 33, 30, -102, 71, -119, 62, -106, -105, 85, 60, -78, -83, 82, -115, 46, 87, 105, -79, 99, 24, -69, 41, -19, 107, 71, -109, -85, 29, -5, -26, -87, 13, 31, -37, -96, 37, 7, 2, 43, -11, 2, 112, 28, -51, 61, 56, 0, 10, 13, -70, -85, -88, -21, 58, 70, -111, 71, 106, -112, -50, -90, 15, 91, -93, 70, -14, 11, -20, 45, 15, 29, 47, 127, 47, -41, -85, 58, -49, -104, -22, 77, -93, -76, 122, -101, 58, -2, 73, -116, -124, -8, -69, 108, 35, 115, 73, -91, -18, -13, 1, 8, 71, -94, -113, -92, -102, 30, 64, -89, -40, 65, -60, -77, -101, -38, -94, 85, 77, 83, 14, -98, -16, -5, -111, 117, 71, -102, 66, 102, 48, 21, -32, -36, 98, -104, 22, 21, -33, 8, 44, 46, 98, 58, 48, 38, 119, 92, -23, 66, -21, 28, -12, 71, -19, -66, 36, -40, 15, -71, -35, -110, -89, 31, 74, -52, 41, -28, 31, 107, -115, 88, -46, -70, 79, 90, -58, 32, 76, 67, 87, 112, 69, -35, 98, -116, -45, -15, -2, 66, -119, -80, -53, 10, 87, 116, -73, -53, -91, 84, 11, -115, 57, -29, 71, 56, -52, 120, 65, -34, -45, 0, -21, 0, 97, 41, -89, -18, 10, -86, 119, -11, -103, -37, -97, 113, -58, -84, -56, -113, -21, 72, 56, 63, 8, 14, 57, -9, -39, 6, 50, 95, 44, 26, -103, -86, -28, -84, -127, 32, -74, 22, 67, 95, 54, 116, -80, 120, 114, -3, 86, -34, -91, -102, 113, 64, -97, 111, -5, 17, 101, 48, 117, -6, -2, 109, -105, 12, -75, 9, -123, 72, -17, 105, -110, 57, 68, 70, -61, -38, 40, -123, -97, 36, 87, -31, 68, 120, 21, 71, 26, -59, -55, 14, 118, -21, 119, -68, 68, -39, -11, -96, -62, 89, 45, -55, -80, -126, -104, -112, -9, 52, -127, -112, -118, 19, -18, -75, 93, 107, -50, -47, -72, 40, -66, 62, 126, 47, 45, -121, 121, -37, -3, 69, -81, 63, -14, -65, -124, 83, 108, 52, 116, 115, 67, 16, -81, -41, -11, 9, 80, 111, 64, -61, 3, 20, 90, -43, -90, -33, -11, -68, 107, -25, 56, -3, -4, 100, 27, -59, 23, 13, -115, -28, -14, -55, 109, -39, 22, 54, -17, -25, 45, -15, -95, 104, 109, 126, 33, 125, -101, 101, 42, 70, 80, 24, -99, 127, 110, 45, -37, 20, -65, 65, -67, 107, 35, 75, -56, 36, 122, 25, -75, 22, -16, -95, 7, 111, 40, 41, -8, -54, 16, -82, 1, 127, -96, 69, 17, 60, 63, 101, -83, 34, -21, -118, 100, -94, 95, -21, 106, -54, 72, 55, -24, 47, 79, 116, -41, -122, 5, 7, -109, 46, 15, 118, 22, -15, -55, -9, -42, -25, -3, 8, -126, 68, -57, 125, 84, 49, 0, -5, -98, -117, 107, -11, -86, 120, 73, 74, 0, -49, -104, -37, -28, -105, 26, -107, 60, -103, 96, 126, -45, -80, 105, 19, 113, 114, 99, -22, -109, 111, 7, -39, -80, 10, -72, 86, -17, 6, -1, -107, -99, -65, -15, -51, -112, 120, 119, 121, -93, -88, -20, -112, -103, 15, 116, -122, -46, 20, 25, -107, 99, -121, 33, 38, 48, 114, 56, 44, 67, 29, -30, 110, -41, -97, 103, 29, -45, 50, 112, -70, -115, -117, -47, 39, 40, 3, -33, -8, -103, -87, 68, 9, -5, -2, 26, -49, 23, 71, 89, -49, -102, 84, 71, 26, -96, -80, 39, 35, 70, 56, -49, -21, 50, 3, 81, 61, 98, 15, -71, -70, 12, -31, 68, -76, -107, -115, -72, 28, 7, 97, -3, -17, 124, 27, -39, -87, -44, -88, 63, 119, 38, -10, 94, -75, -51, 113, -126, -54, -7, -71, -30, 105, 24, -37, 51, 7, 102, -98, -114, -125, 41, -81, 65, 117, 92, -101, 123, -19, -41, -108, 81, 105, -123, -70, -7, -3, -109, 114, -47, -100, 46, -48, -122, -14, 54, 98, 67, -79, 95, -3, 17, 90, 56, 70, -18, 79, -75, 23, -87, -95, 24, 37, -105, -87, -85, -120, -67, 4, 81, 16, 25, -3, -3, 123, 110, 47, -10, 47, 24, 8, -10, -49, 61, -122, -103, 69, -11, -58, -8, 97, -77, -35, 69, -66, 121, 118, -63, 97, -41, 51, 120, 22, -38, -126, 69, 88, 1, 68, -76, -102, 74, -30, -6, -48, -92, 59, -118, -14, -31, 27, 104, 119, 94, -81, -78, 1, -81, -50, -117, -39, -25, -76, 54, -40, -14, 57, -120, -86, -12, -108, 61, -59, 127, 92, -34, 83, -102, -122, 26, 111, -85, 6, -61, -116, -32, -56, -127, 96, 43, 63, -102, -18, -45, 110, -85, 25, 86, -109, 4, 46, -70, -100, -96, 5, 38, -63, 90, -126, 66, 89, -10, 78, 72, 124, 40, -112, -97, -110, 0, 126, -110, -7, 36, 31, -58, 80, 75, 53, 39, -9, -34, -2, 79, 84, -28, -23, -90, -76, -44, 25, -93, -38, -27, 55, 78, 87, -45, 113, -52, -123, 44, -66, 46, 80, -38, -108, -21, 52, -7, 25, 108, -92, -60, -71, 94, 44, 113, -89, -47, 30, 42, -100, -79, -119, -38, -14, -121, -100, -59, -79, 71, -127, -116, 121, 13, 12, 87, -6, 82, 63, 56, 49, 84, -84, -45, 15, -65, 73, -35, -125, 103, 76, -53, 57, 82, -109, -2, 5, 45, -16, 109, 52, 98, -76, 18, -32, -80, 24, 48, -74, -53, -65, 75, -2, 31, 21, -61, -90, 48, 6, 126, 51, 80, 22, 111, -89, -116, -35, 60, -20, -47, 33, 0, -127, -73, 63, 2, 60, 57, -2, 104, 107, 53, -26, 81, 20, 110, -108, -107, 64, 35, -84, 14, 101, -59, -113, -47, 57, -35, -7, -61, 47, -62, -15, 61, 78, 23, -95, 0, 27, -78, -5, -46, 36, -32, -12, -116, 3, 54, 46, 93, -6, -6, 13, -73, 50, -102, -37, -76, -96, 0, -13, -125, 44, 76, 91, -7, -93, 70, 72, -60, 95, 112, 86, 2, 86, -72, 8, -7, -91, 88, 34, -16, -105, -119, 78, 28, -25, -34, -20, 63, 63, -125, 84, 87, 124, -58, 118, 114, 64, 62, 34, -94, 118, 22, -80, -108, -103, -85, 39, -61, 124, -36, -116, -112, 32, 47, 96, -116, 76, 19, -23, -65, -112, 78, -14, 36, -118, 91, -12, -1, 71, 6, 6, 37, -20, 29, -108, -101, 84, -94, -40, 16, 16, -113, 62, -32, -12, -42, 25, -72, 62, 124, 85, 101, 62, -111, 67, 62, -70, -113, -106, -9, 86, -15, 1, -56, -33, 74, 95, 55, 25, -83, -92, -20, 66, 69, -60, -59, -48, 20, 26, 43, 49, 62, 42, -69, 78, 111, 81, 127, -4, -97, -77, -124, -65, -60, -125, -28, -127, -70, -53, 60, -97, -11, 71, 34, -45, -128, -1, 123, 20, -73, 71, -4, 35, -10, -25, 49, 98, -19, -85, -123, 42, -90, 57, 56, 114, 64, 106, 34, 110, 44, 29, -109, 62, 97, -68, 72, 106, 53, -50, -14, 116, 109, -85, -30, -106, 51, 127, 35, 62, -81, 108, -61, -99, -84, 118, -114, -35, -93, 14, 123, -94, -15, 4, 56, 17, -127, 103, -123, -111, 13, 60, -41, -79, -65, 95, 89, -73, 116, -18, -125, 70, -91, 102, 47, 86, 59, 21, 106, -84, -37, -25, -64, -115, -92, -21, 37, -14, -123, 19, -86, 111, -75, 27, 113, 19, -7, -7, -68, 48, -97, 78, -103, 25, 23, -84, -52, 5, 12, -94, -76, 14, 40, 65, 76, 16, 123, 118, -54, -31, -110, -49, -82, 107, 18, -46, 4, 107, -4, -123, 13, 101, 91, 102, 42, 100, 20, 108, -21, -13, -4, -114, -16, 57, 123, 42, 114, 31, -82, -119, -73, 78, 15, -17, -84, -91, 50, -6, 89, 76, -53, -42, 101, 74, -89, -29, 52, -128, -32, 39, 21, -46, 58, 79, 71, -99, -126, 55, 113, -113, 37, 52, -81, -18, -124, 50, -24, -24, -36, 101, 59, -7, 2, 28, -83, -81, -127, 57, -102, -107, -44, 17, -43, 111, 113, -102, -108, -62, -53, -59, -37, -128, 41, 105, -15, 111, 73, -13, 85, -6, 62, -107, 0, -119, -35, -39, 18, -21, 105, 113, -110, 111, 4, -92, -53, 9, 48, 120, 44, 72, 75, 123, -42, 9, 86, 122, 42, -80, 55, 75, -40, -125, 3, 31, -109, -37, -47, -91, -17, 21, 117, 71, 67, -113, -84, -27, 11, -21, 32, -51, -29, -101, 82, 30, -84, 13, 123, -97, 46, 0, 53, 46, 9, -42, 34, -128, -100, 7, -19, 95, -27, -79, -21, 71, 10, 3, -70, -92, 43, 109, 76, -38, -69, -28, 68, -16, 55, -126, -35, 116, 120, 59, -19, 108, 72, 67, -56, -91, -43, 81, 101, -30, 69, -49, 88, -87, 82, -55, -111, -124, -71, 45, -38, 31, 62, -95, 25, -99, 62, 19, -99, 81, -30, 115, 118, 52, 102, -89, -39, -30, 17, -83, -94, -11, -33, 69, -16, -128, -3, -126, -65, 33, 115, -25, -52, -41, 112, -122, 48, -28, -8, 108, -37, 44, 71, 58, 99, 112, 55, -17, 104, -68, 37, 13, -3, -16, 113, -128, -64, -1, -112, 80, 51, 50, 10, -62, 11, -113, -94, -67, 33, -121, -93, -6, -80, -12, -90, 76, -81, -13, 13, 19, -52, -96, 71, 96, -29, -63, 43, 116, -33, 12, -73, 63, 29, -119, 57, 46, 126, 117, -45, 58, -89, 52, 86, 105, -40, -36, 67, 50, -82, -14, 75, 102, -93, -30, -53, -120, 83, -59, 99, 89, -105, 102, -3, -65, 27, 66, -1, -103, -115, -37, -100, 97, 108, -82, -5, -10, 38, -64, 77, -124, 110, -54, -27, -16, -68, -115, -95, 19, -65, -27, 73, -22, -109, 46, 76, -35, 101, 125, 104, -32, 21, 79, -59, 71, 42, -79, 115, -46, 4, 6, 95, -125, 102, 121, -55, 30, -36, 71, -123, -125, -126, 47, 112, 31, -80, -124, -13, 126, 6, 117, 39, -6, 2, 98, 68, -20, -64, 32, -17, -62, 31, 110, -103, 98, 92, -69, 78, -7, -94, -7, 41, -4, -23, 83, -84, 124, 99, -115, 16, 16, -79, -65, 12, 69, 71, -60, -78, 105, -66, 43, -114, 53, -73, 99, -20, 22, 125, -107, 47, -111, 126, 25, 55, 121, 120, 120, -52, 87, -119, -22, -66, 112, 68, 96, -109, -118, -44, 125, -72, 69, -57, -91, 34, -60, -117, 36, 127, 68, -84, 43, 18, -27, 35, -116, -12, -94, 9, -78, 83, 127, -43, 109, 7, 61, -98, 8, 25, -39, -4, -91, -1, 45, -42, -87, 24, -58, 107, -103, 79, -40, 115, 51, 53, 92, 18, -66, -112, -14, 109, 100, 60, -35, -91, 41, -63, -28, -53, -100, -106, 70, 107, -78, 88, -97, -57, -96, 127, -25, -127, -50, -119, -101, 69, 101, 28, 94, -30, -47, -125, -38, 12, 9, 83, -108, 17, 107, -109, -46, 15, -19, -13, 105, 108, -97, -88, 34, -117, -96, -90, -103, 123, -59, 84, -74, -87, -17, -8, 11, 36, 107, -24, 38, 24, 73, -57, 81, -28, 75, 59, -87, -119, -58, 110, 125, -29, 110, -66, 108, -90, -31, 41, 118, -44, -67, -127, 67, -11, 83, -48, -127, -116, 10, -33, -85, 85, -46, 26, -54, -37, 112, -26, -117, 79, 25, 1, -27, 96, -100, 49, 126, 111, -37, 14, 58, -124, 78, -33, 7, 34, -110, 71, 30, 91, 104, -118, -12, 112, 117, -102, -5, 105, -45, -31, 26, 13, -115, -18, 46, 45, -69, 69, -66, 66, 62, 88, 67, -107, 64, -126, 29, 76, 17, 107, 23, -120, 82, -122, -3, -62, -56, -75, -24, -119, -119, 54, -12, -109, 82, 25, -101, -106, -86, -83, 33, 62, -39, -122, -68, 53, 19, -118, 118, 69, 94, -78, -27, -54, 65, -127, 55, 52, -36, 9, -38, 72, 119, 35, 47, -94, 6, 38, 78, -45, -51, 7, -49, -99, -99, 71, -19, -10, -81, 5, 34, 37, -26, 23, -55, -14, -21, -66, -113, -50, -19, 111, 92, -15, 122, 82, 0, 106, 124, 107, 84, -8, 61, -77, 62, 110, 38, 112, 30, -73, 114, 58, -18, -35, -38, -117, -97, 111, 33, 50, 53, -40, 9, 14, 9, 37, 82, -20, 9, 76, 86, -59, 72, -58, -109, -57, -19, -27, 33, -7, 47, -54, -45, 29, -95, -38, -58, -51, -43, -58, 94, 74, -7, 75, -39, -43, -37, -67, 45, 14, -26, 44, -38, -115, 80, 84, -109, 10, -32, -19, 56, 43, -49, -35, -38, 58, -11, 87, 74, -87, -111, 117, 77, -8, 105, -5, 73, 108, -67, -75, 117, -44, 36, 43, -92, -72, -84, 73, -118, 120, -104, 90, -23, -89, 78, 91, 30, -14, 74, -93, 73, -5, -5, 48, -29, -31, -122, -49, -52, 91, -126, -114, 111, 44, 120, 56, -116, -123, 83, -86, -40, -42, 33, 124, -44, 40, -126, 46, -54, 5, 86, -49, -105, -4, -64, -23, -13, -19, -72, 35, -35, -93, 57, -58, 40, 112, 72, -100, -120, -2, -63, -15, 124, 6, -7, 20, -44, -1, -19, -31, -55, 73, -4, 53, 91, -8, 17, -28, -121, -96, 36, -7, 39, -69, -87, 48, 55, 21, 104, 63, -94, -126, 32, -114, 18, 126, -112, 32, 91, -15, 36, -92, -80, -97, -125, -12, -125, -31, 25, -48, 117, -29, -109, -67, -46, 113, -36, -61, -120, -53, 113, 72, 81, 8, -49, -121, 106, 26, -19, -94, 29, 122, -6, 103, 44, -18, 20, 57, 13, -99, 67, -113, -107, -94, 80, 22, -112, -23, 23, 38, 34, 47, -36, 23, -96, -109, -1, -68, 116, -110, -9, -24, -25, 41, -81, -109, -29, 81, -13, 118, -36, -35, -122, -97, -14, 87, -106, -46, -55, -69, 76, 35, 34, -98, 30, 45, 64, 30, 108, 83, 88, -36, -78, -26, 118, 15, -60, -109, 80, -115, 87, 94, -113, 100, -71, 121, 55, -90, -115, 49, 2, 7, 33, -7, -9, -25, -6, -16, -23, 113, -100, 4, 55, 103, -92, -119, 6, 50, -75, 127, 103, 51, 73, -101, -57, -9, 91, 102, 60, 77, 57, 103, -113, 18, 38, -73, 125, 40, -14, -106, -116, -115, 116, -60, -128, -101, -97, 85, -116, -22, -69, 62, -44, 73, 109, 127, -83, 102, -128, 121, 38, -118, 98, 26, 40, -46, -58, 102, -10, -51, 1, -128, -115, -77, -4, -9, 88, -127, 36, 46, 49, -31, 87, -17, 41, 9, -103, 97, 91, -59, 91, 65, 68, -72, -41, -47, 117, -58, 7, 52, -3, 126, -69, -98, -121, 17, -119, 120, 99, 43, -124, 94, 74, -88, -94, 112, -1, 127, 15, 109, 43, -78, 45, -13, -80, -16, -76, 70, -9, -121, -64, -35, 125, -51, 17, 59, 111, -42, -55, 112, -84, 74, -101, -20, 108, 35, 59, 4, 41, 44, 117, 68, 32, 126, -3, -92, 13, -77, 65, 106, 122, -114, -11, -16, 84, -80, 85, -83, 17, 68, 31, -31, -104, 29, 4, -88, 30, -38, 64, -16, -106, 105, 27, -109, -42, 7, -80, 89, -74, 111, 93, 18, 68, -30, 104, 53, -32, 11, -5, 6, -17, -121, -19, -35, -43, -104, 18, 121, -102, -65, 92, 36, -126, -105, -78, 27, -18, 34, 102, 26, 60, -43, -72, -47, -99, 63, -86, 25, 38, 115, 40, -23, -45, -43, -19, -4, -88, -106, 31, -80, -61, -41, -38, -66, 74, -19, 65, 75, -20, -64, 11, 56, -14, 42, 2, -39, -63, 27, 86, 28, -100, -43, 70, -1, -118, 40, -53, -2, 40, -58, -13, 16, 106, 100, 116, 64, -18, 113, 124, -65, -38, 2, -107, 31, 41, -47, 110, -76, 50, 64, -114, 105, -58, 74, 73, -70, 103, 30, 25, 39, 11, -13, -113, -75, -71, -40, 66, -106, -41, -126, -122, 44, -47, 16, -70, -2, -10, 13, 19, 106, 97, -63, -67, 40, -61, -98, 56, -67, 73, 108, 107, 98, -3, 100, 6, 11, -66, 78, 5, -80, 46, -18, -2, -29, 115, 109, -90, -40, -26, 55, 29, 110, 60, -115, 59, -116, -68, 102, 115, 115, 73, -36, 81, 84, 28, -108, -5, 33, 75, -7, 86, 112, -70, 1, 34, 31, -28, 108, 65, 21, -43, -20, 93, 118, 61, -20, 99, -99, -113, -116, -122, -13, -64, 83, 99, 14, -104, -57, -58, -17, 22, 70, 36, -127, -55, 78, -32, -72, 126, -54, 30, 80, 30, 69, -122, 86, 76, 107, -12, -110, -102, 105, -19, -124, 72, -36, -34, -12, -3, -71, 38, 52, -126, 110, -20, -79, 126, 95, -86, 3, -12, -45, 62, 95, 60, 28, 65, 75, -112, 33, 117, -20, -103, 86, -76, 29, 39, -113, 54, -74, 4, -112, -100, 81, 77, 90, 40, -96, -22, -19, -60, 124, 119, -93, -65, 92, 43, 77, -106, 83, -68, 119, 58, -30, -40, 44, -120, -64, 55, 80, -26, 12, 71, 80, 85, -34, -116, -45, -122, 70, -76, -57, 78, -111, 99, 119, -1, -57, -41, 32, -90, 123, -73, -97, -99, 118, 17, 87, -42, 97, -23, 10, -110, 84, 60, 54, 72, 60, 119, -26, 27, -27, 51, 39, -99, 8, 28, 80, -98, 116, 67, 0, 11, -53, 11, -41, -95, 69, 71, 118, -74, 76, 101, -30, -95, 108, -6, -93, 117, -128, -107, 52, 51, -23, -102, 50, 70, -51, -120, -37, 117, 64, -122, 124, 115, -72, 23, 120, -60, 23, 111, -55, 28, 32, 78, 74, -20, 44, -48, 10, 70, 86, 48, -125, 15, -34, -58, 5, -104, -14, -103, 86, 119, 26, -106, -61, -2, 108, -48, -57, 109, -128, 39, 75, -32, 82, -104, 17, -55, 8, -1, -77, -51, 60, -38, 110, 38, -117, 117, 83, -36, -88, 13, -70, 27, -14, -14, -47, -107, 126, 65, 47, -119, 120, -93, -44, 96, 2, -49, 67, 93, 74, -50, -61, 40, 51, -21, 71, -48, -41, -97, -84, -108, 71, 81, 92, 50, -33, -102, 14, 27, 63, 29, -88, 76, -33, -93, 112, -67, -3, -6, 56, 104, 25, 57, 81, -125, 35, -57, -89, -118, 10, 42, 82, -127, 30, -120, 29, -25, 95, -4, 18, -72, -95, -71, -89, -22, -72, 115, 23, -125, 61, -46, -88, -39, 119, -119, 5, 39, -91, 110, -37, 13, 69, 1, -127, 71, -106, -101, -17, 62, 46, -39, 30, -83, 92, -51, 92, 117, -63, 25, 58, -16, -39, 54, 88, -52, 75, 49, 42, -121, 46, -17, -53, -59, 41, -20, -47, 100, 40, -95, -33, 79, -106, 34, -37, 100, -16, 122, 73, 110, 2, 42, 56, 11, -15, 119, -4, -14, -37, -13, 38, 11, 25, -15, 116, 95, -90, -30, 125, -94, -90, -41, -89, -52, -38, -93, 18, 6, 99, 44, -69, -86, 61, 104, 48, 91, 120, -6, -56, -71, -39, -20, -84, -17, 124, -14, -99, -84, 92, -42, 12, -38, 116, -42, 34, -21, 47, 78, -18, -41, -113, 66, -22, -15, 119, 14, 95, 38, 4, -2, 59, 97, 13, 110, -32, -101, 92, 97, -48, -71, -81, -40, -32, -89, -27, 77, 64, 104, -18, -3, -58, -2, 115, -30, 86, -69, -50, -68, -22, -60, 90, 88, 14, 116, -43, 122, -67, 103, -30, 55, 47, 33, -90, 65, -51, -108, -1, -124, -34, 2, -54, -81, -125, 34, 125, 15, 74, -66, -12, -103, 114, 98, -26, 92, 42, 89, -66, 114, 125, 84, 124, -120, 93, 106, 84, -115, 117, 33, 102, 9, 74, 60, 5, -47, -57, 84, 123, -21, -107, -90, -58, -77, -60, -70, -62, 82, -21, 105, 107, 104, -74, -35, -53, 123, -105, -68, 5, 4, -23, 86, -121, -10, -12, 37, -59, -71, -100, -105, -48, 16, -124, -108, 50, -125, 68, 50, 71, -48, -72, -118, -96, -98, 117, 127, 99, -117, -124, -60, -15, 43, -43, -14, 77, 9, 50, 113, 75, 114, 11, -53, -7, -20, -14, 111, 116, 4, -102, -116, 67, -57, -103, 111, 51, 37, -102, -48, -92, -123, -7, 87, -40, -54, -71, -97, 108, -3, 98, -79, -14, 79, 70, 71, 113, 67, -121, -44, 105, 98, -112, -73, 12, -50, 26, -40, 16, 127, 51, -16, -97, 52, -68, 34, 104, 24, 70, -115, 113, -61, -51, -87, 75, 127, 29, -111, -110, -22, 60, -90, 54, -110, 1, 21, 77, -22, -99, 54, 40, 108, 53, -39, -20, -18, 77, -114, 81, -73, 72, 44, 100, 83, 126, 12, 22, -21, 78, -43, 41, 59, -124, 39, 117, 8, -103, 104, 88, -100, -76, 40, -9, 65, -73, -94, -21, -121, -19, -19, 112, -10, -3, 22, 86, 25, 104, -83, 73, 124, -58, -79, 83, -81, -83, 110, 34, -96, -90, 15, 94, -120, -20, 23, -96, 33, -100, 37, 14, 68, 83, 59, 64, -40, -90, 27, 82, -96, 35, 37, 102, -107, -26, 121, 94, -121, -42, -23, -19, 79, -92, -50, -33, -104, 59, -59, 9, 60, 101, 87, -32, 28, -90, 77, -39, 59, 38, 50, 87, -88, -39, -98, 43, -66, -24, -32, 93, -43, -117, 19, -100, 67, -75, 53, 72, 115, -27, -22, 84, -92, -118, 108, 91, 117, -54, 21, -70, -64, 105, 79, -108, -34, -64, -118, 88, 43, -82, 96, 70, 75, 13, -76, -24, -88, 70, -63, -41, 60, -74, -97, -72, -58, 37, 20, -86, 89, 54, 79, 114, 5, -73, -44, 115, 83, 96, 86, 2, 102, -62, 75, -44, -128, 7, 29, -41, 21, -2, 63, 35, -90, 9, 96, -12, -62, 82, 47, 53, 32, -30, -46, -128, 83, 90, 35, -3, 40, -126, -50, -18, -32, -1, -69, -84, -25, 114, 24, -76, -34, -36, -127, -43, 115, 91, 64, 122, 59, 36, 125, 48, -69, -109, -43, 115, -40, -106, -27, -12, -78, -37, 52, 119, -31, 64, 27, 8, 96, -90, -33, 61, -92, 119, -105, -13, -25, -100, 29, -75, -26, -6, 50, -128, 19, 48, 83, 37, 30, -68, -9, 93, 72, 56, 82, -32, -74, 35, 37, 13, 3, 18, -77, -102, -107, 79, 7, 25, 86, -19, -59, 27, -34, 26, 16, 1, -108, -95, -86, -103, 51, -43, 66, 68, 58, -107, 36, 10, -47, -56, -50, 59, -79, 37, -107, 63, 84, 125, -95, -2, -19, -59, 52, 83, -69, 71, 102, 86, 32, 121, 25, -109, 93, -24, 65, -64, 6, -90, 15, 80, 66, 111, -120, 41, 72, 16, -7, 121, 51, -76, 31, 93, -109, -8, -121, 60, -84, -2, 15, -49, 68, 29, -15, 40, 74, 44, -93, 79, -115, 87, -112, -122, 89, 52, -2, -94, 111, 123, -110, 99, 44, -12, -93, 31, 13, 36, 23, -80, -37, -33, 116, 8, 107, -17, -126, 116, -119, -114, 59, -32, -109, -38, 95, -76, 47, -20, 49, 108, 91, 118, 121, -9, 91, 32, 0, 41, -14, 67, -65, 12, 109, -6, 45, 80, 57, -35, -83, -108, 53, -27, -22, -19, 56, 116, -2, -66, -11, -113, 74, -51, -16, 104, -56, 56, 79, -71, 42, -58, 69, -38, -56, -112, -47, 35, 50, 35, -45, -18, -42, 106, 46, -102, 1, 0, -27, -75, 22, -87, 125, -56, -120, -33, -123, -128, 6, 60, -81, -45, 4, 21, -108, 46, -37, 72, 53, 104, -35, -60, 10, 52, 45, -52, -25, 36, -119, 108, 55, -122, -64, -33, 63, -29, 78, 54, 6, -44, -92, -72, 101, 121, -61, -41, -25, 78, -2, -10, 27, 22, -93, -69, 39, -112, 32, -114, -66, 95, -37, 42, 95, 4, -124, -59, -68, 21, 125, -124, -6, -114, 72, -53, 50, 72, 116, -109, 114, -62, 10, 92, 112, 10, 52, -116, 51, -15, 124, 98, 66, -97, 126, -97, -93, -45, 84, -99, 13, 58, 87, -78, 19, 93, -87, -71, -14, 33, -112, -44, -115, -63, -110, 113, 5, -118, -7, 116, 9, 82, 23, -118, 26, -57, 62, 5, -9, -19, -86, -89, -5, 86, -68, 83, -108, 79, -65, -81, -59, -33, -109, -88, 14, -39, 71, -107, -115, -104, 39, 13, 44, -71, 35, 111, 120, 99, 22, 85, -33, 57, 86, -121, -30, 50, -29, -11, -122, 23, 113, -41, 31, 46, -119, -84, 49, 90, -83, -5, 6, 47, -97, -76, 44, 53, -48, 107, -95, -4, -88, 102, -16, 19, 80, 126, -29, 109, 75, 110, 90, 17, -40, -104, 105, -56, -7, 27, -61, -25, -8, 126, -32, -39, 122, -119, 5, 28, -19, 97, 28, 35, -37, 94, 110, -41, 46, -124, 10, 27, 80, 12, 20, 98, 82, 10, -122, -123, 93, 65, 105, -67, 6, 31, 36, -15, -64, -64, 45, 52, -3, -72, -109, 82, 30, -85, -64, 33, 101, 87, 112, -83, -94, -120, 123, 104, 100, 116, -73, -70, -93, -6, -25, 75, 106, 98, 15, -48, -75, 60, -81, -74, 50, -90, 96, 22, 112, -35, -36, -48, -26, 93, -9, 10, -45, -41, 51, 4, 38, -80, -85, -75, 106, -52, -99, -6, 64, 76, 72, -35, 126, 56, 117, -103, 67, -90, 2, 16, -93, -38, 74, -39, -62, 1, -1, 17, -37, -117, -122, 87, 83, 98, -23, -45, 60, 39, -32, 58, 117, -112, -65, -15, -97, -83, 91, 109, 123, 12, 113, -12, -5, -64, -90, -12, 49, 25, -17, 67, 1, 92, -123, 105, -97, -119, 101, -67, 30, 34, -45, 0, -92, 89, -58, -127, 40, 89, -51, 64, 65, 31, 97, -118, 71, 84, -86, 66, 90, -53, 23, 99, -27, -4, 119, 78, 88, 116, -89, 121, 99, 4, 64, 88, -54, 83, 102, -8, -59, -62, -6, 65, -58, -70, 115, -94, -39, 16, 115, 83, -106, -18, 105, -14, 97, -8, -35, 125, 22, -66, 14, 70, 21, 59, -109, 109, -118, -28, -55, 119, 13, 48, -58, -89, -118, -56, 59, -46, -82, -124, -65, 44, 9, 96, -90, 74, -12, -36, -72, -70, -16, 83, -103, 94, -58, 63, -4, 5, 124, 35, 96, 38, 41, 125, 46, -88, 16, 44, 65, -47, -82, 78, 85, 64, 92, -78, -115, 114, 38, 41, -119, -10, -36, 64, -21, 87, -51, -70, -21, -47, 108, 70, -66, -31, -104, 63, -127, 99, -103, -3, -117, -126, -6, -18, -94, 115, -12, 116, 122, -57, -31, -8, -76, -23, 31, 57, 84, 89, -35, 87, -28, -83, -60, 94, 45, 64, 77, -58, 44, 55, -57, 100, 40, 72, -109, -25, 14, -11, 70, -126, 73, -21, -73, 86, 93, 118, -29, 8, -124, 36, 28, -62, -81, -79, -64, -49, 127, -42, 114, -98, -58, 19, 61, 33, -45, -100, 113, -56, 61, 0, -89, 124, 115, 49, 31, 57, -97, 47, 103, 37, -58, -82, 102, -86, -48, 119, -73, -71, -65, -59, 98, 73, 7, -69, -51, -38, -107, -102, -14, -87, -6, -63, -25, -5, -96, -84, -68, -123, 102, -99, 68, 3, 74, -77, -46, 50, 70, 47, -62, -76, -22, 45, -88, 6, -66, 26, 101, -15, 114, -36, -54, -6, 95, -113, 27, -46, -45, 46, 64, -28, -109, 29, -98, -70, -16, 75, -110, -34, -65, -17, -112, -16, 6, 32, 85, 50, -16, -84, -84, 58, 124, -43, -111, -11, 0, -37, -88, -27, 73, 99, 121, -21, 15, -88, -88, 42, -9, -117, 56, -43, -109, 79, -76, 67, -126, -76, 116, 53, -60, -128, -47, 40, 6, 82, 127, 22, -11, -94, -1, -13, 58, 120, -107, 39, 91, 112, 126, -82, -102, -79, -59, -77, 91, 36, 63, -88, 108, 113, 47, 118, 98, -75, -19, -40, 58, -119, -59, -75, 30, 59, 99, 127, 53, -80, -55, 8, -23, -96, -64, 42, 9, -22, 112, 57, -44, 115, -113, 88, -105, -48, 18, -9, -58, 112, 6, -32, 115, -121, -11, 69, -20, 98, 55, 2, 99, -118, 29, -35, 35, 79, -2, -84, 126, 117, -11, -127, -88, -104, -30, -47, -123, -33, -117, 78, -11, 46, -79, 86, 56, 95, -54, 105, -79, -73, 113, 125, 82, 91, 49, 118, 116, -127, 25, 123, 30, 122, -75, 96, -101, 86, -58, -127, 6, -43, 64, 52, -109, 35, -21, 22, 101, 28, -31, 90, 123, -13, 119, -34, -84, -91, 55, -47, -33, 70, 18, -124, -21, 49, 43, -19, -125, 21, -105, -119, -103, 123, -93, 64, -126, -47, 99, -46, -7, -16, -91, 49, -43, -25, -34, -78, -95, 50, -102, -51, -67, -93, -82, 8, -70, -96, 44, 27, -13, 37, 109, -32, -115, 81, 66, 103, 1, -84, -113, -83, -21, -76, -89, -14, -123, 117, -16, 86, 66, -24, 111, 118, 34, -68, -65, -121, 69, 118, -77, -53, 79, 122, -24, 4, 120, 99, -68, 62, -5, 7, 54, -61, -67, 29, -49, -77, -61, -43, 87, -80, 82, 121, 3, 43, -114, -78, -33, 63, 21, -35, 60, -78, 59, 69, 119, 118, 119, 32, -102, -106, -6, 95, -87, 29, -112, -5, 4, -12, 37, 52, 88, -115, -108, -87, 1, -63, 106, 121, -13, -121, -52, -4, -56, 70, 58, -8, -81, -13, 26, 24, -56, 113, -43, 40, 118, -99, 106, -128, -59, 36, 61, 40, 104, -27, -128, -1, 97, 85, 47, -24, 14, -46, -67, 103, -32, 46, 22, 93, 85, 77, 18, 89, -106, -87, 22, -54, -78, -110, 14, -107, -120, 56, 106, 76, -79, 126, -89, 80, 77, 53, -114, 27, 110, 45, -127, 26, 79, -93, -70, 45, 103, -9, -121, 42, -88, 45, -28, -127, 92, 74, 75, -17, -38, -114, 28, 4, 84, -103, -92, -50, -56, -65, -92, 1, 102, -32, 91, -64, -120, 115, 109, 39, -75, -120, -101, -125, -64, -83, 72, -68, 30, 94, -97, 54, -17, 44, -119, 37, -44, 66, 13, 28, 77, -118, -20, -38, 104, -34, -43, 36, 37, -8, 125, -125, 60, -64, -58, -46, -50, 116, -51, 13, -83, 123, -96, 41, -7, 120, -113, -63, 88, -126, -30, 19, -51, 17, -107, 5, 15, 85, 32, -49, -102, -108, 99, -67, -116, 50, -105, 30, 93, 52, 17, -74, 58, -28, -85, -75, 71, -57, -59, -106, -116, 111, 3, 106, -74, -27, 41, 102, -43, 7, 59, 79, -111, -50, 92, 27, -104, -69, -92, 94, 114, -110, -43, 9, 98, 124, 21, 83, 109, 32, -14, 94, -97, -85, -2, 56, -53, -26, 108, 126, -104, -95, 28, 33, -80, -34, 98, 38, 71, 75, -71, 30, 59, 126, 43, -111, 120, 119, -47, 38, 76, -95, -64, 39, -104, -71, 12, -116, -4, 74, -53, -74, 91, -32, 30, -82, -88, -30, -93, -19, 41, -53, 20, -102, 109, -115, -28, -16, -77, -66, 0, 20, 94, -98, 49, -5, -62, -36, 120, -7, -41, 126, -116, 87, -100, -38, 2, 67, 10, 36, 46, 86, -18, -104, -90, -29, -17, -87, -118, -114, -69, 48, 75, -101, -33, -115, -37, -87, 57, 70, 86, -77, -3, -108, 11, 86, -21, 54, 3, -91, -63, 125, 49, -109, 1, 62, -112, -57, 18, 19, 121, -99, 19, 112, 81, -10, -22, 91, 64, -119, 102, 109, -71, -4, 7, 126, -82, 59, -17, -85, -122, 41, 113, 118, 4, 72, 11, -4, 96, 122, -80, 33, -43, -120, 35, -37, 49, 27, 12, -80, 46, 3, 5, -82, 126, 55, 124, 98, 120, -94, -77, 64, -28, -99, -76, -125, -118, 101, 12, -49, -84, -77, -25, -118, 98, -73, 48, 71, -23, -98, -19, -41, 43, -98, 92, 93, 25, -102, -110, 0, -88, 108, 38, -46, 37, -36, -38, 8, 22, 78, -27, -16, -30, 11, -55, -97, 18, 96, 43, -112, 20, -121, -125, -53, -91, -124, -35, 115, -68, 81, 27, -123, 7, -15, -105, 104, -116, 89, -54, -51, -23, 118, 81, -56, 50, 23, 126, 41, 26, 51, 1, 59, -36, 81, 59, -40, 20, 117, -117, 112, 66, -10, 80, 113, 49, 58, -113, -41, -92, 43, 118, -46, 79, 0, 114, 20, -41, -108, 68, -112, -8, 7, 7, -62, -80, 94, -81, 111, -55, -91, 30, 12, -92, -69, -109, 79, 37, -122, 2, 94, 105, -78, -34, 74, 17, -99, 76, -60, 63, 36, -84, -96, -126, -70, -77, -30, -14, -40, 117, -74, 35, 63, 87, -46, 122, -56, -106, 55, 60, -4, -49, -11, 59, 124, 95, -112, -32, -34, 78, -97, 122, -56, -32, 8, 35, -87, 12, 36, 54, -2, 61, 30, -32, -58, 2, 120, -128, -29, 38, -66, -127, 7, -79, -22, 30, 67, 28, -104, -103, 6, 110, 116, -111, -8, -20, -117, -29, 84, -85, -66, 43, 107, -121, 112, 125, -75, 57, -12, -10, 0, -38, -117, 27, 117, -45, -48, -116, -1, -119, 122, -56, 50, -110, -108, -127, 60, -120, 51, -46, -120, -82, -88, 93, -104, 43, 118, -67, 48, 102, 42, 109, 16, 1, 75, 88, 26, 11, 0, 4, 28, 116, -122, 104, 9, 80, 59, 24, 100, 126, 23, -31, 16, -6, 53, -66, -91, -122, -112, 37, -97, 27, -74, 58, 48, 66, 64, -19, -11, 31, -12, -44, -64, -121, 38, 126, 30, -100, -110, 78, -107, -96, -60, -86, -39, -74, 57, 97, -122, -94, -119, 66, -61, 30, -93, -70, -117, -57, -113, 30, -29, -126, 123, -84, -90, -39, 58, -33, 30, -83, 14, -106, 30, 125, 14, 127, -125, -114, -110, 88, 19, -74, -102, -95, -35, -101, -40, -107, 53, 114, 29, 10, 22, 106, -67, 121, -102, -68, -12, 10, 41, -72, 73, -89, -9, 36, 96, 119, -35, 117, -25, 105, -66, -23, 26, 20, -124, 70, -92, 1, -13, -67, 124, 108, -18, -103, -79, 35, -11, -36, 26, -101, 120, -19, 123, -70, 3, 49, -3, 66, -73, -104, 92, 79, -47, 70, 111, 40, 32, 124, -6, 9, -60, -123, 36, -54, -80, 99, 21, 36, -103, -60, -123, -117, -60, 113, -67, -92, -13, 22, 84, 11, -111, 107, -7, -125, 32, 84, -35, -40, 32, 100, -59, 57, 19, -25, 23, -111, 88, 50, 1, 95, -90, 123, 8, 101, -59, 36, -13, -105, 16, 25, -43, 54, -88, -92, -61, 60, -23, 38, -52, -43, 61, 25, -86, 98, -86, 31, -58, 15, 27, -61, -115, 11, 121, 36, 104, 88, -9, 74, -35, 106, -119, 1, 98, 14, 32, 112, 93, 24, -65, -10, -49, 71, -72, 122, -86, 71, -125, -75, 97, 124, 31, 124, -52, -68, 67, -93, -5, -36, 51, 41, 122, 3, -95, -112, -84, -101, -80, -18, -127, -7, -32, 127, 74, -75, -103, -101, 124, -74, -70, 93, 80, 115, 60, -41, 10, -85, -20, 37, -23, -95, 89, 79, 32, 19, 23, 20, 55, -107, 107, -128, -9, 75, -128, -118, 26, -39, -60, 101, 27, 124, 83, 29, 111, -124, 10, 75, 100, -94, -11, 104, 16, 57, -3, 49, -119, -96, -69, 93, 65, 55, 86, 71, -47, -90, -37, -120, 90, 107, -53, 0, 17, 81, 111, 57, -120, 0, 91, -16, -20, 64, -90, -105, -61, 93, 120, -56, 64, 47, -70, -34, 53, 8, -46, 105, -99, 19, -36, 80, 12, -90, -39, -49, -53, 20, 10, -1, 81, 64, 58, 20, 42, 39, 30, -127, -20, -37, -117, -3, 66, 5, -126, -126, 96, -127, 84, -125, -24, -11, 81, 107, -59, 83, -67, -40, -2, -89, 126, 71, -73, 45, 28, 109, 14, 64, 72, 53, 31, -56, -76, 12, 84, 77, 30, -95, 11, 78, 102, 32, 74, 127, 37, 97, -8, -27, -26, 64, 96, 110, -1, -62, -29, 110, 28, 98, -41, 27, -43, 55, -53, -81, 72, -125, 26, -13, -103, 2, -110, -120, 10, 1, -70, -31, -35, 36, -12, 124, -50, -38, 1, -82, 120, 74, 50, 5, -71, 56, -96, -103, -75, -51, -74, 19, -14, 110, 68, -56, -43, -98, -125, 91, 12, 105, -66, -87, 45, -99, -21, -31, -53, 108, -45, -124, 107, 16, -110, 60, -89, -118, -93, 64, 98, 14, 34, -74, -29, 66, 7, -112, 49, 125, 112, -11, 48, 82, -31, -108, -121, 21, -101, -17, -55, 105, -72, 32, -12, 104, 83, 19, -13, -52, 105, -87, 68, -34, -5, -1, 4, 64, -106, -43, -40, -95, -68, -6, 14, 61, 48, -88, -66, -124, -17, -38, 111, -40, -89, 105, 17, 101, -128, -81, 13, -46, -49, 49, -23, 18, 107, -82, -75, 69, 122, 79, -101, 52, -125, -70, 80, -100, -18, 79, 0, 108, -110, -115, -47, -34, -31, -80, -66, 89, 83, 42, 36, -4, 116, 33, -80, 111, 23, -35, -21, 13, 51, 55, -5, 60, 109, 12, -116, 111, 121, -16, 73, 100, -121, 42, -127, 115, 21, 3, -89, -94, -99, -112, 4, 28, 37, -56, -25, 30, 93, -117, -108, 25, 88, 83, 68, 108, 49, -126, 26, -16, 38, 80, -19, -119, -77, -60, -119, 20, -12, 4, -112, -117, 30, 107, 68, -73, 86, 113, -75, 5, -109, -45, -56, -97, -27, 41, 8, -123, 47, -33, -17, 58, 1, -105, 66, -89, -124, 27, 56, 7, 70, 104, -98, 104, -103, 64, 111, -117, -2, 97, -19, 63, 77, -37, -125, 65, -83, 89, 97, 52, 55, 78, 120, 74, 124, 12, 50, -107, 95, -114, -38, -99, -76, 48, 34, -71, 126, -13, -75, -57, -50, -112, -111, 37, 97, -44, -80, 108, 1, -67, -83, 66, 76, 59, 54, -24, -103, -57, 40, -94, -50, 93, 64, -75, -73, -79, -32, -72, -105, -45, 32, 49, 77, 93, -31, -122, 81, -123, -15, 16, -110, -93, 47, -59, 61, -69, -51, -84, 28, 33, 102, 110, -128, -73, 24, -53, 59, 1, 34, 44, 77, 35, -22, 34, -124, 126, 10, -36, -61, 101, -52, 11, 114, 5, -113, 24, -35, 33, 53, 123, 81, 43, -124, -105, -54, -14, 57, 58, -4, 122, 110, 71, -38, -26, -48, -13, -12, 6, 46, 17, 85, -80, 4, -55, 17, 115, 52, 41, 122, 115, 47, -104, 46, -114, -97, 102, -55, 28, -37, -19, 45, -87, -119, 76, -100, 93, 35, 90, 90, 4, -85, -6, -79, -51, 49, -39, -73, 6, -113, 64, 124, 63, 41, -45, 99, -45, -88, 56, -124, 62, 18, -88, 109, 36, -69, 91, 124, -77, 103, 17, -30, -48, -17, 40, 63, 9, -53, 101, -106, -119, -10, -104, 106, -82, 124, -93, -30, 3, -94, -93, -34, -75, 126, 73, -59, 56, 36, 54, -9, 65, -125, 15, -32, 116, 2, 123, 125, -86, 29, -104, -69, 46, -39, -96, -28, -115, -27, 1, -125, -42, 67, 38, -121, 38, -110, 18, -116, 126, 105, 62, -62, -126, 94, 62, 110, -45, -113, 81, -59, -118, 83, 100, -37, 36, -12, -112, -68, 36, -60, 114, 3, 15, -113, -108, 64, -40, 39, -73, 43, -126, -108, 98, 25, 18, 32, -45, 78, 126, 19, -109, 112, 107, 16, -91, -21, -78, 54, -98, -89, 111, 61, -96, -34, 14, -68, -3, -58, 100, -34, -10, -25, 81, 67, 28, 91, -120, 21, 107, -25, 63, -74, -61, 26, -98, -95, 121, 58, 73, -40, 110, 77, -24, 102, 89, 123, -29, 109, 95, 24, -21, -38, 59, -44, -12, 110, -64, -86, 5, 28, 56, -90, -76, -23, 68, -36, 59, -87, 40, 94, 95, 84, 88, -39, 63, -59, -32, 8, -110, -6, 22, -108, 47, -112, 8, 91, 17, 27, -68, 115, 25, -94, 31, 51, -86, 17, -14, -84, 36, 37, -7, -103, 119, 123, -26, 77, 2, 86, -98, -51, 76, -42, 121, 125, 29, -12, -10, -58, 88, 0, 86, 39, -99, -90, 41, -107, -50, -82, -24, 105, -90, 46, -115, 94, 79, 28, 72, 89, -29, -118, 13, 74, -88, -39, -67, -16, -53, 54, -66, 101, -35, 53, -43, -13, -17, -57, 37, 102, -51, -64, -87, -59, -49, 100, 54, 80, -43, 55, -52, -27, -25, -16, 73, -65, 26, -66, 19, -12, -20, -71, 24, -106, 66, -94, 51, 50, 70, 122, 121, -32, 73, -88, -59, -108, -79, 61, 23, 55, 75, 77, 59, -5, 69, 56, -17, -21, -74, 120, -99, -81, -34, 30, 46, -59, -79, -23, 118, -53, -36, -115, 122, -63, -71, -104, -91, 10, 72, -120, -19, -94, -99, -44, -64, 27, -49, -49, -1, 106, 84, 30, 5, 52, -14, 7, 2, 7, -19, 65, 94, 35, -28, -118, -98, -25, -39, -58, -30, -84, 126, 83, 59, -12, -43, -109, -4, 38, 92, 34, 24, 30, -104, 121, -89, -36, -5, 119, -96, -121, -121, 71, -30, 25, -13, 57, -54, 99, 12, -39, 62, 61, -94, 14, -125, 103, -123, -83, 59, 0, -110, 29, -98, -76, 42, -60, 37, 124, -97, 113, 38, 39, 127, 78, 17, 53, 19, 28, 106, -76, 72, -53, 8, -123, -107, -2, -15, 49, -68, 58, -31, 77, -45, 7, 48, 86, 38, 69, -23, -18, -46, -72, -103, 20, -94, -124, -114, 55, 0, 85, -49, -54, -66, 34, -114, -52, 28, -63, 103, -112, -35, -23, -14, 13, 123, -115, 0, 80, 85, 29, -1, 51, 11, 121, 84, 127, 36, -59, -51, 15, 61, -63, -48, 106, 55, -11, 14, 8, -109, 110, -15, -50, 73, 120, -92, -115, 29, -39, -111, -32, -13, -19, 51, 114, 47, 13, 109, 85, 125, -4, -61, 13, -109, 73, -25, 109, 70, -90, 55, -26, -124, -27, -24, -17, -112, 89, -97, 36, 32, -62, 4, 49, -1, -55, -88, 24, -48, 122, -128, -6, 95, 100, -87, 62, -87, -70, 12, 88, -103, 111, -75, -27, -88, 20, -12, 76, 115, -18, -54, -22, -28, 98, 90, -91, 40, -39, -29, -94, 61, -15, -55, -7, 101, -81, 53, -1, 110, -38, -125, 109, -7, 94, 102, -88, 16, -31, 118, -104, 69, -115, -2, -77, -39, 8, 5, 22, -1, 73, 107, 32, 91, 84, 0, -3, 109, -85, -69, 54, -120, -68, 110, 59, -43, -61, 75, 120, -84, -85, 3, -55, 100, 3, -84, 35, 114, 22, 71, 109, -74, -101, -26, 56, -113, 115, -121, -63, 70, -127, 28, 67, 94, -13, -30, -36, -109, 29, 32, -80, 124, 96, 48, -77, -13, 1, -63, 127, 114, 37, -1, 38, -87, -92, -28, -30, 104, 16, 0, -13, -107, 33, -9, -26, 13, 4, -10, 44, -94, 49, -117, -35, -29, 126, -36, 106, 32, -32, 10, 5, 68, -2, 3, 13, 110, -99, 18, 116, -126, -86, 44, 104, 28, 85, -86, -99, -127, 121, -105, -116, 15, -58, -66, -51, -109, -88, -90, -20, -33, -68, 32, -16, -28, 89, -90, -101, 80, -21, 94, -41, 86, -6, -4, 73, 18, -22, 35, 56, 118, -16, -128, -71, 37, 84, 79, 106, 125, -51, 101, -92, 6, -84, 92, -26, 18, -7, -9, -40, -91, 46, -60, 4, -127, -122, 110, -32, 28, -28, -120, -104, -80, 60, -120, -50, 9, 13, -25, 40, -91, 25, 29, 82, 92, 119, 14, 112, 109, 84, 50, 30, 59, 86, -112, -119, -90, 120, -2, -106, 122, -4, -85, -47, 38, -68, -20, 114, -121, 112, -38, 122, -95, -117, 107, 111, 127, -36, -112, 34, 22, -61, 76, 1, 28, 87, 110, -56, -10, -57, -66, -75, 105, -122, -84, -28, -107, 94, -124, -5, 0, 26, 68, 127, -92, 3, -37, 40, 46, 31, 52, 29, 56, -16, -99, -29, -44, 17, -40, -14, -69, 46, -80, -29, 25, 23, 114, 105, 70, 81, 71, 103, -83, 20, -65, -13, 50, 26, -61, -79, 90, 112, -44, -23, 107, -42, -21, 43, -104, -21, 30, -10, 72, 116, 17, -99, -76, -48, 0, -50, 90, 42, 83, 21, 127, 58, 65, 37, 46, -81, 121, 17, 40, 47, 21, -103, 27, 111, -118, -16, -64, -92, 40, 41, -69, -43, -70, -42, 9, 30, 54, 124, 85, -29, -5, 120, 5, 24, -73, 45, -109, -7, -108, 113, -96, -52, -1, -106, 82, 102, -34, 124, 118, 118, -50, 86, 115, -127, -19, 75, -70, 107, 78, -26, 77, -20, 39, 123, -122, -62, 42, -15, 58, -22, 90, -7, 71, 95, -13, 86, -59, -116, 69, -31, -9, -28, -45, 76, -81, -21, -90, -124, 4, 32, -120, 2, -9, -112, 82, 88, 32, -52, -106, -66, -117, -85, 91, 74, -21, 35, -109, 14, 86, -26, 119, -3, 92, 121, -26, -106, -25, 14, -54, -61, 28, -26, -102, -18, 45, -18, 66, 35, -93, -29, 16, 37, -97, 110, 109, -20, -84, -118, -104, 3, -116, 76, 64, 88, -55, -2, 12, -109, 127, -14, -78, -90, 127, 93, -61, 74, -99, 35, -107, -53, 14, -114, 118, 45, -24, -27, 13, -88, 104, 26, -114, 96, -9, -44, -62, -18, 46, -13, 57, -80, -22, -99, -8, -80, 47, 80, -122, 19, 19, -121, -54, 120, 118, -115, 89, 82, 100, 4, -112, -58, -126, 108, -9, -112, -81, 39, 27, 78, 38, 83, -101, 124, -19, -90, 112, 67, -45, -21, -91, -63, -22, -96, -47, -71, 20, -125, 69, -112, 27, 60, 124, 28, 25, 7, -127, -18, 114, -75, 54, -26, 73, 127, 7, -75, -7, -44, 75, 95, -76, 44, -120, 120, 56, -72, 44, 27, -98, -92, 127, -111, 109, -30, 24, 91, -98, 111, 33, 61, 107, -45, -45, -46, 45, -93, 11, -47, -1, -91, 107, -18, -117, -92, -108, 89, -125, -114, -1, -50, 56, 19, -51, -26, -73, 16, 2, 95, 107, -36, -26, 57, 45, -122, 20, 58, -94, -96, 27, 113, 65, 72, 72, 59, 91, 5, -105, 43, 118, 54, 97, 8, 30, -88, -106, -113, 46, -97, 87, -97, -97, 119, -28, -81, 7, 72, -103, 63, -112, -27, 49, 81, 37, -43, 8, 73, -78, -22, -111, 63, -105, -37, 77, -115, -34, -41, 72, -125, -76, -120, -26, -73, -77, 115, -16, -97, -33, 39, 87, -11, -112, -2, -119, -64, 126, 65, -92, 101, 58, 77, 127, 34, 51, -114, -5, 24, 43, -36, -26, -71, 32, -63, -73, 7, 44, -87, -63, 103, 20, -19, -24, -41, 7, 119, 1, -54, -51, 47, 106, -119, -73, -19, 7, -120, -54, 115, -62, 114, -98, 2, 35, -17, -113, 57, -68, -15, 100, -26, 87, -10, -64, 85, -74, -41, 3, 44, 24, -63, -18, 24, -51, -116, -4, -78, 27, 108, -74, -117, -38, 77, -110, 82, -37, 112, -17, -33, 71, -8, 96, 101, -67, 57, 16, 58, -38, 111, 97, 81, 28, -27, -42, 105, -24, 7, -127, 49, 29, -109, 11, -16, 121, 15, 17, 111, 123, -29, -114, 94, 111, -49, -69, 56, 50, 112, 118, 78, -43, 10, 35, 101, 72, 118, 108, -31, 63, -48, -69, -69, 62, -69, 6, 108, 114, -128, 100, -18, -97, 19, -89, -7, 19, 84, 11, -25, -15, 79, -29, 79, -116, -47, 55, 66, -82, -58, 93, -81, 35, -69, 68, -96, -6, -68, 108, 22, -41, 89, 53, -32, 92, 83, -42, -85, 87, -28, 90, -22, -114, -14, -72, -35, 44, 15, -25, -20, -1, 101, -67, -79, -90, -1, 51, -75, 5, -28, -62, 25, -13, -27, 67, -84, -23, -62, -22, -114, 28, 11, -66, 69, -50, 65, 97, 109, -118, 57, -91, -12, 74, 115, 103, -58, 74, 78, 60, 82, -45, 91, 95, 124, 4, -59, -23, -58, 68, 98, -85, -113, 86, -119, 99, 10, -93, 21, 25, -77, 111, -93, -70, 79, -39, -11, 92, 79, -22, 121, 12, 116, -24, 39, -14, 114, -66, -69, 78, 83, 51, 15, -27, -68, 23, -12, -116, -3, 90, -1, 56, 1, 92, 82, -16, 71, -64, -125, -12, 116, 73, -104, 105, -60, -128, 84, -80, 90, 29, 98, -120, -84, 90, -77, 117, 53, -99, 17, 18, -124, -82, 39, -107, -122, 69, 101, -122, -46, -10, -75, 122, -103, 49, 99, 0, 49, 18, -108, -47, -28, -70, 62, -44, 121, 127, 29, -48, -114, -98, -7, 88, -5, 101, 97, -23, -47, 114, 87, -64, 91, 66, -88, -69, -47, 14, 25, -73, 121, 66, -40, -50, 95, -83, -122, 40, -46, 66, 95, -60, -85, 64, 38, -28, -49, -120, 57, -92, 117, -43, 82, -73, -59, 52, 41, 34, -23, -120, 94, 31, -105, 90, 40, -34, -30, 104, -57, 27, 88, 21, 4, 118, -106, -5, -31, -92, 10, -73, 7, 99, 84, -78, -97, 72, -54, 61, 48, 12, 41, 55, 126, -21, -127, 27, 12, 82, -30, 57, -37, -104, -112, 92, 29, -100, -81, -10, 103, -22, -83, 102, 90, -70, -85, -112, 86, 97, 113, 84, 119, -116, -10, -39, -120, 8, -28, -14, -107, 54, -38, 23, 69, -2, 9, -115, 87, -9, 2, 29, -98, 54, 98, 112, 97, -42, -119, 48, -41, 126, -48, 80, 122, 78, -89, 10, -54, 45, 9, 16, 90, 27, -127, -33, 17, -62, 29, -50, 68, 13, 31, 55, -47, -4, -74, -28, -2, 119, -50, -110, -13, 110, 58, 11, 90, -23, 89, -31, -19, -127, -106, -103, -66, 31, -46, -100, -22, 117, -71, 8, -28, 126, 113, -78, 92, -23, 86, 105, 31, 44, 93, -18, -31, -104, -39, -74, 27, 126, 49, -84, -97, -27, -82, 26, 12, 57, 95, 2, 70, -67, -38, 114, -117, -114, -118, 87, 105, 63, -21, -124, -29, -38, -115, 97, -69, 39, -114, 101, 9, -60, -82, -50, 29, 125, 18, -70, 9, -100, 25, 28, 47, 25, -70, -18, 1, -70, -41, -37, 105, -39, -10, -69, -89, 96, 104, 10, -67, -90, -79, 50, -98, -94, -28, -80, 30, 117, -24, 86, 111, -121, -78, 18, 96, 40, -62, -14, 91, -35, -46, 109, -37, -74, 116, -17, 68, 115, -67, -118, -76, -80, 119, -128, -97, 104, -25, -32, 79, -99, -121, 46, -123, -53, 117, 84, -30, -82, 95, 116, 89, 94, 93, -109, -112, -115, -19, 114, -94, 104, 0, 79, 37, 64, -26, -106, 25, 62, 58, 104, 20, -11, -55, -12, 116, -24, -88, -14, 123, -124, 125, -11, -89, -57, -124, 70, -63, -125, 47, 76, -62, 127, 109, -92, 11, -81, -77, 25, 90, -58, -29, 60, -126, 41, -74, 96, 121, -64, 110, 127, 30, 25, -11, 78, 95, 32, 118, -26, -88, -15, -28, -66, 122, -66, 10, 100, -64, 45, 93, 5, -71, -95, -114, 122, -24, 61, -82, 72, -39, -26, 71, -41, 102, 31, 11, -102, 97, -4, 125, -93, 116, -46, -33, -103, 105, -96, -121, 25, 49, 90, 58, -1, -74, 57, 30, 18, 32, -120, -103, -122, 114, 27, -104, 23, 44, -88, -92, -73, 127, -17, 107, 11, 32, 90, 89, 47, -50, -92, 74, 66, 69, 76, 124, -108, -74, 93, -24, 46, 63, -55, -43, -83, 114, -98, -80, 13, -41, -51, -13, -127, 112, -57, -99, 107, 102, -2, 28, 42, 119, -54, 93, -109, 11, -58, 84, -38, -41, 2, -102, 76, 115, -93, 38, -13, -77, -7, -23, 38, 91, 91, -107, -96, -14, -41, -48, 8, 73, 91, -9, 21, -91, -96, 82, 99, 26, 100, 24, 25, -50, -89, -84, -19, 19, -38, 63, -20, -19, 121, -128, 24, -104, -45, 95, -68, -99, -48, -106, 14, -28, 77, -106, -105, 99, -66, -32, 32, -50, -16, 27, 54, 99, 123, 73, -41, -124, 24, 90, -26, -58, 86, 73, -88, 58, -34, 4, -7, -102, 69, 20, 80, -17, 96, 75, 42, -4, -36, 47, -87, 8, 17, 118, 44, 46, -19, -111, 39, -84, 63, 15, 83, -119, 89, 70, -77, -39, -58, -47, 70, -26, -47, -121, -45, -46, -52, -90, -34, 95, -110, 81, -75, -82, 89, -126, 93, 28, -2, -101, -55, -90, 65, -119, -95, -20, 99, -50, -93, 72, -4, -68, 4, -17, 116, -40, -60, 36, 88, -103, 118, -20, -27, -3, 62, -113, 27, -83, -3, -113, -8, -108, -83, -58, 21, 38, 52, 122, 12, -101, 121, 47, 112, 52, -117, -33, -58, -15, 102, 79, 12, 96, -25, 110, -80, 126, 34, -46, -34, -6, 33, 91, 42, 63, -121, -18, -116, -72, -80, -126, 34, 3, -111, 79, -50, -81, 32, -128, -62, 43, 72, -7, -128, -32, -99, 2, 98, -65, -89, 71, 114, 11, 60, 65, -40, -51, 47, 56, -81, 122, -37, -38, -37, 34, 123, 53, 39, -23, 16, -119, -63, -13, -17, -37, -75, -4, -51, 85, -19, -115, 82, 59, -116, 83, -13, 39, -76, -63, 82, -123, -74, 64, 110, -16, 118, 31, -21, 107, 124, 6, -46, 58, 14, -66, 48, -30, -26, 93, -59, 114, 70, 96, 114, -46, -28, -17, 31, 57, -118, -124, 19, -7, -51, 27, 67, -105, -53, -46, -92, -21, 127, 120, -18, -37, -35, 98, -34, -34, -96, -36, 51, 108, 60, -110, -11, -34, 51, 20, -71, -106, 30, 24, -121, 62, 52, 5, 9, -26, 44, -71, 24, 78, 28, -122, 61, -1, -55, -66, 15, 112, 115, -78, -6, 79, -24, 29, -62, -80, 106, -20, 88, 54, -126, -109, 35, -123, -60, 126, -112, 56, 33, -41, 3, -106, 0, -120, 29, 107, 31, 54, -26, 17, 48, 87, 73, 27, -47, -16, -3, -59, 85, 32, 45, -117, -86, 68, 69, 61, 66, 32, 125, -114, 84, 80, 74, 38, -18, -64, -94, 15, 28, -62, 69, 65, -36, 34, -123, 66, 43, 80, -123, 56, 73, -92, -98, -91, 24, 62, -51, -48, 111, 39, 88, -82, -6, -120, -39, -116, -76, -122, 49, 12, 19, -62, 14, -5, -123, 103, -38, 67, 12, 63, 41, -1, 104, -71, 3, 102, -55, -88, 70, -89, -55, 16, -115, -104, -52, -96, 14, -115, -11, -7, -17, 115, 80, -38, 112, 17, -22, -62, 99, 53, 52, 115, -76, 42, -83, -90, -69, -90, -97, -12, 86, -52, -21, -24, -80, -109, 10, 19, 109, 33, -11, 121, 123, -22, 105, 81, -20, 11, 112, -12, 49, 44, -43, 8, 23, 127, 64, -29, 75, 111, -48, 44, 126, 111, -31, -56, -119, -73, 50, -34, -50, 125, 119, -39, -5, -89, 32, 113, -90, 15, -54, -25, 99, 19, 47, -92, 102, -121, 82, -115, 4, 39, -65, 110, -116, 9, -110, -124, -94, 100, 74, -37, 118, 16, 11, 91, 55, 48, -109, -76, -95, 56, -41, -67, 127, -87, -105, 65, -93, -55, -25, -63, 11, 58, 4, 12, -8, -6, 89, 86, 23, 82, 116, -107, 104, -75, 63, 67, -93, 17, 124, -96, -89, 88, -4, -32, 56, -13, 61, 8, 94, 52, 102, -81, -24, 51, 30, -76, -37, -109, 81, -76, -86, 32, 27, 73, -97, -7, 42, -41, -11, 26, -66, -115, 119, -93, 15, -54, 74, 35, -50, 37, 116, -125, -57, 12, 72, 87, 22, 86, -96, 8, 113, -34, -5, -101, 99, -23, -106, -99, -57, 32, -85, -26, 79, 83, 17, -116, 56, -30, -86, -91, 14, -23, 44, -69, 63, -34, -37, -58, 68, 127, -54, 86, 117, 12, -6, 103, 115, -126, -21, -67, -37, 36, -121, 125, 20, 45, 63, -106, 112, -32, 101, 48, -103, 117, -111, 96, 125, -53, 76, 15, -62, -97, 101, 60, 126, -65, 49, -26, -13, -49, 112, -69, -20, -76, -111, 0, 109, -15, -108, 15, -77, 67, 64, 33, 70, 125, -62, 60, -83, -126, -60, 45, -9, -124, -30, -10, 105, -92, 68, 123, -113, -42, 49, -61, 11, -43, 106, -52, 65, -96, 87, -46, 43, -97, 47, 84, -100, -115, -94, 10, -76, -105, -4, -55, -110, 96, -69, -20, 127, 90, -42, 22, 125, -102, -4, -48, -35, 1, 116, -41, 101, 77, 123, 126, -64, 40, 103, -93, -50, -57, 16, 1, -123, 60, -51, 126, -97, 4, 85, -42, -109, -21, 57, -24, -59, 62, 71, -78, 18, 19, 68, 127, 40, 12, 68, 30, 39, -114, 27, -74, 3, 36, 88, -79, 98, 111, 37, 103, 97, -127, 49, 120, 56, 99, -122, -34, 72, 54, -57, 95, 92, 116, 36, -24, 58, -68, 120, 81, -34, -86, 2, -25, 104, 49, -46, 40, -57, 47, -72, -89, -110, 80, -46, 92, 98, 107, -94, 37, 58, -112, -19, -119, -83, -99, -57, -5, 115, -1, 59, 34, -75, 105, -69, 120, -128, -19, 27, 20, 45, 66, -105, -116, -98, 113, -20, -61, -115, 123, -64, 123, -4, -3, 127, -70, 49, 75, -109, 26, -95, 34, 127, -11, -104, 74, 4, 44, -91, 83, -86, -99, 33, 36, 66, -12, 109, 31, 98, 97, 50, 33, -120, 110, 73, -51, 72, -17, -79, 48, 71, -37, -94, -65, 114, 102, 70, -74, -35, -90, 108, 125, -24, -97, 105, -45, 86, -12, -62, -57, 90, -120, 37, 48, -126, -47, 92, 119, 73, -62, 53, 52, -120, -73, 93, 16, -78, -70, 98, 48, -68, 92, -45, -23, 54, -3, -46, -10, 25, -42, -85, 120, -125, 24, -14, -108, -111, 7, -99, 48, 50, 23, -44, 106, 19, 61, -120, -49, -35, -82, 61, -3, 19, -25, -95, 28, -45, 62, 97, 4, 61, -104, 124, -125, 12, 82, -122, -75, -1, -60, 40, -55, -15, 20, -88, -126, 51, -115, 52, -68, 94, -114, 112, 4, 51, -4, -14, 37, 4, 124, -41, 72, -110, 85, -91, 21, 56, -33, 76, -40, -4, 124, 11, -3, -51, 28, -95, -114, 108, -123, -71, 101, 16, 87, -74, -53, -21, 52, -99, -119, 61, 9, 30, 85, 21, -94, -51, -2, -90, 12, 66, -52, 57, 38, -44, -60, -25, 68, -24, -64, 95, -119, -60, 55, 6, -125, -125, -105, -70, 103, -36, -85, -9, 73, 95, 82, -52, 86, -49, 97, -103, 38, -120, -61, -62, 15, 77, -66, 39, 119, -17, -108, 106, -71, 108, 57, 118, -71, 53, -26, 112, 6, -123, -1, 60, 121, -125, -59, -126, 95, -89, 86, 13, 46, -92, 21, -54, -59, 124, -37, -37, -43, -34, 14, -110, -56, 3, -10, -51, 104, -104, 40, -12, 1, -5, -26, -122, -11, -99, -4, -33, 75, 95, 28, -75, 36, -67, 109, -111, 40, -40, -30, -9, 12, -94, -45, -117, -61, 89, 46, 86, -118, 126, -8, 8, 121, -121, 89, -117, 53, 16, -93, -120, 29, 41, -69, 87, -76, -63, -5, -128, 105, -43, 47, -103, 36, -63, 106, -106, -107, 42, 68, -35, 15, 24, 7, -90, 6, 12, -111, 17, -102, 28, 33, -50, -36, -97, 61, -127, -76, -121, 93, -77, -110, -55, 117, -80, 69, 109, 76, 5, 30, -102, -103, -64, -87, -95, 119, -87, -3, 45, 8, 66, 29, -29, -110, -57, 120, 69, -60, -5, 115, 116, 86, 5, -92, 86, 105, 119, -58, 17, 35, 113, -14, -28, -19, 24, 58, -21, 13, 34, -100, -100, -56, -101, -83, 91, -96, -114, -10, -104, -35, 64, -67, -121, -33, 25, -50, -117, -23, 49, 10, 76, -78, -37, -10, -96, -110, -51, -10, -67, -55, -127, -73, -84, 66, 74, -75, -86, 94, 16, 69, -86, 5, -47, -11, -43, -48, 82, -51, 110, -117, 90, 113, -70, 73, 69, 88, 99, 93, 119, 110, 3, -80, 88, 117, -93, 105, 78, -45, 62, -80, 30, 117, 26, 99, -42, -103, -82, -83, 60, -23, 59, -29, 36, -64, -31, -44, 92, -34, 87, -48, -56, 102, -113, -6, 89, -28, -15, -90, -121, 51, -28, 84, -21, 61, -104, 57, 47, 45, 55, -22, -42, 24, 99, 40, 51, -45, 119, -26, 3, -26, -18, 42, 75, 98, 59, 94, -113, 79, 74, 4, 116, -82, -50, -15, 59, 56, -26, 114, -38, 14, 72, 44, -109, -85, 27, -12, 93, -127, 87, 6, 75, 37, -94, -26, -2, -103, 118, -106, -83, 14, -100, 12, -52, -55, -46, -62, -110, -27, -94, -14, 5, 83, -88, -33, 22, 106, -15, 54, -91, 47, -77, -120, 27, 3, 46, 86, -86, -125, 59, -117, -58, 65, -46, -31, 23, -4, -61, -41, 116, 54, -124, -113, 83, 70, -102, -20, 77, 116, -75, 63, -90, 25, 78, 13, -115, -82, -55, 5, -89, -113, -105, 51, 122, -67, 18, 67, -128, -18, 87, -11, 101, -102, -83, -117, -68, 55, 5, -81, 113, 25, -12, 84, 83, -15, -19, 116, -62, -11, 53, -78, 121, -48, 101, -127, 20, -86, 11, -112, -83, 102, -30, 41, 107, 18, -67, -86, 103, 124, 30, -78, 65, -72, -80, 63, -99, 2, 78, -98, 73, -61, -3, 89, 123, 40, 125, -114, 55, 45, 20, -106, 62, -12, 52, -104, 104, -95, -39, -73, 45, 121, -69, 99, -103, 81, 14, 103, 48, 4, -23, -80, -1, 39, 84, 110, -116, -76, -103, -74, -29, 103, -96, -41, -38, 114, 48, -71, 77, -21, -58, 114, -38, 99, 31, 77, 7, -113, 119, -92, 91, -38, 96, 68, -75, 78, -70, 114, 92, -78, 17, 113, 12, -89, -105, 8, -101, 33, -79, -78, -80, 18, -48, 49, -94, 56, -124, 44, 115, -46, -126, -27, 71, -14, -4, 18, -93, 17, 88, 4, 66, -88, 84, 0, -10, -28, -82, -61, -24, 97, 120, -40, 46, 112, 65, 89, 73, 43, -74, 26, -94, -48, -62, 105, -13, 71, -81, 123, -85, -47, 111, 119, 22, 55, -46, 125, 13, 21, -63, 68, -65, 25, 57, -78, -119, -14, -92, 16, -17, 0, -29, -5, -79, 46, -33, 40, -9, -90, 122, -75, 100, 61, -12, -86, 78, -103, 114, 122, -52, -65, 102, 99, 63, -6, -80, -91, 83, -5, 91, -32, -75, -53, 122, -95, 7, 5, -20, 112, 50, -83, 22, -85, 12, -29, 44, -103, -101, -84, -50, 122, -127, -32, -18, 72, 3, -126, 106, -93, 49, 55, -21, -18, 107, -114, -123, -128, -123, -76, 28, 95, -18, -79, -105, 109, 98, 18, -4, 71, 124, 3, 121, 69, -104, -109, -33, -21, -121, -75, -124, 15, 66, -123, 109, 69, -104, -74, -74, 105, -116, 50, -128, 93, -5, 124, -87, 19, 23, -66, 11, -16, 87, 3, -105, 115, 9, -15, -61, 73, -91, -16, 107, -113, 58, -77, 55, -114, 60, 45, -45, 10, -11, -65, 120, 95, -40, -128, -65, 62, 69, -76, -120, -17, -109, 124, 47, 118, -60, 86, 51, -76, -23, -103, 102, -16, 101, -115, -112, 61, 28, -95, 0, 45, -92, 2, -87, -29, -28, -53, -33, -57, 108, -92, -48, -63, -67, 86, 9, 37, 104, 23, 58, 124, -23, 126, 43, 74, -128, -92, -123, 23, 96, -121, 61, 25, 104, -12, 92, -68, 44, 85, -40, 67, 100, -124, -2, -17, 13, -50, 53, -123, -108, -50, -50, -66, -64, -101, 106, 34, -14, -42, -51, -46, 28, -35, -110, 124, 93, 98, -87, 10, 104, 33, 113, 120, 70, 49, -103, -59, 73, -121, 107, 49, -83, 14, -72, -33, -114, 30, 79, 40, -76, -99, -16, -104, 10, -39, 105, -85, 68, -96, -127, -17, -117, -22, 94, 126, 30, 102, 51, -63, -12, 82, -22, 117, -37, -99, -2, -114, -50, -49, -77, 125, 9, 110, 115, -44, -111, 103, 108, -74, 34, -54, 100, -61, 109, -4, -35, -75, 89, 17, 124, -16, 105, -27, 5, 104, 110, 43, 40, -77, 22, -16, 23, 108, 43, 49, 65, 7, 69, 49, -8, 58, 46, -126, 114, -39, -8, -60, 122, 67, -3, -125, 23, -34, -17, 53, 62, -83, 63, 8, -4, 102, 41, -12, -46, -82, -49, -39, 97, 37, -78, -95, 34, 112, -60, 68, -38, -68, 125, 48, 76, -111, 104, -85, -16, -36, -122, -102, 96, 51, -102, 56, 121, -100, -10, 91, -35, 126, -20, 4, -100, -87, 35, -116, 102, 75, -102, -122, 40, 76, 3, -114, -55, 101, 42, 21, 116, 14, -115, -103, -66, -100, -46, -33, 1, -6, -72, -61, -37, 16, -116, 113, -94, -46, 20, 95, -22, 48, -95, -111, -118, 87, 59, 41, -71, -122, 9, 44, -41, 118, 20, -115, 20, 110, -13, 31, -121, 33, 91, 13, -7, 56, 17, -101, -38, 8, 11, -92, 125, 93, 77, 55, -118, -48, 21, 57, -48, -18, -7, 53, -59, -102, 58, 103, -106, -101, 94, 118, 90, -5, -62, -37, -8, 85, -54, -95, -80, -55, 34, 102, -114, 108, 115, -95, 47, 30, 29, 96, 61, 59, -110, 29, -81, 62, -93, -127, -116, -62, 35, -81, 31, 27, -32, -69, -56, 62, -66, 36, -105, -68, 84, 59, 34, -107, -87, 46, -122, 84, 83, -80, 5, -36, 3, -98, -89, -117, -57, -49, 30, 18, -114, -122, -42, 55, -9, -108, 115, -92, 28, -79, -27, 42, 118, -63, 11, 93, 34, -31, -36, 69, 71, 110, -47, 42, 24, -44, 108, -15, 51, -119, 113, -70, 15, -119, 106, 65, -112, 25, 24, -70, -43, -34, -95, -28, -36, -44, -92, -47, 21, 106, -48, 64, -128, -92, -29, 55, -121, -108, -99, -90, 61, -120, 0, 89, -83, 9, -72, 10, 127, -56, 24, -119, -78, -94, 90, 31, 80, -103, -51, 82, 79, 9, 81, 64, -45, -74, -119, -58, -24, 88, -107, -66, 78, 73, 63, 28, -97, -78, 36, -16, 50, -64, -21, 66, -33, -77, 106, -95, 62, 43, 40, -102, 22, -120, -18, 36, 113, -51, -12, 71, -74, 41, 104, -40, 11, 5, 40, 104, -77, -9, 67, 1, -111, 96, 9, 57, 65, 116, 95, 62, 3, 121, 67, -76, -88, -22, -83, 94, -60, -39, 127, -14, 119, 72, -10, -37, 114, 104, 27, 44, -77, -119, -38, -99, 13, -23, 3, -14, -83, 54, 119, -114, -54, 104, 127, -54, 52, 126, 99, -52, 106, -17, -24, 111, -15, 62, -71, -15, 54, -71, -9, -62, -25, -31, -47, -56, -54, 62, -120, -67, 7, -65, 53, 102, 61, -1, 106, -32, -84, -97, 10, -107, -109, -100, -109, 109, 72, 4, 111, -110, 13, 10, -98, 68, -37, 45, 110, 99, 86, -93, -88, 63, -16, -59, -120, -84, -59, -104, 103, 96, -17, 40, 59, 50, -118, 107, 35, 2, 25, 7, -30, -128, 14, 75, -114, -94, 115, 51, -51, 94, 108, -24, 97, -128, -89, 16, -73, 109, -82, 127, 68, 74, -22, -118, 5, 32, 18, -85, -62, 4, 97, 46, -74, 84, -7, -35, 81, 87, -33, -89, 68, 73, -19, -111, 6, 30, 0, -62, 48, -58, -42, -67, -128, -30, -95, -125, 126, -38, -44, -108, -122, 84, 50, 56, 88, -86, -21, -60, -90, 12, 38, -120, 2, 44, 48, 101, -56, -63, 111, -4, 41, 124, 4, -50, 63, -58, -94, 24, 58, -64, -54, 34, -31, -48, -31, -14, -51, 115, 92, -73, 30, 61, 16, 119, -5, 57, 125, 59, 63, 44, 81, -79, 106, -58, -75, -64, 99, 88, -9, -5, 106, -99, -36, 0, 20, 63, 52, 14, -25, -91, -65, 63, 14, 20, -21, -94, -9, -114, 58, -29, -90, -14, -70, 100, -96, 3, 34, 15, -54, -121, -12, 33, 49, 13, -12, -24, -43, 62, 121, 40, -119, -75, 119, -30, -78, -120, -76, -111, 44, -57, 6, 65, -16, -14, 22, 65, -42, -75, 121, 43, 100, -93, 24, -94, 68, 58, -42, 110, 13, 7, 70, -10, 124, 6, 20, 41, 2, 73, -57, 113, 105, 41, -84, 119, 46, -25, 37, 108, -38, 22, 46, 98, 40, 43, -100, -116, 64, 36, -60, -10, -106, 42, 44, 48, 126, -12, 39, -125, -108, -28, -18, 17, -4, 58, -113, -48, -60, -40, -38, 86, 37, -32, -48, 120, -88, -127, 104, -70, 109, -69, -89, -71, 52, -127, -94, 68, 26, 31, -43, 51, -76, -108, -117, -29, 57, 90, -63, -31, -108, -57, 65, 57, -71, 17, 108, 15, 94, 77, 19, -3, -113, -23, -15, -19, 99, 112, 14, 76, -91, 54, 123, 50, -62, 78, 43, -29, -125, 120, -108, -95, 79, 30, -68, -87, -62, 21, -124, 19, 52, 26, -120, 90, -37, -44, 127, -80, -111, -114, -75, -22, 83, 111, -118, -112, 93, 48, -43, -50, -100, 5, -48, -59, 17, -29, 64, -56, 58, 11, 69, -1, 49, 1, 85, -98, -66, 65, 39, -3, 59, -14, -74, -6, -110, 83, -89, -23, 92, 48, -27, -97, 27, 2, -86, -112, 52, 81, 0, -43, -71, 126, 53, 100, -11, -6, 42, -100, -60, -13, -51, 33, 88, -35, -78, 63, 24, -94, 65, 43, -79, 51, 39, 49, 109, -40, -26, -14, 24, -2, -108, 50, 4, -47, 105, -37, -47, -125, 99, -119, 17, 63, -99, -117, 54, 66, 111, -125, 52, -88, -5, -19, -39, 75, 46, -125, -22, -125, 41, 82, -93, -99, -105, -57, -106, -95, 51, -124, 49, 77, 115, 28, 53, 43, -108, -58, 8, -43, 78, 28, -19, -17, -103, 50, -46, 72, -35, -103, 18, -21, 24, 61, 13, 25, 113, 108, 116, 76, -83, -57, -92, -35, 72, 47, 79, -114, -118, 71, -108, -54, 50, -105, -118, -35, -94, 37, -99, 73, 29, -18, -63, 56, 58, -99, -83, -118, 98, -50, 35, -100, -11, -105, 1, -54, 81, 21, 55, 97, -111, 12, -17, 124, 104, -3, 32, 116, 26, 97, 98, -71, -17, 123, 24, -124, 113, -126, 39, -91, -35, 51, 38, -6, 94, 125, 106, 79, 15, -26, 3, -63, 115, -54, 21, -94, 38, -89, -55, -97, 85, -102, 7, 121, -81, 66, -3, 111, 114, 88, 78, -117, -22, -10, 29, -49, 89, 8, 108, 79, -113, -116, -83, 41, -50, -7, 91, 126, -48, -118, 16, 104, -81, -115, -13, 94, 22, 110, -118, -50, -75, -12, -99, 58, 8, 34, -15, -122, 70, -46, 15, -5, 109, 107, 100, -30, -101, 118, 95, 91, -121, 69, -33, 96, -107, 9, -69, 71, -45, -115, -5, -67, -41, 97, -69, -83, 119, -84, 23, -16, -15, 101, 57, -61, 112, -54, -74, 30, 84, -52, 9, 117, -88, -75, -74, 1, 2, 70, 87, -18, -128, -50, 11, 81, 124, -27, 95, 15, 83, -43, -32, 80, 32, -28, -31, -98, -110, -4, -102, 42, 125, 99, 124, 81, -113, 5, -117, 74, 60, 46, -59, 106, -32, 7, -30, -40, 94, 39, -42, 106, -14, 96, 99, -92, -10, -90, -76, -16, -2, -74, -24, -75, -26, 106, 12, -22, 119, 86, 97, -115, -118, 124, 115, -104, -112, -65, -7, 51, 20, 17, 116, 99, -43, 118, -64, -66, -55, -93, -42, -70, -88, -111, 3, -13, 62, -55, 12, -69, 85, -128, 90, 110, -20, -67, -86, 11, -119, -11, -82, 102, 11, 75, 24, -33, -54, 48, 38, -124, 51, 36, 63, 48, 36, 109, -125, 19, 45, -58, 79, 111, 55, -64, 46, 110, -128, -17, -61, 63, 114, -38, 34, -11, 9, 54, 90, -7, 96, 84, -45, -24, 79, 79, 118, -97, 70, -29, 1, 1, 93, -122, -63, 63, -107, -118, 89, -37, 0, -85, -4, -112, -15, -18, 86, -100, 123, 19, 11, 125, 122, 118, 65, 122, 102, -61, 119, -62, 70, -75, -59, 11, -84, -70, 49, -127, -24, 43, -14, 10, -81, 82, -8, 126, 6, -75, 45, -108, 41, -115, -66, 103, 15, -21, 69, 89, -74, 121, -1, -73, 80, -83, 95, -109, -106, 80, 70, -67, 33, -127, 116, -49, 106, 45, -23, -32, -118, -42, -77, 16, 105, 87, -22, -33, 112, 104, -69, -116, -34, -68, -79, -39, -124, -72, 30, 60, -32, 119, -92, 89, 77, -87, 5, -89, 73, -64, -93, 2, -81, 96, 127, 14, 12, 90, -41, 48, -45, -9, 124, 70, -72, 111, -66, -114, -86, -9, 61, -87, 105, -121, -38, 22, 6, 13, 67, 67, 45, -2, 127, 118, -66, 6, -105, -11, -3, -85, -15, 56, 101, -50, 54, -31, 98, -29, 55, -25, 100, 113, -4, 40, 110, -104, 78, -31, -100, -90, 12, 117, 101, 53, 55, -38, 111, 74, 96, -103, 37, -77, -100, -29, -46, -88, 48, 122, -84, -12, -19, -107, -47, -117, 45, -25, 78, 121, -48, -68, -111, -112, -115, -64, 86, -112, -46, -54, -53, -64, -124, 29, 6, 81, -98, 60, -6, 102, 13, 30, -104, -118, 14, 20, 0, 104, -86, -7, -77, -16, 68, 42, -67, -23, 33, 122, 91, 16, 42, 57, 41, 77, 55, 25, 90, 66, 119, -56, -67, 72, -92, -54, -83, -47, -13, 123, 39, 34, 39, 123, 40, 74, -99, -48, 11, 89, 15, 21, -8, -85, -16, -87, 20, 56, -15, -38, 18, 55, 24, 14, 96, 57, 84, 5, -111, 57, 13, 20, 105, 76, -102, -31, 98, 99, -62, 35, -17, 108, 65, -22, -28, 92, -17, -5, 122, -96, 109, -23, 79, -13, 56, -68, 114, -65, -50, -117, 58, 120, 127, -72, -127, 51, -54, 106, 118, -32, 47, -68, 2, 49, -52, 56, -114, -79, 54, -90, 124, -40, -40, -70, -37, -39, 79, -96, -85, 125, -40, -82, -120, -40, 107, 84, 44, 84, -5, -34, -12, -71, 11, -81, -64, 90, -19, -65, -126, 110, -6, 22, -8, 109, -112, -8, -98, -101, 90, 123, -48, 87, 120, 122, 80, 22, -24, -29, -101, 91, -26, -43, 29, 61, 110, 78, -20, 12, -35, -17, 109, -30, -73, -81, -103, -73, 71, -72, -73, 123, -40, -29, 77, 40, -7, 98, -5, -99, 101, 2, 95, -21, 28, 65, 94, 100, -94, 59, 84, 99, -40, 73, 47, -6, -48, 38, -28, -124, 19, 109, 79, 103, 46, -56, 99, 9, 26, 58, -87, -51, 64, 59, 49, 100, 85, 105, -43, -54, -68, -49, 82, -14, 57, -83, -70, -99 );
    signal scenario_output : scenario_type :=( -15, 2, -97, -23, -70, 1, -128, 29, 55, -42, -64, -127, -15, -66, 49, -31, -13, -16, -59, 37, 93, -48, 119, -6, 24, -128, 11, -128, 37, -21, 74, -75, -31, 7, -97, -38, -79, -79, 29, 127, 85, 127, -42, -43, -119, 18, 44, 29, 15, 127, 43, 49, -128, -16, -102, 23, -128, -38, -128, -97, -128, 36, -93, -33, -7, 70, -117, -71, 85, 32, 2, 114, 45, -90, -79, 13, -54, -90, -59, -103, -31, -128, -37, -114, -128, -58, -28, -7, -3, -15, 24, -63, 112, -64, 63, -108, 12, 5, 22, -58, 70, -39, 127, 54, 127, 16, 127, 17, 38, 127, 127, 127, 1, -128, -78, 107, 53, -128, -80, -27, -128, -65, 60, 127, 127, 50, 69, 0, 86, -85, -74, -92, 114, -75, 69, -73, 127, 127, 103, 79, 111, 86, -42, 47, 26, -15, 107, 29, -66, -64, -8, -60, -124, -128, -128, -23, 127, 57, -128, -121, -50, -101, -109, -101, 101, 15, 63, -48, 39, -49, -90, -18, -60, -103, -128, -96, 33, -54, -70, -128, -100, -109, 1, -124, 0, -27, 21, 22, 66, -76, -38, -73, -45, 103, -64, -81, -29, 73, -122, 28, -85, 127, 124, 54, 127, 102, 127, -74, 38, 3, -10, -103, -116, -85, -7, 127, 127, 87, 79, 34, 29, -73, 37, 60, -45, -23, 71, -128, -118, -15, 127, 127, -36, -97, -54, 18, -81, -95, -32, -49, -26, -26, 50, 118, -128, -80, -6, 45, -39, -22, -16, -70, -128, -66, -128, -49, -103, 127, -76, 59, 13, 127, 43, -96, -6, 44, -70, -18, -85, 8, 107, -22, 81, -13, 78, 21, 98, -7, 7, 117, 12, -2, 31, -44, -66, 68, 79, -7, -55, -64, 112, -3, 93, -128, 54, -123, -32, 2, 114, 50, 22, 49, 75, -128, -28, -42, 90, -64, -79, -6, -53, 17, -59, 6, -7, 29, -31, -17, -117, -128, -117, 96, 123, -15, -101, -127, 65, -102, 42, 127, 92, 44, -78, 101, -33, 102, 119, 68, -112, -95, -128, -116, -123, -27, -69, 76, -8, 116, 37, -60, -128, -70, -88, 127, 85, -6, -88, 12, 16, 113, -10, -111, -70, 114, 16, -128, -66, 57, -37, -64, -58, -21, 23, -58, 1, 58, -2, -37, -109, 6, -85, -65, -80, 109, -22, 127, -22, 78, -50, 95, -23, -128, -28, -95, -3, 21, 57, 64, -75, -59, -103, -31, -54, 12, -6, -58, -78, 26, 44, 60, -5, -8, 13, -79, -26, 88, 34, -55, 127, -102, 127, -49, 93, -128, -8, -128, -48, 23, 50, -70, -128, 5, 45, 12, -122, -97, 127, 68, 74, -107, -32, -74, 102, 127, 98, 111, 106, 74, 38, 1, 11, 112, -38, 90, 60, 42, 53, -124, -93, -103, -85, -116, 36, -73, 34, 127, 127, 22, -59, -91, 7, -107, -98, 1, -78, 53, -26, 34, -122, -65, 69, 85, -66, 96, 49, -91, -121, 68, -106, -128, -27, -75, 127, 13, 73, -6, 98, 127, -79, 97, 111, 127, 106, 45, -8, -55, -66, 47, 27, -128, -128, -128, -39, -57, -47, -128, 2, 23, 127, -96, -102, -57, 108, 42, 98, -17, -32, -6, 69, -75, -90, -47, 92, -33, -128, -90, -128, 11, -78, 124, 43, 47, -111, -114, -128, -63, -13, 102, 58, -85, -16, 106, -11, -128, -78, -42, 127, 102, -50, -109, -96, 93, 34, 55, -88, 7, 10, 23, 38, 11, -55, -34, -2, 66, -128, -28, 100, 17, -98, -88, 75, -128, 52, -74, 122, 45, -29, -8, 58, 78, 100, -21, -88, -128, -128, 33, -17, -44, -2, 127, 87, 29, 18, 59, -21, -128, -36, -128, -128, -38, -100, 50, -128, 39, -128, 127, -121, 86, -53, 127, 80, 59, -122, -2, -75, 32, -128, -128, -73, -113, -79, -128, 112, -45, 96, -55, 71, 76, 42, 97, 106, -47, -5, -116, -44, 31, 31, -74, 73, -128, -37, 1, 52, -128, -114, -57, 71, 111, 106, -92, -113, -92, -74, -128, 37, 60, 70, -90, 92, 21, -64, 11, 28, 76, -13, -128, -128, -48, -8, -78, 13, 127, -23, -63, -88, 101, -76, 101, -52, -28, -27, -63, -111, -117, -45, 60, -117, -117, -26, 11, 37, -79, -78, 50, -112, -128, -71, -128, 16, 18, -75, -63, 55, 127, -128, -123, -76, 70, -58, -75, -16, -118, -1, 36, 127, 127, 107, 58, 6, 96, 22, -18, 66, -1, -65, 26, 24, 70, 34, -91, 44, 15, -116, -59, 127, -28, 44, -90, 15, -107, -128, -114, -93, -16, 59, -17, 73, -34, 0, 37, -23, 127, 92, 70, 108, 5, -28, -21, 114, 36, -128, -45, 93, 42, -48, 75, -102, -107, -74, 59, 45, 123, 0, -73, -55, 74, 106, -26, -31, -122, -16, -116, -32, 6, 12, 39, 118, 18, -18, 5, 34, -2, 42, -76, -69, 21, -86, -96, -102, -128, -91, -128, -66, -128, -42, -24, -36, 6, 47, 127, -3, -1, -28, 32, 58, 48, -60, -6, -26, -71, 29, 57, -2, -123, -122, 122, -128, -71, -88, 85, 118, 16, 68, -49, -54, -128, -123, -128, -128, -79, -128, -128, -81, 106, -24, -11, -66, -34, 28, 78, 112, 112, 102, -100, 112, 58, 127, 18, -114, -37, -31, -5, -23, 127, 113, -68, -6, -26, 102, 1, 64, -118, 22, -45, 100, -75, -88, -64, 127, -128, 23, -128, 121, -52, 42, -37, 74, 17, -127, 17, 13, -114, -73, -79, 34, -15, 119, -128, -52, -102, -50, 28, 33, 127, -6, 118, 60, 127, 71, -101, -28, 97, 127, -59, 108, -28, 52, -8, 73, 127, 78, 112, 6, 49, 15, -128, -109, -128, 3, -128, 81, -128, -39, -114, 64, -128, -109, -64, -34, 16, 81, -42, 71, -3, 101, -38, -16, 27, -31, -24, -21, 97, 6, 127, 91, 107, -11, 101, -3, -33, -53, 15, 108, -27, -85, -92, 127, 127, -10, -48, -34, 102, 47, -109, -114, -128, 78, 27, 53, -10, -39, 127, -63, 21, -65, 15, -69, 28, -70, -34, -13, 122, -50, 73, -13, 29, 122, -107, -6, -64, 124, -63, 17, 42, 92, -114, 127, 7, 33, -85, 127, 43, 88, -128, 1, -6, 76, -55, -26, -124, -54, -37, -6, -103, 49, -75, -55, 16, 65, 22, 8, 68, -68, 37, -88, 92, 127, 127, -53, -38, -31, 42, 73, -127, 28, -128, -34, -117, 22, -2, 52, 32, -6, 22, -55, 60, 98, 2, 87, -26, -8, 95, 80, -128, -88, 10, -63, -128, -112, -27, -128, -118, -79, 78, 81, 13, -121, -1, 63, 127, -39, -28, -47, 79, 29, -128, -97, 70, 119, 70, 92, 98, 59, -79, 0, 127, -108, 28, -31, 116, 69, -7, -32, -16, -22, 28, 114, -128, -128, -59, -43, -128, -63, 87, 49, -28, 123, -102, 95, -119, -32, -122, -18, 68, 34, -128, -128, -128, -55, -91, 92, 80, 127, 80, -53, -121, -12, 95, -128, -68, 43, 127, 86, 88, 122, 60, 127, -31, 112, -113, -69, -128, -124, -117, -128, -128, -54, 92, 127, -93, 116, -18, 98, -128, -38, 70, 127, -15, 127, 38, 58, -63, 74, -109, -128, -66, 101, 23, -71, 31, 38, 127, 7, -128, -128, -98, -8, 66, -38, -103, 53, 74, -54, -100, 18, -10, 127, 64, -15, -96, 80, 100, 96, -117, 45, 91, -50, -86, -38, 48, -116, -38, 3, -80, -85, -114, 22, 127, 64, 71, -128, 76, 0, 80, -128, -116, -44, 86, -64, 0, -100, 127, -68, 48, -93, -36, -17, 97, 127, 127, 127, 127, 5, 127, 97, 103, -68, 27, 107, 86, 65, 68, -59, -43, 101, 69, 49, 49, -1, -33, 44, -36, 127, 34, -92, 6, 98, 53, 127, 122, -17, 0, -7, -13, 123, 52, 96, -65, 17, 38, 117, -64, 13, 127, 63, -27, -47, 107, 37, 127, 38, -121, -31, 15, -85, -2, 17, -8, -128, 63, -117, 33, -128, -101, -96, 127, 43, -128, -49, -12, 3, -68, 127, 106, 86, -45, 81, 7, -8, -24, -122, -22, 74, 127, 127, 127, 114, -11, 36, 49, 100, -118, -81, -78, 48, 118, 60, 65, 15, -34, 60, 101, 121, 111, -23, -33, 127, 101, 108, -128, -78, 10, -22, 1, -68, 66, -127, -34, 127, 91, 127, 15, 26, -111, -107, -128, -108, 1, -65, 10, 55, 22, -122, 78, 34, 116, -43, 10, 52, 118, 2, -1, -106, -6, -124, -58, 10, -22, -109, 127, 68, 86, -128, -13, 8, 90, 34, 109, 36, -58, 16, 96, -39, 69, 52, 60, 36, -2, 127, -24, 100, -71, 92, 123, -23, -52, -17, 90, -87, -118, -116, -109, 112, 17, 93, -117, 101, -34, 39, -66, 76, 122, 21, -75, -98, 34, 47, 127, 95, -6, 127, 52, -65, -107, 127, 87, -10, -12, 93, 47, -128, 2, 127, 64, -8, 123, 127, -78, 79, 0, 3, 15, -12, 127, 127, 80, 127, 6, 127, -71, 76, 53, 26, -66, -27, 37, -45, -100, -75, -85, 29, -96, -22, 127, 96, 127, 54, 38, -128, -64, -81, -114, -111, -58, 127, 2, -63, 3, 76, -32, -112, 127, 11, 54, -43, 117, 2, 127, 92, 49, 80, 103, 109, 34, 86, -91, -127, -59, -49, -32, 34, -13, 58, -7, 92, -98, 24, 55, 101, 95, 1, -31, 10, 101, 10, 93, 26, 75, 103, -27, -119, -98, -1, -49, 18, -128, -70, -31, 63, 127, 109, 113, -11, -85, -54, 86, -3, -11, -45, 52, -47, 80, -60, 28, 60, 127, 98, 34, -95, 33, 2, 3, -106, 113, -107, -23, 26, 127, 107, 45, -27, -52, -34, -122, -64, 44, -18, -128, -102, 64, -112, -128, -108, -42, 93, 43, 103, 127, 127, 63, -23, 39, 57, -91, 81, -95, 70, 116, 98, 37, -107, 1, -38, -58, -124, -117, 108, -5, -11, -109, -54, -122, -79, 7, -93, -128, -107, 11, 55, 31, -95, -24, -69, -95, 26, -101, -73, -58, 65, -47, 57, 127, 52, -59, -128, 36, -128, -128, -93, 58, -31, -36, 6, -64, -68, 24, -69, 86, -128, -49, -73, -10, -29, 29, 97, 5, 28, -128, -43, -128, 59, -128, 107, -75, 76, -100, -127, -53, 113, 59, -66, 21, 11, -116, -34, 17, 68, 49, -74, -28, -76, -119, 33, -74, 11, -16, 86, -75, -128, -24, -123, -66, -64, -15, -93, -107, 0, -71, 6, 11, 79, 38, -17, 127, -44, 127, 15, 5, 93, 85, 117, -101, -34, -109, -108, -75, 39, 78, -100, 8, 127, -22, -78, -64, 113, -128, -24, -76, -31, -85, 47, 24, -50, -86, -68, -128, 31, -123, -44, -70, 54, -103, 127, 95, 101, 63, 7, 17, -128, 102, -86, 10, -92, 29, -43, -53, 127, 111, -2, -58, 109, 43, -47, 68, 29, -42, 116, -81, -60, -48, 53, -81, -128, -45, -128, -97, -2, 37, 124, -43, 91, -128, 12, -28, 107, -45, -91, 90, 68, 48, -79, -49, 127, 96, 127, -128, 124, -109, 85, -113, -42, 11, 15, 0, -63, -74, -128, -63, -69, 88, 50, -76, -106, -95, -76, 127, 91, 5, -128, 26, -18, 5, -76, -37, 66, 31, 53, -128, -128, -124, -86, -108, -64, -64, 90, 43, 63, -8, -23, 127, 103, 117, -108, 38, 91, 81, -16, -128, -12, -18, 127, 123, 65, -59, 26, -28, 23, -80, 127, 5, 0, -95, 44, 90, 38, 21, -117, 21, -8, -128, -93, -127, 97, -16, 53, -112, -37, -34, 49, 78, -124, -97, -8, -88, -128, -65, 63, 16, -128, 13, 111, 117, -50, 0, 127, 112, -59, 48, 32, 0, 85, -69, -49, -103, -128, -32, 34, 22, 11, 127, 95, 8, -88, -43, -24, -90, 69, -128, -128, -81, 0, 34, -92, 73, -11, 47, -29, 127, 85, 78, -17, 107, 8, 2, -13, 86, -98, 28, 16, 37, 59, 52, 127, 75, 127, 60, 66, -10, 79, -73, 63, 3, 108, -29, 48, -81, 13, 74, 37, -11, 88, 123, 53, 13, -12, 85, 69, -128, -68, 55, 50, 44, 54, 124, -102, -55, -101, -52, 10, 58, 80, -119, -1, -103, -128, -128, 7, 37, 38, -47, 58, -128, 23, -50, 127, 2, 127, -128, 58, -114, 71, -128, -36, 92, 70, -74, -106, 47, -58, -119, -12, 32, 21, 53, 71, 127, -16, -28, -31, 127, -39, 112, -43, 127, 22, -13, -76, 97, 113, -121, -103, -6, 55, 0, -103, 79, 22, -93, -113, 90, -7, 43, 93, 117, 127, 15, 102, 1, 73, 127, 80, 73, 127, 64, -71, -57, 116, 96, -85, -29, -49, -64, -26, 1, 53, -54, -48, 54, 28, -128, -24, -48, 69, -121, -78, -57, 66, 111, -28, -50, 106, 112, 76, -10, -112, 92, 52, 127, 53, 127, 92, 22, -128, -48, 127, 113, -34, -28, 27, 79, -128, -2, -28, 64, -116, 127, 111, 11, -128, -34, -49, 16, -87, 100, 117, 23, -7, -128, 17, -96, 79, 127, 86, 64, -26, 118, -48, -58, -49, -7, -128, -128, -42, -27, 43, 21, 79, 68, 127, 106, 73, 95, 127, 74, -79, -81, -90, -128, -65, 93, -8, -127, -6, -75, -128, -36, 109, 81, -2, -101, -59, -65, -15, 92, 74, 8, -128, 1, 12, 85, 70, 112, 73, 33, -81, -76, -90, 63, 10, 127, 42, 81, -1, 33, 114, 90, 75, 127, 0, 7, -76, 87, 70, 11, -26, -71, 127, 36, 112, 122, 127, 114, -128, -81, 21, 80, 27, -76, -11, -5, -43, 100, -28, 18, -128, -37, -128, 34, 8, -32, -128, 78, -124, 70, -60, 127, -42, 32, -128, 21, 17, 17, -108, 68, 27, -38, -96, -128, 119, -111, 26, -124, 92, 103, -48, -119, 63, 107, 127, 8, 76, -128, -92, 50, -2, -48, -70, -59, -66, 122, 92, -3, -45, -63, -87, -28, 29, -116, -128, -91, -53, 78, -128, -66, -128, 29, -90, -48, -103, -80, -107, -86, -85, 78, -8, 48, 22, -1, 109, 100, -53, -55, -24, -32, -65, -16, -122, 101, -31, 32, -38, 6, -128, -85, 106, -76, -128, -42, -22, 43, 7, 43, -128, -16, 60, 76, -60, 86, -49, -48, 54, -80, -57, -128, -128, -18, -65, -114, -107, 39, 36, -32, -13, -12, -91, 79, 123, -85, -18, 32, 18, -128, -107, 96, 12, -22, -101, -64, -71, 59, 13, 33, 32, -17, 102, 112, 127, -1, 127, -57, 117, 8, 127, -128, 65, -122, 31, -49, 63, 127, -76, 74, -97, 101, 76, -5, -29, -12, 86, -23, -124, -88, -87, 91, -6, -36, -109, -16, -124, -5, -47, 10, 37, 127, 50, -28, 37, 97, 6, 39, -44, 71, -128, 92, 12, 75, -71, -113, -32, 7, 117, 86, -48, 63, -8, -128, -113, -90, -78, -60, 85, -21, -121, 7, 85, 60, -55, 127, -58, 127, -65, 106, 28, 39, -12, -27, 127, 127, 59, 123, 111, 127, 127, 127, 109, 18, -17, 29, -12, -38, -123, -58, -47, 127, -57, 37, -96, 11, 47, -37, -45, -98, 113, 64, 15, -109, 78, 15, 78, -53, -128, -128, -128, 36, 63, 113, -47, -128, 22, 117, 93, -73, 127, 78, 86, -12, 36, 16, -128, -90, -116, 57, -16, 92, 106, 96, 106, -96, -103, 24, 47, -32, -32, -22, -7, 87, -24, 59, -70, 27, -80, -11, 127, 86, 50, -7, -57, -54, -101, 114, 17, 45, 8, 44, -7, 86, -91, 70, -92, 127, 127, -42, -128, -76, -10, -57, -80, 12, -107, -44, -17, 2, -128, 10, 127, 86, -128, -127, 49, 98, -48, -2, 127, 47, -128, -102, 88, -15, 8, -2, 1, 23, -36, 108, 64, 103, -64, -54, -128, 49, -53, 96, -71, 81, 127, 37, 73, -45, 113, -23, -59, -22, 0, -93, 58, 23, 127, 24, 39, 10, 5, 31, 34, 127, -65, 32, -26, 121, -64, -128, -88, -54, -88, -128, -47, -74, 68, -44, 36, 53, 127, 116, 76, -52, 127, 17, 127, 13, -45, -128, 65, 116, -86, -116, -1, 114, 127, 79, 127, 15, 107, -128, 60, -39, 73, -112, 112, -8, 66, 44, -29, 39, -45, -43, 10, 68, 28, -124, -74, 48, 33, -85, -128, 26, -27, -2, -128, -34, 127, 54, -28, 127, 13, -42, -128, -47, -12, 88, -107, -78, 101, 91, -47, -53, -107, 37, -50, -128, -128, -47, 127, 122, -39, 60, 127, 127, 113, 100, 127, 102, -86, -29, 107, 17, -13, -128, -111, -39, -128, -65, -107, 116, -112, 116, -88, 63, 54, 87, -15, 53, 127, 10, 0, -50, 24, -78, -90, 116, -88, 16, 8, -50, -85, 127, 93, -128, -18, 95, 109, 7, 127, 26, 76, -13, 101, 0, -31, -28, -5, 121, 98, -64, 55, -26, 87, -36, -48, -91, -75, -33, -93, 53, 80, 42, -128, -13, 36, 122, -59, -102, -48, 127, 70, -65, 68, 88, -42, -98, 127, -22, -101, -69, 3, -43, -86, -10, 86, -39, 117, 45, 127, 16, 91, -80, 54, 97, -5, -88, 55, 97, 39, -81, 111, 53, -37, -86, 73, 39, 71, 47, 58, 48, 8, -28, -21, -22, 107, 127, 21, 127, -98, 102, -54, 59, 50, 123, 93, -128, -81, 127, 15, -109, -128, 50, -45, -102, -128, -124, 3, -128, -122, -57, 106, -74, -60, -121, 34, 27, 27, -65, 33, -71, 8, 98, -128, 10, -73, 118, 58, 71, -53, -70, -53, 79, -11, 16, 85, 7, 47, -79, 71, 37, -87, -49, -59, -81, 37, 127, 16, -73, -109, -22, -11, 38, -6, -17, 39, -127, -127, 127, 47, 127, -122, 2, -96, -1, 15, -86, 17, -37, 78, 107, 95, -45, 60, 48, -24, 1, -91, -38, -112, 7, 64, -128, -47, 38, -54, -54, 3, 63, -101, -117, -17, 33, 117, -66, -39, -73, 37, -39, -37, -64, -27, -5, 127, 117, 118, -55, 127, 127, 86, -17, 2, 119, 48, 6, -39, -23, 127, 78, 86, 22, 87, 127, -22, -26, -21, 109, 102, 24, -2, -107, -128, -113, -12, -128, -76, -42, 91, -81, 45, 127, 106, 123, -7, -78, -100, 68, 127, 101, 52, -64, -49, -68, 16, 124, -7, -12, -75, -91, 85, 28, 127, 10, 86, 127, 69, 75, -119, 75, -113, 44, 102, 109, -55, 12, 108, 63, -128, 38, -86, -128, -113, 5, 88, -96, 12, 0, 103, -49, -128, -124, -50, 91, -128, -8, 97, 127, 13, 127, -43, 100, -38, 96, 50, 66, 27, 5, -34, -52, -22, -15, -128, -128, -24, 57, -108, -128, 127, 118, 127, -106, -10, 1, 112, 26, -116, -122, -55, -50, -24, -58, -114, -106, -97, -50, 76, -24, -111, -114, -128, -128, -24, 60, -39, -71, 117, 29, 127, -69, -92, -124, 54, -38, 124, -52, -64, 44, 113, 8, 106, 121, 28, -26, -63, -53, -106, 57, -43, 127, 100, 127, -93, 70, -15, 127, 58, 127, -29, 76, -3, 127, 127, 103, 86, 68, 71, -31, 127, -32, 127, -32, 102, -128, 76, -58, 91, -79, -98, -47, -3, 119, -27, -101, 13, 87, 92, -68, -44, 127, 68, 63, -17, 127, -2, -80, -128, 78, -128, 116, -107, 70, -128, 17, -6, -54, -42, 127, 27, 88, 127, 108, -128, -63, 119, 127, -81, -103, 31, 65, 10, -54, 127, -65, 116, 26, 127, 95, -43, 0, 75, 127, 92, 22, 127, 47, -92, -128, 6, -60, -88, -92, -2, 13, 17, -60, -128, -95, -128, -128, -69, -90, -34, -58, 71, 87, 2, -97, 121, -65, 95, -109, 92, -6, 87, 12, 60, -22, -8, -58, 127, 60, 127, -11, -59, 38, 27, 80, -127, 73, -2, 71, 32, -11, 24, -45, 12, -37, 31, -36, 98, -8, 47, -128, 69, 113, 54, -37, 127, 59, -55, -37, 60, -24, -106, 59, -17, 75, 78, -44, 127, 127, 127, -7, -96, -22, 90, -43, 127, 74, 66, -27, 64, -37, -85, 119, -128, -111, -95, 33, -128, -112, 47, -10, -113, -108, -55, 28, -112, 47, -48, 60, -111, 60, 44, 127, 70, 55, -52, -11, -39, -128, -112, -122, -57, -43, -22, -65, -111, -113, -12, -128, 28, 43, 0, -31, 22, 75, 54, 18, 88, 88, 127, 111, 85, 127, 38, 127, -107, 127, -88, 109, 36, 127, 75, 36, -78, 100, -95, 33, -128, -57, -102, -76, -57, -10, -53, -86, 79, 44, -66, -92, 6, 127, 91, -128, -8, 92, 55, -116, 109, 31, -116, -123, -38, -27, -93, -128, -10, -128, 22, -59, 91, -128, 37, -37, 119, -57, 86, 127, 57, 44, -107, 18, -29, -29, -36, 64, -73, -21, 96, 39, 73, -96, -63, -81, 47, -88, -87, 102, 114, -88, 29, 109, 95, -128, -70, -42, -86, -128, -70, 127, 47, -116, -78, 127, 36, 32, -128, 127, -128, 91, -73, 90, -65, -128, -128, -121, 18, 92, -57, -50, -47, 44, -54, 36, 79, -128, -33, 69, 53, -97, 27, 2, -75, 34, -54, 47, -48, 11, 36, -86, 45, -54, 70, -32, 98, 118, 127, -8, 16, -69, 123, 81, 31, 78, 93, 98, 68, 65, 127, 127, 15, -10, -33, 111, -91, 17, -128, 87, -96, 39, -31, 74, 54, -34, 113, -122, 68, -75, 90, -97, 43, 66, 23, -3, 12, 106, -128, -81, -128, 37, -71, 127, -16, 116, 127, 31, -112, -79, 55, -98, -22, 18, -37, -2, 112, -121, 65, -88, 59, -15, 13, -45, 58, -29, -27, -128, 8, 113, 45, -93, -36, 108, -66, 28, 44, 76, -58, 87, 114, -21, -17, 10, -23, 117, -116, -37, -11, 26, -69, -101, -101, 6, 48, 87, -31, 102, 44, -96, -45, -38, 0, 127, 127, 52, 55, -17, -70, 78, -128, -66, -128, 55, -80, 97, -5, 23, 118, 42, -2, -128, -50, -91, 101, 44, -33, 2, 103, -34, 11, -60, 12, -12, 31, 127, 127, 116, 102, 123, 15, -86, -88, 28, -100, -44, 92, 36, -69, -128, -92, -128, -114, -128, 15, -123, 17, -69, 78, 112, 116, 122, -128, -60, -128, 127, -128, 113, -128, 113, -93, 87, -22, -73, 22, 96, 78, -116, -86, 107, -65, -128, -79, 103, 127, -107, -64, -53, 80, 27, 54, 127, 127, -1, 122, 116, 92, -7, 127, 64, 43, -128, -76, 21, 8, 16, -36, -76, -128, -128, -78, 91, 0, -70, -55, 58, -55, -45, -12, 18, 2, -3, 127, 103, -49, -101, -111, -12, -29, 76, -85, -54, -112, 127, 127, 0, -88, 44, 101, 79, -11, 23, -65, 116, 108, 101, -6, 101, 124, 58, 3, -88, 66, -103, 16, -22, -106, -16, 95, 107, 127, 127, 52, -13, -17, 119, -57, -66, 22, 93, 127, -119, -118, -47, 127, 39, -13, -121, 0, -53, 92, 54, -86, -64, -128, -39, -88, 97, 32, 102, -43, -122, 123, 0, 29, -128, -2, -117, 127, 80, -38, -116, -80, 127, -117, -128, -87, 49, -122, -85, -37, 54, 109, 121, -5, 68, 80, -6, -127, -122, 95, -10, 88, -81, 2, -70, -15, 54, 17, -43, -98, -90, 21, -112, 127, -58, 36, 0, 112, 127, -18, 73, 59, 68, -78, -93, 49, -13, -45, -38, -128, -80, -75, -36, -128, -100, 31, 13, -102, -114, -128, 91, 12, 23, -128, -54, 21, 38, 11, -75, 64, -123, -8, -128, -79, 23, -50, -18, -68, 122, -80, 47, 103, 78, -65, -128, -79, -60, -101, -79, 63, 42, 103, -81, -50, -13, 87, -48, -15, 69, -28, -37, -111, 22, -87, -128, -68, -22, 18, -87, 70, 127, 127, 17, -52, 109, 127, 116, 119, 68, 88, 74, 127, 74, 127, 48, 127, 123, 1, 8, 50, 69, 50, 24, 117, 0, 123, -75, -11, -70, 91, 118, 5, 48, -65, 90, -79, -6, 124, -48, -88, -116, -2, -91, 127, -17, -107, -86, 81, 33, 5, 68, 80, -128, -55, -55, -27, 15, -2, 91, 48, 48, -24, 17, -81, -106, -100, 127, -96, 44, -17, -21, -36, -116, -18, -128, 68, -54, -24, -78, -124, 37, -101, 127, 24, -1, -76, 39, -71, 11, -53, -128, -39, -64, -128, -107, 116, 127, -11, -112, -128, 124, -128, -112, -128, 127, -128, -70, -93, 44, -28, 54, 13, -37, 96, 127, 57, 76, 15, 127, 103, 0, -128, -42, 21, 28, -102, 71, 127, 47, -128, -2, 81, -29, -128, -74, 11, 68, 23, 23, -128, 80, -16, 75, -80, 3, -119, 59, -28, 39, -44, -10, 127, 102, 127, -128, 80, -121, -18, -55, -18, 109, -44, 98, -123, -116, -17, 75, 59, -113, -69, 63, 76, 118, 127, 42, 26, -88, -16, -128, 42, 117, -116, -128, -127, 64, -37, -27, -106, -28, -33, 60, 124, -54, 24, -28, 108, 121, 76, -75, -22, 48, 55, -97, -103, -128, 66, 26, 48, -91, -5, -128, -93, -88, -18, -79, 50, -12, -48, 112, -36, -70, -71, 58, 127, 16, 5, -128, -117, -106, -36, -34, 31, -7, -1, -93, 29, -71, 100, -128, 127, -29, 116, -21, 38, 64, 75, 127, 29, 127, 80, 22, -63, 1, 42, 63, 29, -121, -1, 42, 64, -74, 127, -74, -86, -111, -26, -87, 5, 38, 33, -101, 121, 96, 106, -128, 32, -36, 29, -87, 86, 34, -128, -76, 106, 23, -36, -90, 27, -60, 7, -27, 86, -73, -128, -71, -43, -57, -81, 11, -64, -60, 36, -52, 85, -18, 127, 7, 118, -95, -81, -69, 69, 86, 50, 48, -16, 24, -63, 69, -68, -98, 122, 96, -73, -128, -57, -21, 87, -42, 127, -23, 107, -96, 127, 78, 24, -52, -24, -18, -122, 68, -58, 127, 117, -2, -38, -57, 12, 21, 45, -58, -45, -111, 34, -91, 114, 93, 127, 116, 37, 55, -42, -13, -12, 127, 66, 75, 65, 109, 7, 109, -21, 116, -1, 127, -47, 52, -15, 64, 3, 44, -16, -21, 127, 127, 127, 127, 114, 127, 127, 117, -3, 127, 54, 42, -87, -22, 52, 3, 3, -18, -24, -29, -26, -27, 127, 66, 127, 119, -24, 0, -15, 33, -73, 127, 127, 32, -50, 57, 6, -88, -128, 127, 6, 96, -128, 17, 23, 0, -128, -52, -47, 66, 12, 127, 48, -53, -128, -52, -5, -15, -52, 55, -3, 117, 117, -33, -113, -92, -21, -3, 8, -18, -64, -34, -64, 22, 127, 123, -18, -76, -128, -128, -87, 26, 31, -39, -121, -128, -79, 95, 93, -2, 74, 5, 124, 48, 42, -48, 22, 58, 123, 127, 22, -21, -7, 23, -121, -128, 39, -6, 29, -90, 65, 90, -5, -69, 32, 113, -63, -117, 88, 124, 3, -128, -70, 37, 17, -2, 13, 127, 71, 34, -53, 22, -128, -22, 107, 73, 55, 42, -54, -24, -1, -58, -48, 127, -33, 52, 69, 28, -42, 16, 58, -26, 127, 86, -8, 28, 127, 33, -8, -63, 93, 64, -23, -17, -21, 45, -124, 6, 70, -54, -17, 96, 28, -100, -128, -128, -22, -18, 47, -31, 112, 24, -85, -18, -128, -55, -71, 42, -78, 127, 121, 116, -17, 52, 39, 113, 117, -31, 54, 15, -5, -121, -108, 80, 52, 112, 102, 127, 47, -74, -76, -44, 37, -57, 68, -88, -114, 24, 64, -29, -47, -119, 97, 98, 54, 6, 123, 127, 5, -74, -63, 2, 109, 73, 97, -128, -31, -106, 45, -15, -13, -2, 76, 16, 127, 16, 102, -102, 5, 2, 50, -23, -121, -114, -16, -69, -8, -53, -39, 32, 109, 86, -59, 8, -60, 22, 59, 57, 21, 127, -118, 39, 0, 127, 106, -112, 127, 90, 119, -49, 63, -128, -112, -119, 8, 39, 86, 13, -68, 85, -71, 124, 34, 127, 127, 87, -39, 74, 47, 58, -128, 127, -93, 74, -34, -17, 34, -128, 21, -73, 5, -128, 48, -96, -13, -42, -128, -80, -128, -26, -63, 55, -68, 24, -128, 55, -53, -13, -107, 10, -38, 45, 52, 127, 88, 112, -5, 44, 68, 1, -103, -54, 118, 116, 63, -73, -128, -74, -92, 68, -112, -65, -23, -106, -128, -128, -63, 16, -90, -101, -59, 23, -43, -6, 127, 11, 75, 103, 29, 96, -15, 127, 32, 39, 37, -3, -28, 65, 127, 64, 91, 74, 50, -64, 17, 45, 11, 85, 59, 53, 55, 63, 102, 79, -101, -88, -27, -128, 100, -86, 80, -10, 85, 92, 36, 100, 118, 73, -91, -128, -52, 78, 73, -65, -52, 92, -8, 113, -66, -42, 44, 81, 42, -86, -73, 71, 88, -123, -107, -116, 127, 87, 127, -108, 10, -116, 42, -38, 17, -53, -128, -124, -22, -66, -34, 55, -16, 92, 85, -3, 0, -103, -24, -128, 10, 28, 24, -90, -38, -22, 22, 81, -5, 11, -127, -36, -128, 75, -71, 92, 37, 74, 85, -42, -43, -111, 44, -34, -32, 5, 27, 96, 18, -6, -95, -128, -37, -27, 69, -85, 121, 101, 6, -128, -97, 12, 96, -123, -76, -124, -79, -128, 12, -85, -90, -36, 103, 85, 34, -12, -29, 122, 116, 127, 97, 98, 23, -73, -3, -128, -128, -58, -60, -12, 2, 127, 81, -32, -128, 127, 34, 109, 2, 123, 122, 6, 63, 116, 37, 7, -98, 0, 45, -128, 13, -27, 95, -48, 38, 90, -36, 44, 7, 127, 91, 27, 80, 75, 1, 32, 127, 15, -54, -59, 29, -98, -10, 127, -43, -32, -69, 98, -39, 107, 92, 90, -128, -111, -108, -13, -3, -74, 50, 38, 79, -29, -128, -121, 52, -66, 3, -128, 101, -63, -21, -17, 39, 124, 74, 106, 43, 47, -32, 78, -38, 127, -128, -57, -81, 88, 90, -128, -39, -2, -39, -128, -52, -63, 86, -69, -92, -45, 76, -57, -122, 63, -12, -31, -85, 54, 22, -29, 2, 119, 109, -33, -31, 24, 114, -69, -44, -74, 45, 93, 1, 12, 66, 127, 87, 50, -122, 18, 86, -128, -23, 3, 118, -57, 97, -53, 76, -24, 119, -95, 63, -97, 127, 38, -81, -54, 98, -36, -79, -38, -21, 70, 27, -128, -112, -81, -114, 74, -52, 48, 23, 111, 24, 50, 92, 108, 48, -16, -106, -28, -76, 12, -53, -98, 73, 113, 91, -98, 12, -10, 59, 127, 78, 15, -98, 15, -63, 70, -7, -76, -128, -88, 122, 127, 52, 97, 118, 74, 102, 88, -52, -78, -127, -59, -29, 93, -26, 21, 17, -1, 81, -50, 107, 107, -63, 29, -38, 7, -18, 93, 32, 127, -22, 18, -22, 44, -16, -106, -64, 43, -12, 16, 3, 90, -45, -71, 48, 97, 119, -60, -58, 6, 112, 127, 63, -42, -33, 39, 31, -34, 91, 92, -85, 36, -87, 107, 57, -47, 3, 69, -53, 59, 65, -116, 36, 1, -28, -124, 45, -66, 127, 50, -6, 92, 33, 127, -52, 92, -54, 127, -28, 37, -53, 95, 0, 78, 31, 31, 13, -8, -54, 21, -53, -24, 18, -12, 73, -92, -47, 88, 8, 85, -81, 87, 92, 44, 15, 57, -12, -17, 63, 60, -59, 1, -37, -91, 2, -48, 42, 54, -74, -44, -6, -38, 68, 93, 127, -34, 127, -52, 127, -96, -86, -29, 93, 16, -33, 127, 90, -54, -85, 87, 52, -29, -113, -54, 23, -128, -128, -128, -118, -127, -128, -112, 7, 74, -128, -100, -2, 93, -88, -50, -28, -101, 18, -71, -43, -123, 7, -52, -128, -121, -49, 75, -38, -97, -13, -128, -103, 123, 127, -18, -69, -86, 60, 96, 68, 6, -65, 127, -17, -55, 26, 78, -11, -38, 81, -108, -79, 33, -59, 10, -48, 23, -95, -2, 50, -116, -68, 63, 95, 5, -32, 17, -111, -10, 24, 127, 17, -86, 23, 98, -128, -119, -108, 6, -128, -31, -79, 127, -42, 85, -12, 119, 8, 85, -128, -22, 127, 124, -37, 127, 127, 103, 32, 57, 29, 16, -128, 16, 29, 80, 36, -91, 85, -53, 13, -66, -44, 31, -96, 22, 18, 116, -23, -34, -121, -55, -114, -13, -29, -2, -43, 87, -111, -87, -87, 63, 57, -93, -15, 26, -70, -123, -13, -17, 7, -73, -128, -91, -50, 50, -116, 79, 0, 43, -116, 97, 21, 87, 2, -121, -57, -128, 21, 45, 13, -91, 70, 118, 127, 7, -128, -42, 64, -69, -106, 66, -57, 88, -36, 86, -128, -128, -128, 1, -55, -32, -33, 3, 127, 112, 64, -29, -78, 96, -50, 8, -122, -68, 127, 73, 8, -128, 10, 7, 124, -5, 108, -128, -76, -11, 127, 76, -85, 127, 106, 53, -63, 127, 29, 48, 5, 113, 11, -107, -48, -15, 65, 33, 47, 88, -17, 66, 64, 8, -44, 102, -90, -128, -76, -60, 127, -5, 69, -128, 86, 8, -33, -79, -124, 74, 23, -5, -117, -1, 54, -68, -12, 127, 127, 33, -122, -87, 90, -116, -12, 5, 127, 93, 3, -63, 33, -128, -95, -48, 23, -128, 29, -55, 34, 10, 102, 114, -24, -17, -128, -75, 17, 127, 97, 114, 55, 43, 127, 127, 114, -68, -98, 48, 71, 85, 127, 48, -71, -128, 108, 5, 23, -116, -109, 119, 54, 96, -64, 91, -16, -52, -109, 75, 16, 60, 127, 0, 118, -96, -3, 36, 29, -22, -93, -103, -36, -65, 8, -119, -55, 10, -71, -10, -123, -128, -109, -26, -5, -55, -39, -85, -26, -15, -80, -75, -13, 29, 50, 101, 101, -16, -11, 52, -73, 12, 22, 44, -73, -37, 109, 60, -128, -50, 127, 123, 78, -2, 127, -13, 28, -70, 127, 17, -5, 2, 91, -50, 27, 11, 79, 63, -1, 29, 53, -55, -69, 27, -1, 57, -42, 70, 75, -95, 47, 118, 96, 57, 22, 27, -95, 119, -107, 43, -49, 34, -81, 17, -116, -64, -114, -23, 27, -118, -102, 127, 54, 11, -24, 108, 39, 59, -21, -10, -55, 0, 10, 8, -57, 49, -124, 0, -71, 39, -66, 78, 23, 78, 127, 117, 109, -44, 37, 127, 10, 21, 1, 91, -118, -65, -79, 88, 39, -38, 85, 54, -24, -108, -86, -85, -53, 29, -32, -3, 87, -80, -28, -128, 90, 65, 54, -54, 59, 101, -13, -24, 127, -7, -23, -63, 0, 69, -107, 127, -38, 63, 12, 66, 73, 29, 127, 6, 102, 5, 127, 39, 34, 6, 28, -78, -93, -100, -44, 79, 22, -68, -6, 63, -81, -43, 65, 1, -39, -75, -76, -26, -98, 1, 86, -128, -27, -6, 85, -96, -127, -128, -111, -101, -44, -103, 111, 28, -11, -102, 91, 32, 1, 6, 90, -36, -11, -93, -31, -7, 15, 31, 65, 26, 57, -23, -93, -3, -47, 127, 70, 127, -86, 106, 127, 127, 81, -3, 124, 127, 17, 73, -21, 107, 60, -119, 42, 29, -80, -85, 17, -128, -128, -78, 111, -81, -109, -90, 127, 118, 86, 0, -48, -79, -106, 36, 78, 2, -15, 45, 16, -26, 127, 108, 98, -79, 127, 28, 1, 17, 101, -92, 27, -10, 102, -127, -3, 127, 119, 95, -11, 86, -69, 16, -128, -128, -78, 60, -48, -7, -75, 92, 16, 127, 22, -109, -69, 71, -128, -90, -26, -37, 102, 34, 78, 43, 98, -31, -118, 121, 53, 107, 2, -57, -42, -52, 127, -27, 70, 103, 103, -71, -128, -102, -3, -13, 22, -128, -10, -54, 64, -85, -73, 0, -58, -66, 59, 11, -60, 0, -68, 119, 74, 90, -119, -74, 26, 8, 8, -36, 78, 63, -128, -23, -74, 22, 16, -70, 123, -113, 101, -108, -78, -86, 108, 127, 127, 29, -45, 55, 124, -58, -3, -111, 0, -21, 70, -116, -86, -93, 121, 103, 101, 15, -79, 63, 127, 98, 101, 31, 37, 127, 127, 106, 75, -57, -128, -2, 93, 55, -109, 127, 0, -52, -71, 127, 39, 96, 76, 11, -128, -113, -124, -76, -10, 23, 29, -128, 2, 26, 101, -63, 71, 11, 12, 44, 91, 90, -6, 42, -5, 85, 127, 127, 118, -36, -70, 127, 117, 38, -103, -85, 48, 92, 127, 86, -85, 74, 70, -54, -50, -128, 17, -71, 91, -75, -48, -128, -128, -91, 32, 127, 23, 8, -81, -76, 71, 10, -37, -128, -64, -127, -63, -114, 15, -102, 29, 108, 73, 39, -128, -66, 79, 90, -128, -101, -13, 109, -98, -109, -128, -52, 31, 63, 58, -76, 0, 39, 108, 101, -53, 18, -53, 95, -113, 13, -78, -24, -29, -121, -64, 127, 54, -73, -108, 31, 127, 52, -90, -117, -27, 75, -50, -114, 23, 66, 127, 0, 68, -66, 118, 76, 66, 98, 118, 80, 127, 15, 43, -109, 127, 59, 66, -21, 48, -87, -69, 0, 85, -119, -45, 87, 127, 127, 60, 65, -79, -29, -127, -128, 34, 92, 123, -32, 127, -70, -69, -100, -21, -7, 65, 116, -117, 12, -103, -54, -108, -128, -21, 39, 119, 26, 91, -12, 44, 7, -128, 58, -128, -48, -116, -45, -78, 69, -39, 22, -97, -87, -93, 64, 127, 27, 44, -103, 93, -69, -15, -23, -8, 114, -50, -22, 111, 127, 118, 81, -100, 45, 74, -32, 31, -38, 33, -98, -27, 79, 47, 113, 44, 127, 122, 70, 81, 103, 63, -1, -80, -11, -102, -128, -21, 23, 113, -90, 96, -102, 53, 16, -63, -2, 103, 63, -88, -2, -59, 34, -80, 33, -121, -71, 90, 127, 109, 57, -45, 24, -95, 7, -11, -128, -53, -106, 1, -64, 100, 55, -116, 18, -44, -26, 75, 44, 69, -76, 63, -121, -26, -128, -98, -117, -79, -13, 48, -26, 107, 27, 57, 118, 95, -90, -49, -17, 107, 21, 36, -57, -117, -100, -27, -39, 116, 116, 97, 3, -28, -76, 76, -66, -34, 127, 80, 127, -54, 74, -96, -47, 6, -80, 43, -98, -127, 36, 95, 5, -112, 53, 65, 17, -23, 127, 96, 75, 34, 65, 17, -15, 69, -128, 33, -45, 95, -76, -128, -103, -118, -97, -96, 22, 111, -26, -75, -128, 64, -44, 44, -49, 21, 79, -68, -10, 78, 127, -27, -63, -86, 102, 28, 118, 58, -1, -11, -1, 1, 91, 3, -91, -88, 34, -127, -128, -109, 80, 36, -3, 15, 114, 11, 31, -69, 5, -95, -78, -86, 3, 127, 127, 8, -8, -16, 127, 86, -47, 57, 97, -7, 127, 101, 127, 73, 127, 127, 124, 127, 88, 127, 101, -23, -1, 50, 42, -128, 12, -97, 48, -48, 90, 64, 114, 127, 70, 26, -128, -18, 23, 54, 38, 127, 127, 96, 127, 64, 127, 58, 17, -53, -5, 68, 127, 121, -38, -17, 127, 85, -123, 98, 127, 96, -128, -113, 22, 118, 119, -76, 17, -113, 17, -64, 86, 127, 127, 58, -111, -128, -106, -76, -3, -64, -28, -103, 26, 79, -114, 6, 127, 74, -22, 93, 0, 127, 13, 114, -3, 127, 63, -75, -42, 50, -71, -119, 127, 5, -42, -24, 48, 127, 43, 87, 1, 32, 33, -26, 65, 47, -3, -96, -108, 24, -108, -95, -17, 23, -63, -24, 5, 74, 91, 12, 127, 127, 76, 39, -128, -36, -49, 81, -18, 8, -37, -47, 8, 127, 53, 111, 48, 127, 43, 97, -43, 27, -44, -70, -7, -92, 109, 127, 75, -68, 33, -15, -2, -97, 18, 28, 70, -34, 29, 127, 127, 47, -95, -17, -18, -16, 38, 102, 50, 127, -58, -59, -36, 107, -128, 87, -128, 34, -1, -17, -116, -73, 74, -127, -33, -11, 78, 70, 17, 88, -13, -128, -33, 44, 121, -87, 86, -124, 78, -128, 0, -128, 50, 29, 127, -98, 48, -60, 1, 34, 55, 109, 7, -113, -2, 98, 127, -6, 44, 22, 111, 117, -128, -65, -112, 123, -69, 55, -117, -66, -95, 59, 88, -75, -114, -100, -121, -26, -26, 92, -122, -6, -128, -114, 70, 33, 8, -108, 70, -70, 108, -37, 54, -128, -44, 79, 2, -95, -49, 118, -23, -32, 55, 127, 38, -27, -71, 81, 64, 18, 97, -53, -29, -128, 11, -8, 18, -128, -64, 74, 127, 127, 81, 127, 66, 69, -106, -34, 33, 27, -128, -57, 79, 127, 49, -76, -101, 34, 127, 114, 79, 100, 90, -42, -10, 48, -10, 2, -36, -38, 66, 127, 109, 127, 91, 86, 121, 107, -128, 7, 12, 108, -74, 65, -17, -31, -128, -55, -29, 118, -118, 58, 127, 58, -128, -128, -121, -1, -118, -78, -8, 113, 55, -96, 6, -10, -63, 68, -8, -117, -96, 5, 78, 15, -36, 38, -24, -59, -100, -59, -128, -65, -68, -128, -38, 68, 37, -17, -128, -112, -78, 111, -93, -17, -18, 53, -13, -33, -16, 127, 23, 127, 22, 70, 113, 24, -128, -81, 23, 127, 127, 57, -109, 75, 121, 73, 15, -128, -52, -50, 87, 0, 127, 107, 38, -124, 118, 15, 93, -45, 109, 127, 36, 17, -128, 18, -33, 88, -74, 5, 97, 63, -8, -31, 59, -70, 5, 10, -128, -11, -50, 127, 27, 127, 58, 32, 127, 127, 79, -119, -52, 54, 58, 108, 54, -85, -26, -18, 47, -118, -28, 101, 88, 47, 127, 80, 8, -128, -24, 93, 122, 5, 54, -49, -50, 42, 65, 63, 108, 3, -65, -128, 54, -76, 3, -76, 27, 97, -74, 123, 97, -81, -123, -3, 68, -2, -55, -43, 81, 127, 0, 5, -107, 86, -128, -107, -128, 36, -57, 127, 63, 81, 95, 36, -128, -59, -23, 47, -22, -44, 58, 11, 76, -102, -2, 49, 111, 81, -88, -128, -71, 2, 74, -37, 21, 28, 73, -74, 127, 13, 122, -18, 127, 76, 59, 54, -3, 6, -108, 29, 50, -102, -66, 93, 127, 96, 45, -32, 24, 0, 57, 127, -124, -13, -97, 53, -128, -42, 32, 31, -55, 27, 27, 65, 38, -54, -59, -63, 100, -79, 10, -107, -87, 86, 24, -128, -81, 88, -109, -70, 66, -15, -36, 13, 78, -39, 13, 113, -45, -55, -128, 3, 0, 103, 68, 127, 107, 127, 53, 101, -85, -85, 2, 78, 55, -17, 127, 21, 10, 50, 86, 15, -26, -13, -128, -107, 50, 63, -93, -88, -101, -74, 100, 97, 123, 10, 81, 78, 116, 24, -54, -68, 34, -39, 127, 113, 0, 15, -78, 6, -7, 112, -103, 127, 26, 57, -128, -90, -48, 58, 69, -16, 57, -21, -128, -127, -128, -66, -15, 123, 108, -119, -102, -75, 39, -106, 16, 50, 12, -8, 122, 79, -101, 127, 76, 5, -90, 109, 48, -1, -3, 64, -22, -38, -116, -44, 127, 37, 92, 10, 90, -73, 64, 15, 59, -68, -52, -87, 127, -103, 31, -87, 127, 18, 103, -65, 59, 38, -7, -31, 23, 75, -98, -128, -64, -128, -21, -118, 96, -15, 65, -55, -98, 106, 42, -117, -78, -1, -128, -128, -128, -71, -7, 26, -33, -111, 39, 81, 103, -128, 57, 100, 53, -44, -12, 15, -60, 127, -47, -13, 43, 116, 127, 102, 81, 127, 21, 50, -107, 66, -86, 111, -21, -16, -59, 54, -47, 127, 60, -90, 55, 114, 6, -45, -8, 96, 23, -87, -6, -128, -101, -52, 80, -66, 127, -12, 24, -24, 97, 7, -86, -113, -128, -112, -112, -78, 16, 12, 114, 71, 53, -128, -44, -11, 93, 60, 44, -45, 37, 73, -10, -6, -28, 91, -98, 79, -11, -69, -42, -24, 80, 98, 17, 127, 47, 69, 16, 121, 127, 16, -91, 75, 123, 37, -75, -73, 127, -69, 74, -68, 65, -73, -28, -23, 55, -59, -26, -128, -128, -112, -15, 113, -48, -10, -36, 93, -24, 60, 28, -128, -55, 103, 103, 58, 95, 75, -70, -27, 127, 97, 26, 108, 106, -55, 27, -109, 66, -38, 93, 6, -58, 63, 3, 66, -81, -128, 42, 5, 81, -107, 66, -34, 103, -52, 127, 66, 45, -31, 117, -3, -128, -7, 5, -33, -128, 112, 29, 38, -111, 75, 88, 127, -27, 53, -49, 103, -64, 101, 57, -18, 32, -128, -119, -32, -45, -66, -11, -75, -58, 0, -60, -78, -49, 24, 3, 6, 127, 49, 42, -80, 11, 2, 118, -128, -43, -52, 75, 23, 29, 74, -7, 34, 0, 44, 60, -128, -8, -27, -81, 0, 48, -38, -128, -32, 37, -13, -90, 96, 76, 116, -128, 76, -34, 5, -60, -128, -58, -47, -44, -109, -128, -1, -18, 127, 98, 112, 1, 33, -5, -76, -74, -128, 17, -79, 96, 127, 68, 52, -3, 44, -96, -123, 127, 79, 80, -43, -66, 118, 13, 127, -86, -11, -92, 90, -103, -38, -128, -81, -60, 39, -7, 38, 76, -73, -86, 76, 27, 47, 127, 85, 123, 45, -6, 26, -88, -65, 28, 71, 47, -128, -59, -60, 65, -69, -128, -42, -21, 78, -31, -95, -15, 6, -34, 43, 127, 16, 38, 96, 127, 97, 127, 98, -73, -128, -54, -85, 1, -50, 127, 48, -113, 0, 5, -118, -22, 33, -74, -128, -70, 127, 95, -87, -103, 55, 0, -10, -128, -32, -111, 43, -128, -64, -68, -8, -101, -15, -55, -58, 1, -48, -42, -111, -65, 127, -11, 55, -6, 103, -128, 79, -63, -10, -90, 54, 49, -43, -70, -57, -71, 66, 75, 127, 100, -33, 101, 123, 16, -48, -57, -48, 127, -36, 43, -103, 102, -97, 118, 52, -58, -54, 48, -13, -122, -70, 107, -107, -80, -45, 18, 0, -3, -15, 29, 95, 48, 93, -16, 37, 88, 17, 18, -13, -66, -5, 106, 0, -70, -106, 12, -91, -23, -91, 112, -6, -86, -63, -65, 122, 16, 48, -39, -97, 24, -106, 100, 12, 108, 6, 85, -54, -74, -74, -33, 127, 18, 127, -71, 45, -63, 69, -1, 28, 36, -48, 8, -101, 92, 88, 21, -128, -95, -57, 127, 127, -54, 127, 27, 95, -48, -3, -92, 5, 13, 52, -128, 27, -128, 21, -128, -95, -80, -50, -58, -103, -64, -121, 114, -24, 96, -128, -27, -112, 36, -6, -69, -53, -24, -128, -128, -45, 7, -34, -93, 29, 12, -128, -96, 26, -47, -73, -6, 53, 93, -86, -59, -11, 127, 127, 75, -64, -112, 122, -90, 22, -64, 127, -64, -17, 65, 107, -43, 98, -70, 0, 3, 59, -108, 127, 118, 16, -73, 29, -109, -42, -18, 69, -128, -97, -52, -45, -27, 106, -10, 113, 73, 91, -78, -122, -111, -128, 75, -88, 16, -38, 69, 24, 21, 127, 112, 121, 76, 3, 23, 80, 73, 10, 28, -123, -128, -80, -45, 68, 34, 127, -3, -128, 74, 100, 27, -128, -88, -114, 31, -122, 127, -32, 109, -103, 93, -43, 86, 127, 85, 26, -43, 42, 36, 64, -116, -45, -54, -48, -116, 7, 127, -59, -59, -73, 127, 15, 112, 26, 127, -112, 8, -90, 96, 127, 102, 0, 22, 8, -49, -78, -49, -119, -88, 7, 44, -128, 18, -128, 107, -38, -10, -81, 42, 114, -128, -29, -128, 55, -114, 55, 5, 69, 38, 127, 32, 69, 26, 80, -119, 26, 32, -57, -91, -90, -128, -128, -60, 127, -16, -52, -3, 86, -128, -24, 31, 64, -128, -22, 127, 116, 121, 127, 12, -66, 127, 32, -128, -34, 87, 71, -128, -24, -96, 48, -114, -79, 116, 28, -128, -109, 85, -55, -109, -128, 15, -117, 57, -64, 71, -59, -101, -42, 127, 90, -66, -28, 54, 80, 16, 16, 18, -7, 85, 127, 127, 117, -2, -123, 43, -95, -71, -65, 18, -98, -57, 60, -32, 54, 37, -78, -42, -54, 1, -32, -128, -45, -6, 100, -91, -39, -1, 57, 96, -85, -43, 101, 42, 98, -128, -11, 3, 17, -79, -38, -63, 49, 127, 65, 52, 28, 86, 22, 103, -97, -28, -80, -103, -64, -21, 127, 38, 127, -18, 76, -97, -3, -128, -128, 34, 42, 47, -90, -68, -34, 22, 127, -106, 95, -95, 13, -128, -81, 18, 21, 45, 36, -34, -78, 73, -15, 107, -128, -128, -42, 24, 49, 53, -64, -128, -32, 116, 127, -75, 50, -29, 11, 13, -95, 43, 15, 78, 34, -16, 127, 18, -16, -49, -45, 2, 12, 114, -70, -36, -54, -116, -18, 11, 103, -96, 73, 106, 11, -33, 48, 29, 47, 32, 121, 0, 76, -128, 85, -128, -31, -107, 127, 17, -65, -106, 127, 64, 127, -33, 26, -58, 32, 58, 32, 86, -60, 5, 79, 29, 79, -28, -75, 111, 24, -8, -23, -106, 121, -128, 43, -26, 71, 24, 90, 93, -8, 74, -12, -80, 18, -70, 88, 90, 88, -43, 36, -38, -6, 95, 5, 15, 45, -108, 79, 127, 116, -5, 31, -8, -73, 13, -111, 7, -57, 114, -128, 22, -128, 75, -108, 0, -78, 31, 127, 106, 93, 127, 71, 65, 95, 96, -60, 11, 111, -5, -1, -28, -111, -75, -3, -33, -27, 111, 102, -12, 28, -127, 74, -97, -92, -103, -34, 127, 127, 12, 63, 44, 57, 36, 5, 127, 127, 127, 64, 108, 121, 63, -93, -66, 26, -3, 3, -81, 127, 24, 45, -128, 6, -78, -60, -28, -57, 0, 55, 127, -7, -128, -103, 76, 59, -87, -128, -128, -43, 15, 43, -52, 100, -6, -76, 10, 57, 102, -128, -69, 59, 71, -37, -106, -12, -119, 69, -21, -59, -128, -48, 17, 127, -34, 64, -64, 49, 1, -122, 8, 75, -24, -60, -58, -33, -123, -128, -96, 12, -93, -128, -128, -128, -97, -39, -128, -29, 85, 64, -128, -32, 52, -33, -31, 113, 123, 65, 127, 117, -37, 49, 81, 127, -7, 7, -10, 64, 103, -128, 13, -111, 2, -128, -58, 74, 0, -12, -8, -2, 98, -5, 24, -65, 31, 5, 127, 22, 57, -36, 107, -90, -128, -57, 8, -86, -124, -27, 24, 50, 47, -64, 21, 3, 76, 90, 0, -95, 12, 37, 49, 71, -103, 117, 2, -42, -2, 0, 127, -5, 80, -93, 73, -65, 122, -68, -76, 23, 127, -79, -18, -87, 58, 0, 127, 50, -31, -80, 127, 118, 86, 66, -113, -90, -93, -22, -90, 65, 127, 73, 49, -69, -106, -119, -128, -13, -122, 11, 85, 127, 81, 54, -50, 127, 87, 52, -92, 127, 127, 127, 22, 55, -23, 64, -75, -128, -33, -71, 10, -48, 108, 127, 123, -45, 53, 109, 86, -3, 97, 92, 55, -15, 68, 127, 21, 78, -111, 12, -29, 44, -3, 79, 92, 53, -68, -45, -114, 42, 69, 57, -6, 37, -123, 106, -11, -90, -128, -100, 0, -1, 36, 13, 121, -49, -106, -69, 29, -128, -96, -11, 48, -124, -58, 127, -76, -34, -60, 118, 48, 26, 26, 55, 85, -122, -32, 15, 127, 73, 64, -60, 85, -68, -128, -59, -13, -116, -78, 44, 26, -11, -1, 32, -128, -3, -106, 127, -37, 92, -113, 103, -97, 123, 66, 24, -39, 57, 76, 78, 127, 10, 42, -13, -49, -112, -128, 11, -116, 45, -118, 69, 93, 16, -128, -70, -5, 106, 27, 71, -102, 45, -128, 31, 44, 116, -128, 11, -43, 114, 63, 107, -1, -13, -87, -97, 127, 6, -93, -55, 36, -127, -65, 22, 63, -102, -3, -68, -76, -79, 111, -60, 68, 8, 127, 6, 26, -88, 31, 127, 87, -18, -107, -54, 122, 57, 127, -86, 47, -23, 76, -32, -16, -103, 124, 74, -5, -128, 8, 5, 97, -10, 42, 2, 78, 88, 59, -90, 21, -116, -86, -22, 21, 78, -55, -8, 65, 119, -13, 123, 87, 28, -128, -103, -128, 44, -87, 80, 15, 103, -81, 127, 68, -80, -106, -116, -54, -52, 63, 88, 127, -18, 32, -29, 127, 10, 79, 60, 92, 26, -18, 127, 103, 53, -2, -66, 88, 65, 76, 5, 88, -128, -95, 85, 66, -128, -128, -93, 43, -45, -128, -86, 42, 21, -100, 57, -128, 88, -63, 90, -60, -81, 81, 22, 29, 39, -37, -16, 15, 76, 15, 127, 127, 114, -21, 127, 22, -31, -27, 34, -109, 53, 53, 127, -60, 50, -60, 102, -47, 13, 68, 78, -128, 16, -71, 107, -113, -33, -58, 127, 68, -33, -5, 31, -114, -128, -98, -128, -10, -85, 3, -31, -80, 44, 48, 18, 127, -86, 75, -16, 118, 76, -21, 76, -33, -123, 16, 32, 68, -107, -101, 10, -24, 127, 24, -5, -52, 127, 91, 106, 101, 48, -34, 59, -11, -128, 57, 127, 57, -128, -93, 91, 71, -103, 59, 48, 124, -116, -7, -93, 43, -58, -128, -6, 63, -7, -73, -13, 37, -128, -90, -79, 127, 88, 73, -7, -54, -92, -55, 33, -106, -53, 91, -108, 0, -123, 127, -32, 70, -128, 34, -86, 97, -113, -81, -71, 127, -65, 78, -81, 127, 101, 27, -49, 100, 74, 2, 0, 49, 31, -36, -44, -128, -31, 96, -75, -79, 59, 65, 127, 37, 90, -114, 127, -8, 81, 32, 57, -48, -128, -42, -13, 12, -66, -128, 122, -21, 127, -119, 64, -128, 2, -86, 86, -112, 93, 63, 53, 45, 33, 12, -97, 60, 88, -32, 10, -108, -39, -128, 63, -96, 79, -24, -123, -91, -73, 127, -13, 73, -38, 127, 1, -128, -75, -13, -86, -64, 12, 58, -60, 127, -39, 95, -128, -68, -78, 127, 101, -119, 16, -124, 123, -54, 78, -128, 88, 73, -49, -128, -128, -81, -70, -34, -5, 66, 119, 3, 93, -78, -123, 91, 29, -44, -103, 53, 127, -2, -2, -16, 93, -71, 102, -124, -111, -128, -36, 28, 23, -128, -85, -2, -7, -93, -128, -60, -81, 122, -54, 66, 13, 73, 127, 31, 60, -66, 113, 127, 81, 127, 24, 93, 69, 23, -103, -128, -111, -22, -26, -70, -7, -38, -27, 88, 127, 127, 122, 50, -31, 100, 21, 127, -68, 127, -53, 127, -78, 109, -128, -5, -128, 47, -17, 87, -128, 107, 7, 58, -74, -34, 59, 57, 36, -119, -101, -55, 24, -93, 50, 36, -36, -12, 55, 34, 34, 32, -76, -128, -65, -52, 49, 44, 65, 24, -3, 78, -95, -60, 117, 10, 127, 57, 58, -127, -36, -108, 117, 81, 32, 10, 103, -34, 18, 27, -64, 6, 127, 127, 0, 127, 81, 64, -128, -60, -21, 59, 49, 127, 118, -21, -57, 127, 12, -71, -21, -11, -109, -91, 0, -128, -53, 97, 64, 18, 108, 81, -22, 8, -3, 75, 50, -18, -122, 44, 22, 127, -64, 95, -12, 92, 11, 88, 26, -119, -102, -17, 124, -24, -112, -80, 24, 10, 127, 93, -10, -38, -26, 108, -47, 49, 68, 0, 127, -37, 42, -81, 116, -128, 43, -1, 74, -128, -1, -102, -8, -128, -73, -58, -68, -128, -64, 92, 80, 18, 10, 127, 73, -69, -38, -81, -52, -33, 60, -128, 102, -65, -38, -71, 127, 49, -32, -128, -63, -121, 7, -53, 76, 109, 127, 127, -29, 123, 102, 10, -97, -73, -22, 73, -5, 127, -11, 88, -100, 76, -43, 127, -128, -7, -8, 96, -16, -92, -80, -38, 11, -13, -75, 113, -68, -128, -95, -34, -26, -123, -74, 92, 118, 95, -24, 50, 0, -10, -128, -47, 55, 75, -23, 15, 102, -128, 39, -127, -119, -128, -29, 6, 75, 17, 92, -50, 79, 127, 79, -13, 28, 60, 116, -70, 58, -15, 17, 21, 106, 107, -21, -48, -27, -38, -26, 109, 33, 22, 18, -13, -6, 53, 97, 79, 27, -22, -60, -7, 88, 50, 27, 43, 42, -24, 127, 127, 18, 79, -50, -28, -106, -128, -45, -127, 44, 21, 108, 17, 127, 88, 21, 91, 127, 44, -31, -31, -52, -52, -116, -29, 18, 42, 18, -3, -122, -123, 127, 127, 1, -69, 13, 88, -128, -48, -91, -8, 10, 93, -13, -50, 37, -37, 127, 32, 28, 22, 18, -45, -47, -7, -45, -21, -42, 124, -128, -71, 22, 127, 127, 86, 44, -8, 127, 127, 33, 85, 119, 85, -96, -21, 49, -5, 45, 90, 63, -106, -48, -100, -109, -50, -106, 50, 64, 122, 38, 127, 127, -33, 11, -43, 101, -73, 3, -54, -48, 106, -88, 95, -13, -33, -114, -64, -63, -47, -96, 37, -71, -63, 13, 38, -34, -128, -45, -58, 92, -118, -75, -15, -1, -80, 76, 127, 54, 75, -116, 27, -43, -128, -97, -98, 29, -107, -66, 63, -52, -39, 11, 70, 17, -128, -53, -16, 108, 7, 37, 92, 96, -117, -54, -128, 2, -71, -34, -128, -33, 10, 114, 44, -128, -6, 88, 59, -65, 0, 29, 45, -128, -44, -49, 127, 26, 48, 58, 127, 93, 42, 127, 33, 7, 36, 127, 42, -128, -58, 95, 5, -112, -60, 47, 42, 118, -49, -5, -22, 16, -34, 116, 127, 127, 91, 76, -79, 121, -128, -23, -43, -66, -64, -124, -17, -78, 47, 39, -117, -6, 127, 18, 64, 22, 109, -74, 8, -85, -16, 127, 98, 93, -50, 33, 0, 15, -12, 93, 127, 68, 69, -81, 23, -27, 69, 93, 75, -24, 123, 117, 47, -111, -85, 8, -38, -44, 103, 127, -55, 85, 28, 26, 76, -128, -111, -86, 33, -118, -119, -128, -64, 6, -48, -16, -81, -32, 49, 127, 32, -121, -80, -24, -128, -32, -8, 12, -49, 80, -12, 57, 42, -22, 50, -6, -95, 64, 65, -1, 70, 127, 127, 106, 81, 98, 52, 68, -128, 39, -52, 108, -128, 28, 15, 92, -87, -43, -100, -128, -37, -15, 124, 15, -6, 59, 34, 127, 127, -39, 2, 54, 127, -128, 123, -101, 79, -39, 81, 63, -68, 123, 45, -128, -36, -47, 127, -28, 80, -15, 127, 98, -31, 127, 8, 22, -43, 64, -70, -128, 31, -37, 111, -48, -11, -23, -10, 91, -66, 42, 24, 78, -91, -21, -39, 5, -80, 127, 106, 12, -28, 69, 60, -44, 59, -12, 95, 44, -117, -6, -128, -1, -42, -66, -53, 66, 23, 2, -71, 38, -98, 65, 44, 127, 81, 127, 0, 116, -78, 127, 113, 75, 96, 127, 114, -101, -52, -28, 117, -73, 17, -37, 117, 109, 23, 70, 0, 92, 127, 103, 34, -81, 52, -119, -70, -128, -78, -128, -37, -44, -102, -128, -81, -70, 73, 65, 52, 31, -2, 24, -52, -91, -6, 0, 43, 63, -70, -3, -16, 32, -128, -128, -128, -103, 10, 70, 8, -112, -63, -1, 100, -97, -128, -128, -128, 17, 85, 88, -103, -29, 34, 37, 65, 102, 127, 37, 127, -36, 117, -65, 88, 80, 58, -90, 108, -10, 24, 98, 127, 36, -102, 15, 87, -27, -36, 16, -60, -78, 112, 22, -96, -32, 107, 70, 109, 42, 45, -49, 49, -47, -114, 36, -73, 86, -74, -57, -38, -78, 57, 88, 60, -70, 69, -31, 92, -22, -93, 34, -18, -57, -128, 49, -128, 33, -109, 26, -65, -69, 43, -69, 45, -114, 58, -73, -13, 34, -34, 47, -23, 26, -27, -58, -37, -124, -6, -128, 74, -16, 122, -53, -33, -127, -26, -118, 42, -112, -128, -65, -39, 127, -44, 127, 34, 44, -95, 122, -13, 17, -80, 3, -47, 5, 127, 127, -66, -6, -21, 44, -75, 55, 92, -128, -12, -12, -3, 127, 90, 102, -114, 127, -32, -26, -73, -28, -36, -128, -107, -122, 81, -15, -10, -57, 127, -17, -71, -119, 32, 3, -79, 58, 93, 127, -73, 85, -111, 31, -27, -24, -64, -27, -107, -12, 88, 127, 33, -108, -108, 127, 44, 127, 57, -34, -13, -8, 127, -93, 33, -96, 3, 91, 44, 101, 15, -24, -66, -60, -44, -52, 59, -128, -119, -10, -85, 59, 64, 127, 64, 60, -60, 69, 55, 127, 111, 69, 44, -34, -37, -128, -65, -18, 106, -50, -64, -23, -97, -34, -98, -65, -32, 122, 118, 16, 100, 2, 79, -66, 42, -101, -93, -47, -48, 70, -47, 44, 122, -119, -13, -28, 37, -71, 54, 38, -48, 78, 97, 96, 13, -86, 127, 39, -79, -86, 108, 75, -10, -103, -128, 12, -85, 81, -66, -34, -128, -92, 10, -34, 1, 111, -128, -47, -108, 87, -128, -128, -71, 27, 127, 17, 39, -39, 118, 17, -36, -128, -87, -127, 127, -7, 114, -33, 11, -48, 0, -108, -68, 103, 91, -128, 3, 16, 69, -54, -54, 47, -37, 71, -98, 22, -47, -13, 55, -128, 97, -122, 100, -63, 60, 66, 48, 23, -95, 1, 81, -68, -91, 127, 98, 127, -63, 69, -93, 93, 127, 114, 80, 18, 15, -27, 0, 18, 16, -33, -128, -70, -78, -39, -44, 107, 70, 26, 127, -79, 93, 5, 100, 86, -58, 127, -13, 116, -116, 45, 78, 92, 43, 123, 21, -44, -59, 29, 73, 112, 64, -49, 127, 44, 78, -54, -21, 28, -60, 68, 44, 113, 59, -90, -64, 27, -39, -111, 47, 119, 118, 79, 95, 32, 98, 55, 21, 101, 117, 31, 127, -79, 49, 75, 109, 15, 112, 66, -107, -29, 32, 122, 45, 81, -38, -29, -128, -68, -55, -127, -91, 68, 81, -22, -17, -34, -34, 78, -6, -121, -81, 90, 13, -57, -128, 3, -53, -73, -64, -53, 54, 81, -31, -128, -36, 127, 55, -128, -128, 68, 22, 44, -128, -50, 21, -87, 0, 127, 73, -112, -97, 53, 127, 15, -2, 127, 71, -1, -69, -44, 127, 27, 55, 34, 119, 111, -43, 69, 95, 48, 122, 80, 31, -36, -6, 68, 113, 68, 38, -15, -5, -39, 68, -90, -112, 66, 18, 48, -50, -36, -3, -64, 116, 127, 127, -80, 6, -13, 127, -73, 31, -121, 74, 127, 59, -65, -60, -66, -27, 93, -24, -128, -80, -96, 2, -58, 3, 58, -127, 100, 54, 71, -79, 127, 127, 127, 90, 127, 64, 3, -53, 127, 76, -38, -128, -58, -47, 12, 6, 10, -27, 127, 75, 37, 7, 109, 63, 39, 81, 13, 98, -49, 55, -47, -111, 127, 75, 109, -55, 90, 32, 66, -70, 70, 34, -49, 29, -17, 85, -2, -33, -60, -57, 0, 117, -10, 85, 85, 36, -22, 13, -48, 39, -76, 118, 27, -78, -79, 53, -128, -92, -128, -5, -128, 50, -96, 0, 0, 118, -128, -128, 11, 127, 116, 2, 93, -108, -31, -28, 96, -128, -79, -53, -32, 3, 58, 106, -88, -75, 10, 97, -127, -109, 26, 44, 21, -111, 59, -52, 107, 127, 45, 60, -63, -78, 58, -68, -59, 21, 55, -18, -121, 16, -88, 127, 58, 127, -8, 91, 87, 49, -78, -128, 23, -128, 12, -66, 127, 12, 22, 127, 59, -81, -128, 8, -128, 0, -122, 111, -24, 127, -44, 70, -54, 0, 6, -45, -6, -88, -33, -71, 118, -49, -78, -32, 124, 57, -68, -26, -76, -52, -90, -97, -15, -21, 107, -102, 7, -23, 48, -39, 16, -128, -85, 96, 114, 7, 33, 127, 113, 127, 8, 47, -128, -76, -24, 118, 127, 60, -128, -53, 92, 58, 15, 111, 109, 127, 127, -114, -12, 59, 88, -103, 127, 103, 18, -121, 8, 7, 63, -58, -68, 92, -117, 13, -52, 127, -47, 91, -22, 127, 88, -127, 10, 58, 71, -76, 127, -124, -95, -87, 33, -88, -44, 65, -16, -13, -128, -28, 127, 101, -42, 18, 59, 101, -38, -2, 55, 80, -31, -16, -37, -31, 8, -55, -121, -16, 27, -79, -39, 3, 5, 7, 92, 108, 127, -37, -74, -12, 76, -68, -95, 127, 111, 44, -7, -91, 91, -87, 17, -17, 0, -78, -21, -44, -74, -128, -3, 71, 71, -54, 117, 107, -22, -1, 66, 76, -128, 127, -60, -13, -12, 117, 127, -13, 42, -108, -88, -124, -53, 101, 5, 45, -1, -5, -23, 118, 127, 127, 86, -54, -12, 102, 48, -48, 116, 75, 127, 39, 75, -96, -117, -75, 37, 60, 37, 49, 44, -128, -55, 76, -92, -119, -79, 32, 3, 28, -70, 95, -31, -17, 8, -24, -75, -85, -128, -81, -58, -103, -128, -113, 17, -88, 32, -24, -21, -43, 18, 88, -32, 70, 10, 79, 65, 127, 55, -28, -85, 27, 3, -34, -13, -90, 76, -79, 80, 22, -111, -91, 29, -75, -111, -91, -128, -86, -88, 27, -69, 119, 92, 5, 5, -37, 127, 80, 75, -49, -95, -128, 117, 95, 39, -55, -13, 111, -42, -32, -75, -47, 18, -128, -47, 43, 27, 10, 33, -39, -103, 3, 53, 52, 13, 55, -90, 0, 127, 54, 85, -73, 76, 100, 88, 107, 2, -102, -88, -58, -12, -33, -63, 2, 34, -32, -53, -112, -43, 27, 127, 81, 95, 97, 127, -31, 64, -74, -64, -128, -79, -103, 13, -128, -117, -1, -113, 76, 127, 26, -100, -66, 53, -114, -34, -28, -128, -106, -78, -29, 11, -107, 127, -32, 113, -18, 127, -121, 2, -100, 118, -90, -95, -15, 70, 24, -11, 127, 57, -71, -80, -16, -100, -124, -38, -85, -29, 98, 2, -3, -128, 24, -124, 85, -59, 27, 48, 123, 47, -78, -15, 109, 117, 127, 127, 119, 27, -28, 127, 127, 88, -13, 50, 42, -107, -116, 98, 33, 55, -26, 29, -66, -128, -11, -43, 87, -88, 0, 12, -49, 92, -93, 37, 91, 73, -128, -128, -95, -128, -128, -65, 5, 79, 29, 0, -21, -128, -128, -71, 86, -6, -42, -71, 88, 68, 71, -6, 58, -116, -11, -47, 6, -38, -102, 11, 42, -8, 29, 96, 69, 0, 27, -97, 29, -48, -37, 36, -22, -37, 8, 69, -128, -107, -128, -42, -128, 66, -122, -45, -128, -79, -13, 71, -128, -102, -68, 71, -52, 71, -81, 64, -128, -69, -57, 52, -90, -116, 7, 58, -28, 47, 76, -31, -122, -63, -8, 5, 34, 47, 32, -8, -128, 75, -101, -5, -117, -66, -66, 38, 27, -2, 127, -128, 111, -128, 2, -96, 13, -97, -74, 29, -64, -127, -93, 100, 98, 13, -13, 116, -64, -36, -128, -1, 29, 64, 21, 81, -10, 45, -27, 127, -75, 23, -128, -76, -37, -27, 68, 127, 55, -95, 6, 60, -128, -76, -78, 28, 106, 100, 93, 17, 127, -50, 100, -22, 76, -128, -97, 24, 45, -128, -44, -128, -128, -65, 42, 101, -128, 33, 26, 113, -10, 58, -60, 23, 10, 34, 127, 127, 32, 36, 50, 113, -128, -128, -66, 127, 96, 38, 127, 76, -36, -88, 127, -1, 34, -43, 106, -87, 95, -47, -71, -97, -128, -68, -100, -44, -23, -28, -80, 65, 52, -128, 6, 33, -58, -91, 103, 127, 127, 42, -54, -12, 10, 22, 55, 122, 73, -79, 7, -11, -8, -28, 59, -38, -127, -69, 68, 103, -107, -88, 6, 103, 66, -38, -65, -96, -34, 28, 7, -80, -18, -97, -86, -111, 22, 68, 107, -1, 38, -36, 107, 127, 113, 86, -43, -63, -86, 0, -1, -128, 8, 38, 98, 68, 66, -128, -100, -52, -34, -23, 65, 38, -63, 127, 38, 39, 78, -15, -106, -48, 65, -59, -3, -96, 127, 116, 118, -36, 91, -128, -106, -86, 100, -128, 34, 103, 74, -101, -69, 127, 29, 54, 27, 66, -73, 90, 87, -31, 68, 123, 15, -128, -91, -71, 42, -101, -23, -32, -128, -42, -101, 36, -59, 66, 6, 127, 93, -10, 15, 127, 121, 112, 127, 52, -21, -93, -52, -31, -8, -33, -128, -124, -52, 0, -45, -48, 42, 16, 22, -3, 127, 87, -86, 60, 43, -24, -49, 37, 21, -42, -11, -121, -128, 28, -87, 23, -60, -128, -2, 73, 86, -64, -92, -38, -16, 91, 107, -54, 10, 70, 47, 108, -42, 113, 5, 5, -37, -128, -128, -47, 103, 117, 16, 117, 102, 112, 78, 32, 57, -5, 37, 8, 6, 118, 127, -10, 108, -47, -8, -113, -90, 5, -65, 127, 90, -24, -78, 88, 34, 121, 96, 73, 65, 127, -128, -34, -73, 127, -6, 16, -58, 50, -38, -39, 121, 2, -31, 107, 127, 60, 39, -75, 53, -57, 81, -95, -123, -8, -87, -108, -112, -16, 127, 127, 79, -22, -108, 127, -34, -39, -31, 28, -103, -92, -69, -52, 10, 43, -28, -80, -74, 48, 44, 127, 80, 55, -13, 102, 28, 27, -127, -65, -76, -1, -63, 54, 118, -13, 65, -74, -73, 79, 103, -10, -16, -15, -29, -117, 127, 44, 86, -128, -74, -96, 127, 37, -8, -16, 127, 127, 127, 60, 70, 127, 127, 76, 37, -7, 127, 71, -118, -50, -33, -108, -26, -124, -53, -88, -69, -42, 69, 74, 11, 10, -49, 75, 71, -128, -36, 10, -64, -69, 127, -34, -7, -76, 15, -128, -54, -73, 60, -5, 74, 71, -16, -52, 114, 50, 49, -65, 2, -53, 12, 48, 91, -85, -36, -128, -36, -95, -45, -97, 127, 127, 8, -44, 57, 37, -39, 52, 127, 57, -66, -50, -87, -71, -24, -128, -114, -87, 48, -100, -63, -70, 127, 74, -86, 11, 87, -36, -96, 116, 118, 54, -71, 70, 7, 45, -39, 66, 13, -102, -78, 22, 86, 15, -24, 106, 7, 70, -47, 43, 37, 98, -6, -81, -74, -75, -17, 47, -10, 95, -10, 114, 75, 127, 71, 11, 26, 127, -57, -128, -86, 44, 36, -93, -79, 34, -128, -109, -119, -7, -53, 38, 12, 24, 92, -87, -52, 68, 127, 107, -86, -36, 32, 70, -44, -69, -65, 127, -128, -122, -128, 8, -128, -118, -128, -44, -7, 79, -111, 16, 106, 127, 81, 119, -23, 48, -128, 78, 127, 127, -98, -45, -76, 113, -64, -39, 74, 71, 127, -128, 43, -24, 87, -81, 0, -24, -66, -23, 17, -31, -5, 48, 119, 92, -59, 127, 1, 13, -1, 118, -68, 65, -7, 28, -17, 29, -109, -128, -128, -109, -22, 108, -66, -44, 97, 127, 98, 3, -88, 1, 6, 57, 3, -87, -109, -59, -10, 108, 118, -1, -74, -60, 81, 64, 36, -39, -45, -43, -103, -78, -42, 16, -101, -128, -113, -100, 34, 127, 127, 127, 127, 95, 127, 48, 127, 64, 37, -33, 111, 11, -97, -33, 95, 127, -60, -111, -23, 68, -74, -17, -45, 28, 15, -55, -116, 90, 85, 127, -49, 74, -108, -88, -128, -92, -128, -37, -128, -48, 17, 54, -92, -93, 57, -116, -128, -48, 75, -36, -114, -119, 92, 60, 69, -59, -128, -5, -48, 73, -127, 127, 96, 96, -111, 117, 101, 63, -32, -118, 108, 38, -66, 3, 2, 108, -73, 127, 117, -17, -74, 66, 117, -7, -87, -66, 13, -64, -1, 127, -80, 63, -128, -102, -70, -90, -33, -73, 119, 58, 50, 98, 127, 124, -8, 7, 0, 127, -34, 52, -90, 58, -58, -108, -38, 50, -17, 114, -63, 98, -36, 98, -27, 1, 127, 54, -7, 13, 107, 63, -26, -98, -98, -71, -66, -128, -113, 95, 27, 127, 68, 48, -128, 8, 58, -52, -116, 26, 101, -45, -128, -117, -128, -48, -128, -44, -79, 10, 15, 12, 127, -37, -87, -128, -60, -117, -23, 127, 127, 73, -74, -24, 63, 79, 80, -39, -26, -128, -60, 85, 0, -128, -11, 79, 23, -16, 127, 0, -48, -24, 57, -76, -119, -48, 127, 73, -73, -69, 93, -10, -64, 124, 43, 127, -73, 38, 28, 1, -128, -34, 7, 22, -29, 127, 117, 127, -28, 127, 87, 38, 16, 8, -128, -73, 127, 127, 114, 45, 73, 85, 78, -65, -111, -45, -118, -103, 29, -117, 36, -49, 127, 23, 127, 13, 28, 12, -66, -103, -88, 87, -114, 15, 88, 54, -50, -95, -128, -45, -123, -122, -128, 37, -23, -128, -128, -11, 81, -91, -55, 103, 118, 11, 13, 122, 57, 49, 98, -10, -23, -128, -79, -36, 127, 81, 47, -11, 42, -52, 85, 66, 65, -109, 29, 37, -18, -128, 90, -50, -7, -85, -6, 0, 37, 16, 127, 127, -2, -5, -102, 59, 76, 21, -66, -24, 8, 90, 91, -73, -128, -80, 75, 52, 54, -90, -8, -31, 127, 2, -128, -128, -79, 6, -128, -88, -69, 76, 118, -11, -81, -128, 57, -111, 70, -66, 93, -57, 81, 127, 127, 59, -8, 0, -3, -76, 117, 13, 49, -32, -42, 79, -91, -31, -121, -128, -64, -90, 127, 54, 27, 23, 91, 123, 36, 0, -16, 43, 127, 21, 127, 49, -57, -128, 95, 13, 49, -100, 95, -15, -2, -21, -116, 1, -85, -101, -91, -128, -96, -91, 6, -97, 64, -71, 38, -15, 0, -49, 114, 87, 10, 97, -88, -79, -15, 6, 81, 11, 127, 114, 68, 27, 127, 127, -5, 127, 11, 85, -59, 102, 22, -42, -2, 90, 78, -114, -107, 65, 28, -48, -128, 47, 28, 23, -55, -33, 97, -60, -121, -123, -128, 34, -58, 95, -91, -128, -97, 68, 2, -91, -43, 118, -27, -80, -58, 74, 92, 37, 112, -48, -16, -92, -69, 69, -109, 24, 75, -32, -60, 63, 103, 127, 86, 52, -114, -106, 112, -27, 53, -85, 100, -70, 113, -86, 85, 47, 31, 127, 127, 85, 16, 87, -13, -65, 63, 60, -75, -93, 15, -128, -128, -78, -10, -29, -53, -2, -42, -52, 60, -128, 93, -65, -21, -53, 70, -116, -128, 98, -23, 50, -55, 127, 127, 127, -64, -128, -24, 127, 87, -7, -128, -42, -128, -39, 5, -23, -128, -47, 43, 44, -39, 70, 0, -48, -74, 38, -101, -70, 39, -75, 38, 100, -24, -3, -47, 12, -43, 18, -128, -57, 118, -21, -1, 92, 80, -31, -119, -13, 43, 102, -128, 106, -60, 127, -63, 28, -55, -32, -1, -128, 127, -52, 60, -128, -69, -74, -128, -106, -128, 65, -97, 127, 7, 73, -128, -87, -93, 127, 87, 52, -113, 44, -23, 96, 69, -27, 91, 127, -106, -128, -48, 63, -10, -33, 59, -23, 127, 0, 93, 26, 7, -96, -128, 50, -128, -10, -27, 92, 12, -29, 45, 43, 103, -22, -3, 26, 127, -64, 74, -128, 102, -97, -7, -128, -63, -64, -107, -12, 93, 107, -8, -128, -128, -16, 48, 106, -6, 92, 23, 81, 127, 43, -48, -111, 91, -107, 127, 91, 65, -87, 70, 127, 86, 127, 54, -79, -122, -24, -96, 53, 87, 121, 75, -49, -34, -18, 87, -36, -71, 124, 18, -17, 47, -23, -128, -42, 123, 111, 17, 116, 127, 69, 121, -121, 43, -57, 98, 91, -1, 22, -50, -59, -128, 37, -87, -12, -100, 42, -59, 15, -86, -57, 118, 127, -16, -109, -128, 53, -124, 43, -109, 127, 11, -44, -128, 97, 68, 127, -57, 6, -75, 111, 127, 91, 34, 27, 95, -81, 16, 15, 71, -22, -87, 47, 108, -118, 16, -37, -1, -92, 101, -111, -128, -70, -11, 11, -50, 111, -43, -6, 5, -37, 85, -50, -87, -128, -90, 127, -48, -128, -69, 92, -23, -95, 80, 8, -26, 12, 127, -27, -21, -68, 63, -78, 39, -60, -128, -50, -81, 106, -32, 91, -38, -68, -88, -55, -27, 127, -52, 127, 21, 117, 92, 71, 86, 127, 76, -28, 54, 101, -71, 21, 127, 127, 127, 93, -47, -59, 87, 127, 7, -38, -22, 119, -128, -74, -101, 127, -2, 57, -28, 106, -53, -70, 24, 0, -1, -79, -128, -39, -39, 116, -22, -60, -49, 74, 68, -11, 109, 117, 109, -81, 27, 26, 92, -28, -23, -42, 32, 3, 80, 23, 52, 74, 127, 57, -53, -128, -100, -52, -128, -111, -48, -128, -128, -103, -124, -10, -47, 26, -88, -122, -113, -111, -17, 45, -128, -28, 37, 22, 95, 123, 65, -116, -64, -60, -47, 29, -27, -3, -36, -73, -92, 33, -69, -65, -70, 49, -48, 101, 121, 75, 7, 42, -37, -8, 0, 55, 64, 1, 122, 69, 48, 70, 57, 6, -95, -85, -1, -52, 34, 69, 55, 42, -29, 5, -13, -24, 96, 68, -76, -64, 101, 0, 48, 0, -57, -47, 78, 12, 23, -38, -7, -128, -37, 116, 48, -123, -116, -29, -88, -22, -128, -54, 53, 52, -90, 32, -24, -42, 127, 34, 127, -108, 127, -98, 57, -85, 39, 68, -128, -66, -73, 24, -66, 68, -59, 1, 22, -45, 63, 38, 127, 55, 6, -38, 121, 92, -111, -73, -128, 23, 127, 127, -74, 81, 78, 0, -18, -128, 76, -28, 112, -8, 58, -33, -47, 73, 122, 26, 91, 8, 44, 48, 44, 8, 31, 73, -50, 69, -68, -128, -16, 127, 106, 37, 52, -21, -118, -13, 12, -5, 57, -15, 49, 18, 27, -68, -28, -66, -71, 11, -15, 81, 127, 117, -32, -15, -15, 91, 48, -65, -47, -42, -128, 8, 102, 117, 37, 69, -48, -93, 86, -24, -95, 32, 11, 116, 127, 122, 127, 64, 100, 59, -11, 24, -98, 32, 127, 71, 45, -108, 34, 103, 114, 27, -128, -75, -127, 33, 73, 118, -128, -32, 58, 45, -53, -128, -32, -128, -38, 29, -69, -7, 6, 113, -59, 127, 127, 63, -80, 1, 118, 6, -22, -66, -13, -32, 29, 32, 90, 127, -15, 65, -92, 109, 45, 37, 17, -29, 127, 78, 39, -100, 13, -107, 53, 58, 127, 86, 15, -49, 102, 76, 59, 78, -118, -34, -24, 92, -74, -70, -101, -48, -128, -111, -106, 76, 87, 12, -128, 57, 36, 107, -27, 42, -63, -128, 113, -76, 49, -128, -8, 114, 102, -45, -7, -8, -33, 15, 18, 0, 55, -12, 0, -112, 127, -18, -90, -78, 127, 73, -10, -50, 21, -128, -128, -60, -66, 113, 49, -37, -128, -128, -47, -128, -73, -59, 66, -5, -32, 64, -128, -11, 11, 127, 127, 108, -79, 74, 127, 103, 114, -85, 127, 3, 49, -79, 50, -128, -86, -128, 95, -60, 55, -109, -32, 114, -111, -64, -1, 55, 28, -65, 29, 74, 36, 127, 118, 127, -36, 2, -71, 127, -85, -36, -70, 17, -68, -33, -34, 28, 37, -117, -102, 57, -124, -68, -85, 127, 23, 17, -101, 18, 16, -60, -2, -124, 127, 80, 127, -2, 118, -128, -98, 2, 106, -128, -22, 66, 90, -128, -24, -128, -73, -102, -15, 64, -13, 5, 114, 52, 59, -53, 12, 127, 43, 2, -128, 68, -43, -119, -58, 7, 80, -122, 57, -39, 86, -1, -128, -55, -92, -17, -69, -112, -124, -78, -81, -97, -3, 92, -16, 96, -128, -122, -123, 127, -31, 43, -101, 63, -68, 86, -17, -98, -3, 75, 79, -2, -8, 107, -8, -15, -34, 55, 74, -109, 24, 90, 88, -39, 70, -85, 22, -124, -128, -26, -64, -8, -116, -52, 36, 13, -7, 22, 54, 127, 13, 37, 113, 86, -64, -87, 127, 45, -85, -8, 127, 114, 58, -17, -15, -44, -114, -34, -23, 38, 127, 43, 98, -70, 88, -42, -66, -124, -31, 38, 81, 60, 10, 66, 116, 118, 0, 117, 50, 79, 24, 47, -66, 3, -97, -75, 47, 43, -15, -52, 12, -54, 0, 58, 74, -58, -107, 12, 127, 0, -33, 13, 114, -7, 43, -3, -48, 54, -17, -54, -128, -128, -128, -45, -29, -128, -81, 52, 52, 36, 64, 1, -74, 27, -66, 12, -17, -85, 98, -79, -3, -74, -76, 37, -117, -38, -11, -42, 13, 50, 127, 127, 66, 66, -27, 113, 113, 127, 127, -48, 58, -3, 73, -18, -1, -3, -54, -128, -54, 91, 39, 12, 49, 87, -63, 28, -106, -128, -122, -121, -3, -128, 12, 11, 24, -58, 3, 81, -75, 15, 29, -18, -128, -106, 112, 16, 11, -44, -101, -74, -47, 91, -33, 114, 28, -128, -128, -128, -74, 34, -128, -87, -13, 124, -36, -65, -55, -43, -116, -103, 79, -44, -36, -37, 6, -128, -93, -21, 38, -5, -128, -96, -64, 22, -50, 127, 127, 124, 127, 27, 58, -118, -87, 13, 127, 63, 64, 37, -53, -91, 22, 127, 1, -28, 13, 38, -119, 24, -13, -128, -32, -70, 117, -102, -97, -128, 76, 127, 47, -65, 39, 117, -63, 65, 17, 17, 53, 8, -8, -26, 65, -101, 55, 22, -128, -70, 69, -5, 13, 18, -111, -128, -39, -85, -92, -32, 114, -98, -69, 11, 96, -43, 34, 3, -34, 127, -32, 58, 32, 121, 78, -90, -121, -88, -2, 69, 28, 55, 13, -128, -88, 88, 76, -128, -15, -109, 109, -73, 37, -128, -10, 29, 26, -16, 127, 33, -90, -88, 5, -21, -86, -108, -38, 33, 127, 66, 96, -5, 38, 45, -50, 88, -128, -128, 48, 18, 88, -18, 86, -128, 127, 90, 97, -128, -10, -103, 52, -128, 37, 0, 76, -116, -108, -58, -121, -76, -128, 23, 0, -7, -52, -32, 127, -71, -29, -68, 60, -124, -85, 16, 15, 27, 6, 37, 111, -128, -103, -96, 60, -128, -64, 58, 31, -47, 13, 59, -78, 127, 114, -93, -39, 64, 106, -71, -75, 93, 127, -49, -128, -21, 63, -128, -73, 34, -66, -85, 23, -45, -122, 39, -32, -78, -78, -91, 2, -45, 38, -2, -128, -70, -12, 123, 27, 34, 100, -13, 116, 37, 98, -128, -124, -17, 127, 53, -52, -43, 15, 42, -70, 88, -13, -107, 47, -74, 117, 11, 55, -17, 47, 50, 53, -36, -39, -108, -7, 97, -128, -44, 38, 109, 0, 78, -3, -22, 48, 53, 109, -128, -17, -44, 80, -80, 107, -1, -107, -3, 44, -98, -128, -60, 74, 24, -27, -57, 28, -50, 90, 45, 127, 95, 87, -93, -97, -124, -31, 45, 103, -5, -80, -37, -3, 36, -22, 28, 81, -117, 55, 5, -33, -100, -80, -81, -38, -48, 127, -29, 93, 109, 127, -60, -8, -87, 127, -33, 127, -44, 23, -91, 12, 23, 102, 127, 59, 124, 55, 8, -86, 8, 121, -74, 124, 63, 22, -69, 75, 26, -45, 59, -98, 54, -68, -13, 24, 122, -49, 127, 118, -17, -44, -79, 74, -55, 59, -65, -2, -127, -100, 57, -57, -63, 44, -11, -69, -95, 65, -128, -29, -11, 127, -54, 52, 71, 23, -23, 45, 10, -124, 24, 69, 47, -93, 127, -75, 17, -128, -6, -128, -112, -118, -15, -92, -38, -23, -5, -127, 1, 28, 31, 10, -76, -18, -3, -34, -128, -29, 90, 11, -79, 127, 121, 91, 93, 80, 36, 98, -11, -27, -128, -29, 90, 44, -113, -116, -79, -117, -118, 29, 100, 78, 26, 68, 95, -5, -128, 76, 101, 85, -123, 76, -36, 28, -128, 27, -21, 3, -44, -107, 63, 59, 75, -45, -12, -8, -128, -43, -127, -54, 0, -52, -60, -106, -74, -101, 70, 78, -106, -81, 81, 118, 93, 39, 55, 73, 18, -117, -75, -114, 0, 43, 16, 8, -128, 29, -71, 108, 39, 79, 33, 0, -90, -128, 0, -128, 49, -128, 47, -112, 37, -107, -18, -5, 70, -7, 68, 127, 49, 127, 60, -3, 71, 127, 88, -39, -128, 0, -106, 85, 39, 37, -128, -128, 28, -128, -66, -97, 3, -116, -128, -111, -121, 127, -128, -103, -100, 102, -128, -64, -114, -24, -88, -87, 0, 74, 42, -112, -108, 71, 127, 127, 93, 76, 109, 45, 38, -107, 12, -128, -119, -124, 127, 28, 29, -93, 127, 44, 39, -28, 23, -70, 127, 13, 26, -2, 91, 106, 127, 127, 36, 69, 113, 122, -42, 127, -86, -44, -47, 96, 75, 127, 103, 100, -128, -128, -60, 127, 127, 55, -7, -22, 24, -24, -92, -54, -75, -128, -116, -112, 2, 31, 3, 23, -5, -128, -128, 64, 127, 71, -33, 66, 106, -128, -31, 7, 117, 70, 127, 124, 0, -60, 24, 109, 55, 113, -128, -28, -87, 68, -31, -111, -69, -123, -128, -39, 127, 3, -128, -49, 121, 97, -13, 23, -11, 29, -33, -128, -8, 11, 80, -32, 32, -24, -128, 8, -60, 117, -128, 71, 75, 86, -107, -128, -2, 127, 85, 58, -68, 95, -45, 127, 1, -66, -59, 17, 90, -65, -78, -119, -64, 90, -24, 49, -96, 114, -97, 48, -121, -66, -128, -112, -128, 7, -47, 1, -37, -2, -58, -21, 127, -113, -114, 37, 70, -128, -47, 101, 101, -38, -3, -8, 90, 127, 23, 127, 5, -10, -128, 15, -36, -10, -128, -55, -66, 58, -128, -70, 74, 34, -44, 117, 60, -128, -17, 127, 60, -27, -38, 106, 59, -31, 113, -29, 86, -53, -50, -80, -97, -93, -58, 97, 50, -34, -88, 127, -73, -79, -80, 127, -26, -128, -60, 119, 88, 12, 15, -32, 85, 102, 37, 92, -64, 45, -17, -114, -96, -122, 63, -39, 81, -88, 6, -43, -70, -42, -91, 127, 52, 108, -52, 107, 38, -5, -39, 37, 127, -31, 93, -76, 79, -92, -124, -74, 33, -27, -50, 95, 117, -128, -96, -111, 27, 2, 112, 18, -102, -32, 92, 74, 109, 58, -92, -47, 59, -111, -101, -52, -22, 127, 34, 64, -23, 78, 42, -26, 96, 127, 109, 12, -28, -24, 44, -102, -75, -114, -128, 16, 58, 0, -128, -128, -91, -128, 5, -80, 31, -53, 92, 118, -2, -38, 38, -3, -34, -81, 1, 91, -59, -87, 8, 37, -95, -60, -34, -59, 54, 71, 108, -127, -65, -50, 8, 1, 127, 78, 34, 37, 0, 111, 98, -8, -112, 23, 85, 29, 71, 127, -15, -128, -128, -128, -128, -66, -59, -128, -50, 127, 127, 12, -96, 90, 117, 24, 16, 111, -12, -74, -127, -8, -37, -52, -36, -42, 48, 79, -74, 90, -76, 95, 58, 38, 109, -21, 127, -3, 5, -36, 127, -45, -54, -111, -58, -15, 55, -34, -103, -91, -95, -69, 48, 65, -50, -21, -3, 13, -18, 127, 117, 75, -70, -15, -59, -64, 17, 60, -21, 53, -24, 5, 50, 122, 127, 86, 98, -55, 53, -122, -65, -27, 109, -28, -11, 101, 38, 85, -80, 80, -38, 127, -123, -100, -97, 80, 3, 55, 6, -76, -87, 44, -128, -121, -88, -108, -96, -33, 123, -116, 42, -71, 64, 8, 60, 0, -128, -88, -87, 111, -95, -71, -7, -49, -128, 1, 42, -8, -106, 127, 13, 123, -27, 60, 10, -6, 17, -88, -31, 23, -102, -32, -75, 127, -57, 76, -43, 127, 122, -128, -50, 53, 8, -124, -109, 107, -128, -26, 23, 90, -17, -29, -27, -31, 117, 2, 26, -114, -79, -39, 37, 92, -57, 127, 103, -65, 101, 86, 42, -106, 53, -57, -22, -103, -128, -128, -128, -128, -27, -95, -58, 17, -64, -13, -36, 34, -49, -122, 0, -60, -79, -68, 91, 107, 108, -63, 16, 37, 2, -96, -86, -15, 116, 22, 80, -32, 16, -8, -74, 10, -45, -100, 95, -33, 68, -60, 54, 88, 124, 49, -57, -45, -54, 64, 44, -5, -107, -16, 122, -12, 43, -1, 122, -1, 58, -74, 106, 127, 71, 127, 122, -15, -39, 127, 13, 24, -26, 108, -68, 37, -97, -88, -102, 47, 71, -32, -70, 3, 8, 39, 11, 87, -111, -37, 127, 42, 23, -64, 13, -80, -48, -16, 66, 127, 31, -128, -128, 92, 37, 0, -80, 26, 1, -38, 44, 81, 116, -21, 96, 28, 106, 34, -85, 44, -73, -74, 17, 127, 127, 27, -5, -128, 127, 1, 102, -88, 76, -128, -52, -128, 75, -119, 64, -60, -90, -128, 6, -66, 109, -70, 3, -128, -58, -58, 85, -122, 127, 75, 29, -78, 127, -58, -90, -38, 65, -36, -75, 127, 65, 45, -2, 127, 38, 127, 106, 70, -128, 39, 90, -13, -107, -58, -54, -23, 127, -18, 47, -47, 6, 13, 32, 127, 49, 34, -124, 98, -64, 108, -55, 119, 109, 70, 88, 112, 127, -5, 47, -55, 127, 127, 123, -71, -33, -45, 43, -71, -128, -128, -128, -49, -47, -5, -78, -39, 127, 52, -69, 28, 65, 91, -50, -76, 28, -49, -18, 127, 49, -63, -85, 119, 0, -24, -17, 127, 26, -10, -75, 59, -128, 127, 1, 53, -124, 26, -92, -112, -128, -11, -128, -109, -122, -128, 38, 43, 86, -76, 52, 7, -39, 101, 11, -52, -69, 2, 24, -92, 93, 0, -44, 6, -128, -43, -13, -18, -80, -128, 47, -33, 127, -32, -70, -95, -22, -26, -116, -113, 37, 127, 127, -128, -91, -100, 73, -6, -33, -44, 36, 86, 65, -44, -79, 44, 116, 92, -98, -18, 96, 29, -34, -128, -92, -128, 124, 101, 68, -128, -128, -112, -108, 116, 74, 91, -5, 2, -108, -128, -128, 36, 64, 53, -1, 57, 91, -69, 95, -122, -37, -107, 26, 70, 37, 17, -96, -3, 13, 39, 55, -52, 3, -44, 127, 107, 47, -100, 71, 91, -1, -128, -86, -108, 39, -128, -37, -124, 103, -23, 87, -13, 32, 106, 16, -57, 50, 76, 17, 12, -29, 80, 127, 117, -121, -128, -91, 38, 6, -87, 2, -1, -78, -64, 127, 52, 39, 96, 64, -128, -127, -128, -23, -106, 11, 21, 93, 98, -22, -44, -54, 45, -128, 36, -70, 75, -34, 97, 109, -78, 49, -8, -60, 92, 28, 53, -74, 113, 87, -59, -90, 8, -43, -128, -45, -49, 63, -93, -50, 45, -103, -63, 29, -73, -97, 1, -50, -119, -128, -112, -107, 32, -128, -90, -63, -92, -74, 32, -107, -106, 15, 103, 64, -38, -1, 53, 50, -118, 106, 57, -70, -128, -37, 73, 12, -117, -43, -79, 15, -10, -128, -2, 43, 0, -128, 27, -65, 117, -121, 127, 12, 48, -124, -1, -27, 78, 127, 127, 69, -42, 66, 127, 118, 95, -97, -2, -86, 91, -64, 24, 43, 127, 24, 42, -102, 107, -97, 16, -54, -33, -33, -128, -91, -109, -39, -100, -128, -37, 103, -24, -87, -50, 54, 42, -79, -106, -124, -49, 88, 123, -128, -23, -33, 127, -15, 52, -68, 2, -59, 39, 88, 43, 7, -100, -86, 127, 2, 127, -68, 127, -66, 111, 54, 127, 95, 47, -6, 60, -103, -36, -128, -93, 60, 34, 21, 69, 0, -36, -122, -85, -85, 21, -106, 64, 78, 24, -95, -96, -81, -50, 7, -43, -70, 68, -128, -49, -39, 101, 66, -60, 31, -39, 87, -68, 11, 66, -128, -91, -128, 47, 34, 127, -28, 1, 100, 75, 127, 23, 69, -128, 17, -100, 117, 63, -22, -109, 23, 28, 97, -95, 0, -57, 7, 45, -128, -107, -96, -48, -36, 95, -69, -128, 24, 63, 37, -42, 90, 37, -93, 71, 98, 76, 44, -122, -66, 36, 100, 66, 102, 127, 127, 32, 101, 48, 78, 45, 60, 88, 127, 52, 127, -113, 119, -87, -27, -59, 85, 47, -69, -81, -36, 117, 63, 43, -43, 80, 24, 15, -22, -114, -12, -128, 96, 16, 16, -73, 102, -16, 69, 47, -85, -13, 52, 117, -15, 127, 55, 26, -52, 127, 38, 87, 39, 107, 11, -15, -44, -93, -63, 29, 127, 74, -100, -106, 85, 127, 8, 0, 52, 74, 17, -128, -108, -118, 7, 28, 127, 50, -2, 48, 79, 0, 29, 127, -76, 43, -21, 127, 64, -128, -37, 108, 122, 21, -42, -39, -100, -128, -1, 17, 80, 39, -45, -90, -119, 75, -39, -128, -128, -96, 127, 102, 117, 55, 86, -128, -48, -54, 26, -128, -117, -102, -128, -103, 127, 13, 55, -42, 127, 60, 47, -53, -78, -128, -128, -18, 117, 59, -7, 63, 118, 24, -37, -1, -48, -78, -109, 76, -114, 103, -53, 127, 10, 8, 12, 0, -66, -33, 6, -73, 92, 0, -75, -34, -71, -101, 5, -95, 111, -13, 34, -101, -76, 23, 68, -128, -90, 47, 127, 127, 113, 87, 47, 127, 37, 127, -122, 12, -57, 81, -128, -36, -100, 3, -92, 85, 18, -128, -128, -127, -76, -127, -128, -81, 85, -22, -128, -7, -128, 101, -69, 73, -44, 68, 127, 28, -3, -50, -42, 90, -24, 11, -79, -124, -12, -38, -96, -128, 0, -128, 92, 102, 68, -33, 79, 0, -73, 11, 127, 29, -86, 7, 58, 127, -23, 127, 101, 127, -128, 70, -1, 123, 34, -71, 26, 44, 29, 96, -23, 66, 18, 103, 93, 113, -7, 127, 69, 127, 127, 69, 24, 98, 74, -70, -5, 8, -100, -92, 33, 108, -98, -80, -93, 28, 127, 127, 95, 81, 54, 127, 1, 102, -118, -45, -114, -70, 0, -128, -103, -44, 91, 127, 92, -117, -114, 108, 11, -128, -128, 36, -75, -128, -101, 45, -42, 0, -27, -13, 87, 73, -5, 52, 127, 27, 21, -66, 33, -80, -128, 0, -24, 127, 92, -3, -36, -49, 27, -71, 47, -109, -111, -128, -128, -128, -15, 127, 76, 28, -101, 101, 0, 109, 0, -18, 36, -57, -53, -60, 127, 100, 90, 18, 48, -128, -113, 64, 116, 60, 16, 50, -97, -53, 28, 102, -32, 3, -45, 15, -71, -24, -5, -124, 80, -79, 127, 24, -34, -64, -85, -107, 54, 122, -22, -128, -85, -36, -6, 31, 31, 52, -128, 12, -73, -50, -128, -70, -96, -43, -36, 127, 111, -17, 123, 119, 97, 12, 127, 127, -128, -75, -116, 60, -124, 98, -128, -98, -24, 127, -90, -122, 13, 117, -53, -66, 127, 74, -101, -58, 6, 127, -2, 43, -22, 38, 117, -121, -71, -95, 48, 43, 127, -37, -10, -43, 127, 127, 60, 65, 116, 52, 8, -96, -24, -68, 87, 107, -128, -108, 10, 121, 127, 117, 127, 57, 63, -24, 18, -24, -98, 127, -88, 43, -45, 127, -43, 12, -34, -47, -22, -80, 127, 17, 3, -98, 48, 0, 3, -93, 23, -108, 127, -32, 52, 113, 29, 54, -128, 108, -38, 80, -128, 127, -64, -34, -43, 108, 55, -42, 127, 64, -28, 64, -10, 116, -5, -24, -79, -47, 127, 127, 69, -34, 66, 111, -28, 93, -42, -128, -29, 6, 73, -69, 88, 102, 88, -39, 45, 124, 97, 127, -128, -31, -108, 106, -6, -74, -109, 73, -39, -95, -38, 127, 24, -75, -28, 127, 127, 48, -119, -109, 112, 42, -70, -128, -128, -50, -128, -80, -39, -5, -75, 127, 78, -32, -54, 91, -12, -128, -96, 127, 85, -53, -2, 65, 0, -95, -90, -92, -88, 68, -31, -128, -128, -6, 50, -128, -86, 27, -63, -13, 111, 59, 24, 108, 71, 39, 122, -38, -29, 45, 87, -86, 32, 18, 102, 102, 76, 81, 47, -76, 114, -24, 100, -66, 127, 34, 39, 76, 107, -47, -17, -69, 92, -75, 47, 63, -27, -69, -43, 69, -127, 112, -76, 123, 21, -24, -93, -7, -39, -60, -76, 57, 127, 119, 57, 55, 117, 127, 127, 39, -28, -58, 127, 39, 127, 39, 100, -103, -55, -92, 79, 47, 80, -21, -71, 8, -85, 36, 127, 8, -128, 11, 101, -10, -29, 103, 97, -64, -57, -109, 97, -55, -128, -79, 39, -53, -102, -18, 71, -127, -128, 116, -45, -10, -106, 91, -74, 36, 102, 119, -108, -128, -128, -47, -92, 12, -59, -102, -93, 54, 8, 50, 127, -33, 44, -85, -10, -1, 95, -95, 15, -26, 43, -128, -60, -128, -128, -73, 127, 71, -26, 74, 100, 127, 127, 112, -97, 6, 111, 68, 127, 15, 103, -75, 73, -75, -45, 33, 127, -13, 39, -27, 96, -114, -107, 37, 95, 127, 21, 43, -101, -31, 36, -27, 29, 53, -26, -32, -80, 52, 36, 16, -2, 85, 117, -71, -59, -10, 127, 42, 127, 127, 64, 127, 91, 26, -85, 26, -66, 23, 88, 58, -15, 127, -93, 108, -106, 71, 66, -37, -128, -108, 53, -78, -69, -128, -71, -21, -90, -10, -47, -2, -119, -7, -27, -27, -100, 64, -128, -73, -32, -81, -128, -31, -52, 123, 90, 39, -53, -128, 43, -90, -10, -128, 44, 42, 113, -43, 127, 13, -33, 54, 28, 107, -85, 44, -87, 100, 90, -3, -15, 127, 123, 69, -96, -18, 127, -45, -128, -78, 107, -17, -38, -31, 97, -49, 50, -45, -5, 127, 127, 127, 106, 55, 78, -13, 15, -122, 86, -103, -45, -85, -2, -103, 87, 101, -76, -70, -2, 42, 18, -119, -128, -93, 127, -15, 65, -79, 74, -118, 93, 8, -8, -24, 93, -44, -48, -53, -7, -75, -43, 98, 27, -23, -68, 127, 8, 16, 92, 127, 3, 88, 33, -44, -78, -12, 124, 127, -68, -123, -68, 112, 6, 90, 119, 2, -75, 127, -3, -64, -63, 53, -124, -123, 65, -45, 36, -7, 3, 95, 102, -28, -123, 108, 29, 127, -10, 127, -116, 78, -43, 127, 103, 127, -18, 123, -13, 53, 127, 65, 65, -44, 57, -79, -111, 22, -68, -128, -92, -128, -21, -31, -103, -102, -34, -34, 43, -74, -22, -128, 101, -122, -58, -118, -69, -58, -128, -128, -32, 53, -11, 17, -16, 86, 127, 127, 127, -45, 107, -27, 50, -68, -76, -92, -52, 26, 13, -2, 3, 57, 106, 127, -65, -128, 48, 127, 114, -28, 127, 127, 64, 98, 96, 50, -49, -93, 127, 101, 127, -57, 90, -2, 127, 87, 127, 109, 66, 34, 49, 112, -116, 127, 81, 57, -74, 69, -37, 75, 22, 54, -12, -128, -16, -124, 127, 127, 106, -78, 6, 127, 127, 127, 37, 116, 70, 85, -92, -128, -2, -73, 5, -116, 49, -97, 118, 97, -24, 24, -49, 63, -70, 76, 12, -116, -100, -128, 45, -128, 1, -92, 106, -22, 21, -16, 127, -36, 57, 6, 31, 44, -128, -114, 65, 127, 64, 0, -28, 71, -54, 118, -128, -8, -106, 48, 12, -48, -39, -38, 113, 49, -124, -74, 12, -128, -112, -73, -47, -112, -13, 43, 98, 93, 0, 54, 88, -118, 5, 5, 127, 74, 127, 127, 33, -96, 78, 108, 23, -90, -53, 27, 64, -107, 54, 116, -63, -93, 71, -5, -43, -92, 34, -29, -55, 39, -2, 64, -68, -113, 7, -122, 95, -128, -13, -74, 33, -21, 50, 81, 12, -15, 45, -44, 127, 90, 71, -60, 1, -15, 79, -10, -18, -42, 101, -101, 90, -1, 70, -33, -22, 102, 79, -50, -128, -97, -111, -128, 43, -107, 6, -70, 106, -48, -117, -31, -55, -128, -81, -32, 109, -29, 87, -109, 102, -122, 57, -45, 127, 8, -106, -128, -80, -73, 45, 78, -65, 103, -16, 37, -59, -60, -113, 48, 127, 127, 127, 111, 117, 13, 127, 24, 2, -128, -91, 127, 119, 53, -107, 65, 42, -117, -128, -108, -64, 42, 24, 109, -21, -22, 37, 66, -122, -96, -52, 5, -80, 31, -68, 88, -36, 127, -12, -13, 127, 91, 1, 12, 33, -128, -95, -108, -128, -53, -101, 127, -57, -116, -68, 73, -5, -128, 6, -63, 11, -39, 127, 101, 27, -128, -73, -75, -107, -24, 34, 113, 85, 78, -117, -118, 38, -12, -16, -128, -128, -11, 114, -37, -55, 22, 16, -60, 117, 127, -1, -119, -98, 32, -87, -18, 87, -10, -8, -33, 50, -116, 117, 0, 10, -66, 18, 100, 63, 63, 28, -24, -26, -23, -118, -88, -73, -1, -74, -21, 24, 127, 32, 76, 127, -2, -95, 93, 108, 127, -98, 127, -75, 127, 45, -54, -71, -114, 47, -43, 34, 59, 32, 28, -128, -87, 75, -86, -65, -128, -39, -74, -86, -69, -24, 70, 69, -16, -128, -91, -22, 95, -59, -128, -117, -91, -97, -128, -58, -117, 5, 12, 13, -95, -128, -128, 31, 34, 24, -128, -31, -118, 65, -15, 8, 8, 36, 96, -26, 112, 18, 49, 106, 45, 127, 121, 3, 6, 96, 2, 63, -53, -15, -93, 17, 54, 0, 52, -128, -117, -8, 11, 78, -17, 127, 119, 111, 38, 76, -8, -21, -108, -36, 43, 102, 96, 127, -107, -52, -48, 71, 101, -11, 79, 66, 50, -8, -69, 91, 69, -66, 13, 119, -52, 124, 127, 59, -69, -118, -31, -3, 103, -15, -75, 3, 108, -114, -128, -102, 7, -53, -87, 108, 127, 127, -28, 127, -3, 52, -127, 66, -37, -18, -123, -124, 28, -21, 63, -106, 79, -64, 22, 39, -16, 0, -16, 127, 59, 71, 107, 69, 22, -34, -42, -33, 127, 69, 127, 23, -18, -79, 24, 114, -128, -37, -48, 127, 69, 17, 44, 18, -10, 6, -59, -100, 95, 79, -128, -93, -70, 85, 23, 124, 48, -44, 70, 43, -91, -15, -68, 127, 127, 65, 23, 57, 90, 32, -114, -128, -42, -29, -69, -106, -21, 52, -124, -22, 33, 21, -49, -85, -50, 2, -128, -112, 21, 54, -128, -91, -47, -43, -128, 127, -28, 127, -119, 0, 44, 114, 127, 127, 127, -18, -39, -38, 106, 10, -58, -69, 127, 91, -75, -119, -81, -128, -97, -36, 117, -11, 18, -55, -57, 80, 127, 122, 87, 127, -7, 2, 21, 127, 127, -102, -128, -31, 23, -78, -109, 102, 43, 127, 63, 92, 127, -12, -8, 11, 108, -28, 54, -28, -11, 28, 81, -36, 127, 100, -57, -31, -81, -39, -128, 78, -48, 55, -100, -68, 91, -26, -87, 15, -116, -21, 23, 121, -58, 44, -128, -128, -79, -116, -107, -128, -75, -128, 34, -50, 127, -64, 122, 75, 127, 21, -23, -22, 48, -116, 59, 111, 63, 79, 127, 106, -95, -60, 64, 66, -128, 21, 78, 54, -81, -81, -74, -53, 90, 114, 33, -10, 127, 24, -95, -42, 123, 116, 97, 53, 102, 107, 21, -34, -59, -128, -27, 32, 123, -23, 127, 2, 47, 108, 123, -43, 70, -58, 96, 49, 66, -3, -79, -128, -55, 127, 90, -29, 34, -79, -11, -47, -81, -49, -88, 52, -15, 108, -128, 36, 24, 22, -78, 60, -64, -91, 3, 112, -43, 18, -65, -60, -128, -79, -2, 127, 122, 60, -37, -80, -79, -22, -128, -121, -65, 54, 37, 45, 17, -12, 12, -79, -10, -85, 66, 11, 32, -76, -128, -76, -58, -128, -80, -26, 75, 24, 112, 101, -101, 43, 10, 50, -13, 28, 69, 127, -88, 69, -108, -52, -128, -64, 16, 85, 50, 100, 33, -1, 23, 74, 15, 85, -91, -128, -42, -33, 2, -38, 23, 106, -13, 71, -45, 6, 26, -128, 2, -6, -101, -119, 59, -112, -13, 36, 55, 11, -92, -16, 0, 31, -37, 100, 127, -24, 127, -121, 65, -79, 113, 38, 47, 86, 122, 59, 12, -128, -78, 53, -95, -7, -90, 23, -73, 127, -55, -5, -102, -73, -117, -117, 78, 22, 127, 58, 0, 55, 123, 93, 118, 24, 37, 127, -6, -27, -38, 127, -65, 127, -8, 100, -128, -128, -28, 64, 127, -113, -123, -58, 80, 69, -63, 103, 73, -97, -76, 29, -36, 71, 92, 91, -44, 65, -116, -21, 49, 119, 127, -87, 81, -23, 45, 11, 127, 80, -97, -60, -36, -18, 37, -128, -128, 1, 96, -128, -87, -16, 127, 37, 43, -13, 127, 49, -127, -15, 97, 57, -31, 107, -1, 47, -119, 38, 6, -21, -60, -117, -54, -45, 86, -15, -114, 6, -10, 96, 28, 16, 98, 81, -128, -73, -66, -24, -128, -108, 12, -128, -124, -128, -1, -128, -123, 5, 16, 3, -15, 42, -17, -93, 78, 117, -16, -34, -44, 127, 54, 44, -97, 21, -54, 60, -88, -113, -128, -78, -96, 27, -17, 52, 43, 48, 86, 53, -23, 100, -11, 98, -11, -128, 0, -2, 16, -121, 18, 65, -24, -16, 66, -3, 36, 98, -92, -31, 38, 36, -128, -128, 45, -100, -33, -34, 66, 31, -75, 1, -128, -124, -55, 37, -10, 44, -75, -21, -109, 29, 116, 114, -15, 109, 117, 49, 49, -128, 98, -28, 71, -128, -79, -36, -116, -85, 91, 106, -6, -57, 124, 37, 109, -12, 78, -75, 69, -112, 32, -31, 32, 7, 54, 42, -44, -86, 87, 65, 118, 47, 42, -128, -47, -86, 42, -39, 44, 64, 1, 29, -80, 78, -10, 80, -31, 58, 0, 121, -37, 108, -64, 59, -87, -60, -128, -121, -128, 47, -44, 97, 107, 114, 54, -86, -50, -78, -127, -97, -58, -17, -69, -93, 78, 23, 59, -102, 124, 112, 29, -39, -53, 118, 69, 26, -128, 119, 53, 117, -97, 85, 100, 127, 66, 10, -33, 127, 66, 114, 127, 60, 60, -33, 59, 39, -33, -128, -86, -44, -13, -53, 17, -27, -12, -6, 1, -73, -98, -18, 79, 127, 114, 59, 15, 81, 29, 55, -128, -79, -69, 29, 55, 117, -18, -70, -78, -93, 24, -31, 91, -128, 127, 33, 1, -119, 127, 127, 123, -88, 49, -65, 21, -50, 8, -107, 18, -1, -31, -90, 127, 0, 100, -54, 127, 48, -15, 24, 102, 26, 97, 54, 7, -7, -44, -128, 43, -128, -60, -96, -128, -100, -54, -28, -73, -17, -116, 102, -57, 55, 42, 127, 127, -27, 31, -68, 87, -74, 10, -86, 42, -43, -59, -112, -44, -53, 49, 18, 109, 113, 127, -8, 127, 127, 127, -66, -5, -88, 109, 60, 64, 18, 93, 102, -39, 58, -75, 127, 16, 73, -26, -44, -111, 116, -27, -123, -92, -66, -12, -93, -42, -128, -123, -128, -27, 98, 42, -53, -36, 71, 10, -123, -28, -36, 22, 8, 64, -122, 57, 28, -118, -70, 127, 112, -3, 75, 112, 18, 16, -5, -114, -128, -88, -32, -128, -128, -93, -17, 97, -28, 102, -54, -38, -102, -33, 71, -29, 60, 127, -2, 87, 5, 111, -54, 76, -47, -10, 69, -2, -63, 44, 37, 127, -52, 16, -107, 127, -60, -78, -92, 75, -52, 127, 11, 17, -92, 112, -114, 107, 26, 74, -6, -12, -109, -106, 6, 59, 50, -32, -95, -78, 112, -57, 76, 54, 79, -76, 66, 16, 3, -123, 100, -48, -66, -66, 28, 97, -91, -49, -100, -123, 127, -60, 59, -128, 127, -47, 127, 27, 86, 42, -29, -23, -24, -50, -114, -122, -68, -128, -49, -12, -33, -44, 96, 39, -12, 127, 43, -128, -58, 88, 32, -111, -78, 75, 114, 13, 10, -116, 24, 47, -85, -102, -45, -100, -98, 127, 57, 79, -53, 85, -38, 106, 57, -58, 127, -55, -88, -70, 1, 54, 86, 58, -28, -29, 65, -128, -103, -12, 43, 15, 2, 22, -128, -102, -36, -1, 0, 90, 122, 22, 6, -91, -38, 27, 38, 100, -26, 15, 10, 16, -34, 50, -42, 108, -52, 127, -7, 13, -128, 0, -114, -43, 42, -23, -23, -97, 39, -44, -49, -44, 80, -50, -96, 127, 47, -39, -121, -21, -103, 127, 127, 100, -66, 127, 127, 27, 90, 108, 86, 127, 127, 87, 48, 49, 39, 10, 17, -12, -36, 79, 117, -123, 21, -103, 3, -80, 2, -27, -87, -37, 28, -39, -90, -121, 44, 127, 38, -86, -93, -128, -96, -128, 65, -122, 127, -8, 74, -93, 32, 0, -8, 55, 45, 127, -24, 36, 71, 127, 119, -88, 36, 0, 48, 127, 113, 78, -27, 127, 33, 18, -33, 27, -38, 75, -59, -49, -128, -128, -128, -57, -128, -128, -118, -27, -48, -63, -88, 127, 127, 17, -88, 27, 79, -128, 54, 90, 18, 27, 10, 39, -128, 127, -117, -17, -97, 98, 109, -128, -128, -108, 78, 78, -17, -27, 28, -98, 8, -74, -97, -95, 78, -1, 127, 71, 66, -45, 114, 127, 21, 111, -74, 121, -17, 24, -79, -78, -128, 98, 0, 12, -55, -73, -36, -49, -49, -32, 33, 127, 34, 63, -27, 85, 17, 64, -24, 63, 12, -49, -76, -128, -128, -68, -128, -66, -100, 78, -1, 81, 6, -85, -11, 98, 42, -128, -75, 32, -7, -66, 29, 16, -8, 91, 0, -26, 0, -106, -112, 10, 127, 60, 63, -15, 31, -128, -60, -121, -59, -128, -54, -128, -21, -54, 48, -128, -6, -79, -59, 44, 69, -22, -73, 114, 43, 108, 79, -29, -18, 86, 63, 74, 15, -26, -43, -106, -128, -63, 6, -2, -128, 33, -29, 109, -64, 127, 11, 95, -60, 76, 59, 37, 38, -116, -128, 16, -128, -128, -76, -2, -119, -57, 90, 10, -59, 11, -111, -101, -10, -32, -12, -71, -79, 121, 71, -75, 21, -90, -8, -87, -48, -68, -93, -32, -37, 75, 117, -57, 12, 54, 18, 59, -39, 85, 55, 127, 106, 8, 21, 90, 8, 29, 102, -96, -93, 12, 93, 112, 109, 127, 43, -78, -100, 11, 6, 64, -10, -128, -13, -114, -16, -128, -112, 73, 122, 13, 17, 88, 49, -18, 66, 87, 12, -24, -10, -71, -15, 127, -21, -17, -10, 74, -124, -91, 43, 127, 113, 124, 1, 122, -119, -85, -49, 7, 39, 8, 96, -128, 45, 114, 21, -112, -121, 95, -64, 102, 27, 75, 79, 6, 87, -128, -12, -8, 49, 22, 21, -79, -5, 107, -98, 15, 74, 45, 37, -60, 32, -50, 124, 23, 108, 63, 34, -50, -24, 116, -43, 7, 127, -31, -128, -122, 102, -102, -116, -66, -12, 127, 101, 111, -117, 49, 118, 74, -74, -13, -128, -17, -64, 36, -111, 45, 54, -109, -54, 63, 74, 112, 97, 37, 127, 26, 127, -26, 123, -70, 116, -64, -96, -111, -52, -37, 63, 95, 17, -128, 50, -43, 7, -121, -114, -12, 76, 38, -8, -53, -128, 96, -8, 65, -128, -18, 66, -81, 57, 59, 111, -128, 76, -73, -31, -21, -100, 54, -108, -63, -78, -114, 96, 32, 65, -33, 127, -39, 87, 31, 75, -78, 22, 127, 117, 95, -32, 127, 127, 18, 33, -42, -17, 74, 18, 60, -6, -42, -128, -102, 71, -17, -60, 10, 123, -42, -45, 121, 69, -71, -128, -111, -90, -78, -113, -102, 17, 66, -69, -128, -54, -98, 7, -22, 127, 96, 127, -29, 52, -26, 122, 63, -122, 86, 38, 28, -71, 96, -45, 122, 18, -87, -106, 0, 23, 8, -88, 127, 31, 95, 5, 97, 43, -71, 127, 31, 63, -45, 127, 121, 106, 79, 98, 48, -117, 29, 122, 36, -78, -42, 34, 97, 45, 127, -12, -128, -71, 44, -122, -108, -80, -128, -36, -31, 127, -6, -15, -50, 75, 47, 64, -15, 112, 69, -38, -2, 98, 39, -106, -21, 3, 53, 34, -32, -128, 1, 109, 23, -63, -75, 127, 74, 0, 64, 85, 80, -128, 44, -87, 122, -38, 10, 28, 91, -17, 33, 11, -100, -22, -47, 8, 50, -74, 90, 54, -23, -50, 8, 87, 2, 23, 63, 114, 53, 74, -52, -102, 127, 81, 60, -101, 124, -91, -7, -96, -8, 8, -54, -55, -111, -112, 73, -108, -29, -73, 2, -128, -121, -121, 6, 15, 54, -128, 44, 47, 97, -34, -37, 127, -28, -38, -128, -10, -42, -128, -117, 73, 88, -128, -97, 39, 39, -90, -75, -128, -128, -93, 34, -52, -79, -118, -128, -124, -108, 29, -69, 107, 66, 43, -59, 103, -97, -101, -86, 93, -59, 26, 107, -13, 103, -2, -42, -109, 15, -6, 42, -97, 8, -54, 127, 26, -93, -5, 64, 74, -113, 123, -44, 88, -86, 127, 17, 12, -112, -10, -13, -108, -38, 11, -128, -42, 23, 93, -75, -2, -54, 49, 119, 39, 87, 23, -48, -31, 64, 12, -2, -92, 92, 127, 73, 7, -24, 66, 17, 44, 39, 11, 1, 36, -50, 127, 16, 92, 64, 85, 1, -29, 47, -81, 68, -128, -78, -108, 107, -52, 80, 6, -128, -128, -109, 18, -81, -128, -85, -106, 28, -124, -128, -113, -11, 64, 64, 42, -122, -21, 59, 127, -53, 79, -95, 31, 49, 24, -23, 37, -59, 100, 36, -75, 47, -55, -96, -124, 15, -128, -26, -128, 52, -49, -31, -101, 74, 44, -102, -91, -69, 7, 68, 49, -24, 55, 95, -8, -128, -16, -55, -55, -88, -74, -6, -69, 101, 127, -69, -92, -47, 52, -42, 45, 127, -103, 103, -118, -70, -26, 92, 86, -63, 23, -122, -1, 97, -24, 55, 127, 57, -7, 127, 87, -81, -52, 100, 109, -18, 49, -96, 68, -71, -85, -21, -38, 27, 103, 90, 0, 54, -59, 11, -128, -128, -13, 71, 127, 65, -18, -87, -27, -128, -92, 47, -24, -128, -58, 36, -98, -47, 114, 103, 0, -5, -6, 42, -128, -15, 54, 12, -42, 88, 114, -10, 27, -113, -70, 87, 75, -50, -58, 93, 27, 127, -85, 108, -124, 13, -59, 80, 53, -44, -91, -2, 69, 59, -86, -6, 85, -128, 1, 10, -1, -92, 42, -80, -53, -57, -7, -79, 101, 47, 38, 85, 1, 92, -33, -128, -28, 70, 92, -68, 26, -86, -81, -5, -49, -113, -107, 29, 127, -63, -8, -69, 33, -74, 91, 127, 95, -98, -18, 127, 88, -48, -96, 58, 57, -106, -103, 103, 92, 79, -128, -96, -128, -91, -73, 111, 47, 68, 127, -28, 68, 18, 93, -38, 21, -10, -114, 33, 1, 96, -60, -24, -7, -26, 69, -73, -124, -128, -54, 27, 127, -90, 2, -128, 45, -128, -119, -81, 107, -6, 24, -44, 6, -54, -91, 24, 123, 57, -31, 74, -33, 24, -58, -36, -21, -50, 58, -1, 117, 28, -32, -124, 86, 109, -42, -113, -103, -6, -106, 34, -78, 65, 68, 127, 127, 127, 58, -36, 113, 78, 13, -128, 70, 13, -53, -128, -128, 52, -96, -17, -128, -107, -53, -45, -96, 54, 45, 106, 63, 79, -55, -128, 0, 97, 124, 31, 64, -23, -58, -55, -114, -42, -3, 70, 42, -114, 127, 127, 102, -101, -128, -36, 78, 102, 92, 31, 127, -128, 96, -12, 106, -101, 2, 65, 111, 44, -76, -100, -24, 86, 3, 97, -18, -52, -47, 10, 76, 32, -7, 117, 31, 33, -90, 16, 31, 93, 71, -118, -97, -3, 127, 114, 78, 1, 112, 96, 69, 32, -69, -85, -12, -116, -96, 127, 85, -54, -127, -1, 58, -34, -53, 42, -11, -70, 17, 34, -95, 0, -90, -78, 69, 127, 85, 34, -54, 127, 55, -60, 33, 0, -1, 119, 100, -10, 127, 28, -128, -80, 32, 34, -128, -118, -123, -95, -66, 127, 127, 66, 23, -128, 76, -128, -7, -80, -73, -54, 44, 79, -37, -91, -78, -119, -38, 50, 58, -22, -128, 100, 24, 27, -100, 102, -95, 5, 127, 100, 93, -48, 117, 66, -64, -45, 0, -124, -90, 90, 2, 127, 57, -57, -34, 27, 60, -74, 122, -5, -1, -128, -117, 17, -128, -128, -45, -28, -45, -86, -111, -69, -100, 63, 59, 69, 11, 27, -81, 28, -38, -85, 58, -58, -75, -18, 127, 90, 124, -128, 44, -55, 53, -39, 3, 24, -78, 38, -128, -1, -32, 127, -128, 17, -128, 97, -128, 114, 55, 73, -75, 113, 114, -43, -65, -128, -47, 8, 53, -34, -34, 5, -34, 127, 127, 74, -118, 21, 106, -16, -52, 127, 65, 63, -128, -26, -128, -29, -49, -111, -128, -26, 55, 60, -123, -52, -112, -128, -71, 102, 50, -75, 5, -42, -88, 124, 50, 58, -70, 127, 81, 32, 8, 111, 39, 73, -96, 85, 54, -128, -128, 21, -91, -22, -128, 68, -103, 127, -6, 38, -47, 13, 43, 50, 45, -85, -88, 79, -18, 18, 70, 0, 39, -70, -113, -45, 127, 102, 15, 43, 53, -47, -71, -90, -15, 3, 117, 44, -106, -128, -38, -102, -16, -7, 79, 127, 68, 36, -18, -3, -6, -18, 39, -107, 117, 38, 119, 29, -49, 81, 127, 50, 127, -11, -12, -5, 119, 86, -65, 68, 24, -27, 36, -11, -54, -78, -123, -128, -64, 91, 121, -73, -81, 59, 0, -75, -71, 87, -28, 2, 18, 3, 106, -117, -39, -95, -8, -119, -107, -7, -10, 37, -54, 96, -34, -42, -119, -81, 0, 11, 127, -48, 114, -124, -17, -43, 90, -91, -45, 75, 80, 68, 58, -68, 63, 92, 127, 59, 47, 124, 49, 60, -78, 73, -7, 42, 95, -73, 127, -108, 0, 5, 127, 73, 88, -50, 127, 103, -27, -64, 79, 69, -58, -10, 102, -10, -22, -119, 91, -3, -17, -85, 79, -128, 65, -5, 29, -54, 127, -23, 127, 33, 127, 32, 127, 92, 28, -22, -45, -128, -108, -27, 74, -121, -97, -103, -26, 114, 48, 57, -43, -108, -128, 5, -128, 24, -101, 48, -128, -27, 39, 36, -24, -23, -128, -13, -34, 127, 76, 124, 121, 127, 87, 5, 22, 86, -21, 60, 78, -2, 127, 73, -74, -33, 26, 127, 90, 100, -47, -90, 95, 44, -112, -113, -29, -93, -55, 75, -8, -21, -55, 64, -128, 29, 50, 8, -63, -128, -29, -42, 32, 23, 127, 86, 11, 50, 28, 108, 27, -1, -66, 71, 52, -65, -58, 127, -88, -12, 29, 79, 37, -59, 127, 12, -79, -122, -45, -128, -26, -11, -128, -119, 12, 8, -37, -3, 34, -8, -13, 15, -114, 10, -123, -117, -122, -116, 48, 66, 11, -52, -5, 127, 113, -21, 50, 31, -24, -21, 122, 47, 65, 107, -22, -128, -128, 57, 33, 36, -97, 39, 47, 106, 44, -106, -106, -52, 127, 31, 33, -71, 11, 127, 65, -18, 1, 103, -70, -71, 21, -27, 12, -26, 91, -85, -58, 2, 122, -69, 0, 60, 86, -73, -128, -81, 59, 10, -73, -10, 18, 43, 63, -80, -2, -113, 26, 127, 87, 49, 92, 50, -100, 92, -33, -42, 90, -2, 111, 33, 95, -45, -128, -49, -66, 11, -37, -68, -118, -76, 0, 23, 32, -1, 71, -103, -55, -10, 127, 55, -96, -124, -36, -128, -50, -123, 91, -111, -96, -71, -44, 45, 108, 64, -16, -5, 23, -47, -102, 49, -28, 127, -128, -53, -28, 114, -54, -58, 124, 127, 85, -66, -36, 31, 50, -128, -21, -81, 127, 42, 127, 49, 127, 100, 127, -70, -2, 21, 16, 31, -3, 119, -124, 22, -76, -59, -42, -71, -36, -63, 70, -49, -47, 66, 76, -11, 112, 68, 43, 127, 127, 59, 117, 16, 95, 13, 13, -55, -121, -86, 21, -128, 0, 17, 12, -90, -111, -43, -101, 86, 0, 127, 114, 88, 127, 88, 2, -58, 76, 21, 58, 87, 119, -24, -85, -128, -26, -66, -128, -124, -21, -128, -60, -12, -38, -107, -13, -58, -64, 44, -16, -90, -128, -43, -23, -122, -119, 44, -87, -128, -102, 42, 117, 127, 31, -44, 55, -1, -128, -128, 33, 60, 49, -29, -102, 71, 11, 37, 28, -128, 28, -85, 127, -112, 118, -36, 76, 43, -64, 90, -76, 127, -1, 127, 127, 27, -102, -88, -11, -128, -36, -7, -117, -39, -39, 127, 106, 50, 2, 49, 21, -63, 106, 108, -24, 103, 60, 48, 52, -22, -64, -27, -15, 2, -45, -128, -64, -107, -60, -128, 95, -68, 32, -96, -6, 79, -68, -76, 117, 53, -74, -12, 29, -88, 0, -98, -2, -128, -81, -81, 107, 3, -27, -44, 127, 60, 87, -53, 81, 114, -65, -42, -34, 93, -3, -11, 58, -31, 48, 58, 123, -128, 108, 2, 15, -101, 17, 17, -58, -98, 127, 53, -60, -63, -128, -54, -42, 76, -6, -128, 74, 34, 93, -85, 48, 127, 107, 42, -15, 93, 24, -128, -55, 16, 122, -55, 74, 97, 121, -42, 43, -34, 70, -78, 33, 75, -5, -109, -119, 18, -128, -128, 21, -52, -103, -90, 127, 79, 23, 65, -36, 87, -109, -87, -18, -90, 95, -95, -43, -54, -87, 85, -78, 45, -116, -114, 48, -114, 15, 50, 106, -128, -69, -128, 70, -78, 73, 0, 50, -85, 71, 29, 127, 123, -44, -71, 10, 118, -5, 43, -112, -50, -97, -64, -111, 58, -43, 127, 127, 39, -27, 16, 127, -13, -17, -50, 52, -102, -71, 109, 54, -70, 98, -42, 60, -128, 79, -76, 119, -116, 39, 7, 90, -49, -63, 127, 127, 93, 37, 124, 79, 68, 63, 69, -81, 81, -36, -128, -43, 2, -26, -107, 112, -5, 88, -12, -24, -128, -3, -111, -128, -128, -86, 37, -45, -92, 122, 95, 21, 24, -18, 127, -88, 17, -87, 108, -29, -78, 90, 122, -11, -50, 59, 17, -71, -71, 54, -23, -53, -124, -128, -59, 0, -112, 0, -29, 118, -26, 106, -63, -57, -79, 22, -128, -97, -113, -128, -73, 88, -44, -128, -87, -70, 127, -22, -87, -71, 31, -128, -128, -101, -80, 21, -42, 44, -128, -55, 26, 100, 5, -23, -95, -68, 73, -24, 73, -54, 127, 76, 96, -98, 49, -128, -123, -58, 66, -7, -29, 127, 59, 127, 92, 127, 27, -21, -108, -55, -23, -74, 116, -128, 54, -93, 127, 1, -3, -31, -39, -68, 127, 127, 97, -128, 91, 31, 123, -128, 6, -91, -37, -26, -87, 24, -24, -79, 100, 12, 96, -100, -103, 13, 121, -122, 33, -27, 65, -53, 100, 106, -81, -42, -103, -26, -128, -71, -101, -128, -39, 0, 60, -111, -59, 13, -68, 49, 76, -60, -90, 65, 96, 53, -128, -97, -92, 90, 66, 68, -128, -81, 2, 101, -101, 31, -109, 80, 34, 52, -32, 101, -59, -26, 127, 33, -128, -128, -32, 42, -85, -1, 127, 55, -124, 16, 109, 7, -78, -50, 38, -73, 54, 6, -55, 29, 59, -31, 47, 17, 88, -75, 127, -23, 85, 113, 127, 10, 100, -100, -37, -42, 55, -128, -13, -11, 117, 85, 42, 80, -47, -18, 16, 22, 88, -12, 1, -53, -128, 48, -81, 81, -58, 114, -24, -29, 127, 109, 3, 54, -1, 74, -6, 55, 85, 127, -68, 127, -100, 86, -102, 102, -124, -26, -45, -27, 34, -85, 10, -128, 79, -81, 100, -53, 57, -7, -69, -7, -52, 24, -15, -128, 24, 23, 16, 58, 109, 76, -59, 113, 79, -124, -28, -80, 127, 65, -7, -2, 118, 93, -63, -3, -58, -88, 29, 95, 54, 45, 58, -18, -48, 42, -65, -38, 81, 69, -18, -10, 21, 39, -53, 127, 58, -33, 44, 127, 127, 127, 43, -107, 48, 75, 1, -128, -87, -119, 81, -121, 79, -88, 124, -13, 127, 107, 28, -45, -47, 64, -112, -69, -10, 103, -128, 75, -128, -63, -128, 81, -36, -18, -116, 3, 127, -38, -50, -128, 127, 42, 127, -102, 101, -122, 6, -23, 59, 28, 53, 42, -116, 45, 85, 47, 39, 23, 127, 26, 49, -18, 54, -93, 103, -33, 37, -11, 53, 43, 127, 11, 100, 7, 23, -128, -71, -53, 127, -66, 78, -95, 112, -31, 75, 27, 43, 12, 98, 90, 112, 78, -128, -27, -86, 66, -85, -53, 24, -128, 127, -48, 123, -70, 18, 127, 80, 2, -36, 54, -32, 49, 117, 0, 127, -128, 71, -66, 127, -29, 29, -78, 127, 81, -58, -63, 52, -37, -13, 42, 69, 36, -11, 127, 18, 97, -10, -47, 118, 49, 127, -63, 127, 109, 114, -100, 127, 80, 26, -117, 60, -118, -106, -76, 2, 18, 127, 95, 127, 81, 73, -98, 70, -5, -48, -6, -75, -43, 69, 127, 10, -128, -66, 43, -28, -128, -128, -90, -7, 93, -128, -128, -128, 73, -38, -60, -121, 13, 44, -1, -42, -27, 21, -7, 18, 127, 100, 127, 124, 65, -29, 123, 119, 68, 127, 18, -43, 122, 127, 23, -10, 91, 106, 42, -69, -18, -32, 106, 50, 45, 127, 127, 90, 32, 114, 70, 127, 118, 69, -113, -33, 70, 98, -128, -6, -57, 107, 11, 31, 54, 7, 86, -128, 32, -66, 53, -117, -124, 34, -116, -124, -128, -128, -127, -128, -118, 43, 2, -109, -95, 36, -93, -102, 21, -37, 37, -37, -128, -39, -70, 54, 127, 78, 93, -80, 34, -64, 37, -47, 107, 1, 54, -97, -10, -26, 29, 29, -57, 107, 7, -69, 15, 71, 92, 127, -78, 47, -124, 21, -50, 81, -64, -63, -69, -65, 34, 15, -36, -128, -21, -66, 28, -121, 16, -5, 12, -1, -92, -69, -128, -71, -73, 59, -63, -100, -23, -112, 97, 60, -38, -43, -80, -8, -113, 58, -36, -90, 0, 108, 127, -81, 22, -98, 116, -75, -38, -75, 11, 59, 91, 10, 79, -58, 112, 116, 11, 114, 15, 93, 68, 101, 86, 127, 33, 127, -5, -21, -81, 119, -2, -15, -128, 43, -24, 70, -6, 96, 107, -1, -11, -91, -10, 108, 112, -1, 127, 42, -47, 66, 27, -48, 31, 95, 12, -128, -11, 127, 75, -111, -60, 127, -43, -65, -128, 63, -38, 107, -45, -66, 16, 127, 113, 78, 5, 118, 127, 63, -87, -73, 38, -37, -18, 100, 39, -102, 17, -70, 123, 127, 127, 16, -33, 2, 31, -128, -18, -17, -128, -47, -5, -11, -76, 16, 42, -90, 109, -128, 70, -96, 127, 0, 68, 52, 108, 48, -95, 23, -60, -128, -1, 88, 69, -128, -97, -13, 49, -2, 68, 66, -5, 57, 21, -79, 73, -76, 59, -63, -81, -128, -55, -112, 127, -106, -22, -18, 127, -114, 55, -52, 112, -103, 100, 88, 10, -23, -128, 74, -116, 92, -100, -39, -107, -59, 3, 28, 65, 23, -79, -85, -74, 127, 88, 127, 63, 23, -113, 124, 58, -24, -103, -34, 22, -37, -11, 48, -128, 21, -96, -100, -22, -34, 127, -128, 79, -73, -24, -75, -107, 68, -49, 13, -128, -65, 85, -34, -128, 52, 95, 127, 16, 119, -18, 127, 78, 119, -43, 93, -68, 86, -5, 127, -80, -112, 98, 127, 7, -44, -5, -2, 12, 64, -7, -128, 6, -58, 76, -71, 7, 26, 31, 92, 85, -34, -128, -122, 1, -91, -128, -76, -128, -48, -34, 95, -31, 127, 28, 73, -128, 49, -76, 33, -113, 97, -6, -128, -128, -11, -69, 33, -128, 17, -33, 50, -31, 69, -43, -1, 95, 127, 31, 103, -15, 39, -15, 59, 1, 87, -26, -16, 11, -24, 78, -114, 64, -128, -8, -23, 76, -43, 68, -128, -114, 54, 38, -124, -111, -87, 54, 70, 100, -88, -10, -116, 103, 54, 42, -101, 66, 0, 8, -32, -93, -52, 106, -18, 124, -3, 39, -5, 111, 127, 68, 43, -114, 127, 57, -44, -15, -15, 117, -81, 78, -91, -3, 18, 22, -55, 127, 127, 127, 127, 74, -36, -128, 48, 103, 71, -128, -127, -8, -60, -103, -116, -33, -128, -29, 127, 127, 76, 38, 127, 127, 69, -10, -21, 93, -109, -73, 127, 48, 112, -128, 127, -68, 127, -128, -12, -93, 69, -8, -32, 81, 3, -49, -58, 7, 95, -128, 37, 7, 32, -6, 49, 36, -121, 127, -86, 86, -21, 90, -63, -23, 6, 0, 32, 48, -128, -96, 76, 127, 58, -86, -10, 64, 127, 2, 112, -128, -66, -97, 27, -69, -73, 123, 5, 127, -112, -21, -57, 127, 85, -66, 22, 76, 24, -31, 113, 31, 103, 54, 11, 114, 27, 55, -76, 88, 90, 60, 28, -88, -45, -90, -100, -93, -76, -128, 28, -128, -27, -57, 127, 127, 74, -23, -103, 127, -112, -17, -128, -11, -64, 23, -74, -44, -8, -70, -80, 127, -15, 60, -2, 53, -3, 127, 127, 91, 36, 112, 85, 85, -113, -22, 17, 76, 80, 0, -5, 33, 109, -128, -128, -74, 49, -52, -128, -81, -128, -128, -97, 23, 65, 69, -36, 76, -92, -36, 119, -16, 88, 59, 127, -45, -93, 13, 88, 127, 7, 127, -48, 64, -87, 71, -1, 122, 127, 33, 127, -38, -128, -128, -71, -128, -16, 23, 23, -81, -13, -70, 57, 127, 48, 98, 96, 24, 38, -123, -33, -128, -102, 93, 53, -106, -128, 111, -75, 60, -101, 50, -128, 34, 12, 78, -128, -21, -128, -28, -116, 16, -50, -119, -128, -34, -34, 55, -15, -10, -65, -124, -85, -69, -71, -47, -86, -21, -60, -23, -39, 127, -128, 55, 13, 52, -128, -36, 27, 117, -18, 60, -33, -48, -52, 45, -60, -13, -16, -103, -33, 37, 45, 112, 70, 21, -123, -26, 127, 47, -32, -106, 10, -42, 24, 73, -128, -12, -79, 113, -63, 106, 5, 88, 127, 45, -118, 5, 59, -96, -78, 55, 17, -113, 33, -124, 12, 68, 76, 101, 11, 98, -128, -45, 127, 127, -66, -96, 38, 119, 1, -106, -37, -45, -108, 43, 127, 127, 96, 124, 73, 37, 10, 23, 127, 23, 96, -10, 98, -109, 127, 12, -8, -92, 37, -49, 127, 127, 118, -95, -81, -13, 121, 85, 0, -23, -11, -128, 24, 90, -10, -128, 7, 2, 109, -73, -93, 5, -15, -54, 10, 127, -7, 1, -12, 50, -128, -128, -90, -31, 127, 32, -28, -58, 78, 27, -26, -39, 121, 85, -109, -79, 119, 79, -128, -128, -88, 3, 103, 42, 0, -59, 75, 111, 127, -10, -52, -54, 48, -128, -109, 65, -59, -58, -27, -128, -36, -68, 127, -3, 93, -24, 127, 127, 112, 68, -8, 86, -31, -32, 87, 55, 87, -54, 45, -1, 116, 73, -106, -78, 39, 87, 95, 0, 80, -87, -75, 114, 7, 66, 29, 127, 117, 127, 98, 52, -26, 7, 127, 127, -12, 2, -3, 127, -111, 90, -27, 118, -12, -85, -106, 60, -34, -124, -27, 13, 38, -127, -93, -97, 1, -21, -47, 59, -128, 57, -57, 127, -128, 92, 33, 65, -112, -23, 108, -18, 15, 80, 73, 68, 127, 42, 50, 53, 127, 3, 1, -109, 47, -38, 127, 102, 43, -3, 127, 127, 97, 78, 0, 97, 10, -90, 68, 39, 37, 0, -124, 81, -21, 127, 75, 111, -121, -64, -55, 119, 2, -111, -76, -28, -76, -49, 80, 92, 127, 50, -7, -60, 113, 42, -81, -95, -78, 15, 101, 100, -47, -3, -13, 75, -26, -7, 5, 70, -102, 111, -106, -5, -34, 111, -11, 127, -12, -75, -74, 22, -10, -36, 42, -60, -112, 18, 15, -42, -73, -78, 100, -48, -38, -1, 87, -128, -37, -95, -103, -128, -113, -55, -33, -128, -21, 69, 127, 27, 36, -53, 21, 13, -128, -17, -128, -74, 10, -11, -124, -108, -36, 8, 97, 127, 57, 109, 8, 0, -5, 73, 49, -102, -103, 127, -8, -128, -128, 52, -128, -128, -107, 0, -81, -11, 27, -128, -2, -18, 59, 27, -42, 91, 34, 81, 45, 28, 112, 58, 48, -7, 119, 63, 1, 48, -117, -97, -65, -8, -109, 98, 121, 124, 43, 112, 127, 127, 49, -90, -117, -12, -66, 78, 18, -13, 73, -75, 5, -53, -128, -128, -38, 122, 100, -52, 50, 122, 116, 114, 91, 55, -128, -107, 34, -111, -45, -34, 88, -119, -32, 16, -47, 3, 101, 124, -57, -28, 127, 31, -128, -32, -12, -74, -123, 3, -34, 117, 127, -59, 68, -123, 60, -128, -108, -59, 52, 127, -13, -34, -10, 109, 74, -68, -87, -36, 32, -90, 24, 17, -128, -75, 60, 90, -107, -59, 50, 127, -34, 0, 7, 71, -8, 69, 100, 122, 108, 106, 116, 127, -106, 27, 95, 124, 88, -74, -90, -54, -55, 88, 43, 119, 65, -11, -15, 102, 8, -68, -103, -64, 45, 15, -103, -12, -98, -100, 10, 24, -47, 107, 87, -45, -23, 81, 53, -22, 58, 23, 39, 39, -7, -128, -78, 32, -27, -102, -65, -128, -33, -101, -128, -52, -128, -21, -74, 70, -121, 86, 96, 28, -128, -48, -12, -8, -87, 101, 31, -8, -36, -63, -52, -18, 65, 100, 58, -53, -28, 24, 12, 127, 44, 100, -24, 17, 127, 0, 57, -80, 112, 6, -47, 6, 81, 127, 1, -44, -45, -28, 5, 34, 45, -102, -128, 24, 127, 71, -108, 86, 96, 127, 90, 101, -17, 48, -26, -74, 36, 8, -73, -36, 24, 80, -128, -27, -119, 106, 5, 38, -64, -68, 0, -108, -58, -3, -96, -27, -128, -34, -5, -93, -16, -74, 42, -128, -100, -27, 38, -128, -21, -10, -66, -124, 32, -53, -47, -109, -70, 0, 127, 95, -42, -48, 78, 24, 71, -38, -91, -42, -128, 11, 6, 127, 127, 15, 52, -32, 13, -24, 127, 44, 85, 50, 18, -128, 16, 42, -8, -49, 69, 127, -100, 60, -109, 127, 106, 50, -3, 127, 95, -102, 0, -15, 55, -28, 108, 127, 127, 0, -49, -78, 66, 65, 127, 17, -95, -31, 32, -49, -127, -47, -95, -98, 0, 36, 101, 18, 17, -37, -100, -128, -38, -58, 87, -124, -128, -34, 65, -128, 27, 47, 86, -79, 127, 87, -78, -15, 127, 78, 70, 6, 127, -78, -16, -7, 71, -37, 43, 37, -97, 123, 127, 127, 118, -6, -128, -66, 127, 93, -87, -49, 87, 81, 98, 24, 42, 87, -44, 29, -78, 54, -88, -18, -101, 26, -65, -31, -53, 117, 32, -64, -33, -17, -21, -3, 127, 10, 85, -58, 100, 12, -128, -23, 69, 109, -45, 24, 123, 103, -64, -121, 28, 26, 54, -128, -91, -70, 3, 5, 0, 107, 58, 43, 44, -78, -66, 71, 31, -55, 12, 50, -66, -38, 45, -43, -70, -71, -111, 54, 52, -18, 0, 31, 68, -18, -3, 52, -128, 117, 39, 116, -43, 124, -48, -29, 109, 127, -124, -45, -109, 127, -26, 71, 16, 54, 0, -43, -44, 127, 81, 118, -37, -50, 127, 127, 114, 127, 95, 97, -47, 119, -98, -117, -103, -52, -59, 1, 101, 71, -1, 22, -64, -50, 59, 8, 124, -33, 15, -42, 49, 97, -10, 1, -65, -79, -48, -70, -128, -128, -114, -55, 93, 90, 81, 52, -91, -87, 1, 127, 103, -5, 127, 50, 8, 122, 127, 18, 112, -16, 95, -106, -21, 58, 47, -42, -66, 127, 85, 127, -112, 85, -27, 127, 7, 127, -10, 17, -55, -71, -57, -111, 113, -10, -36, -128, -102, -42, -74, -112, -74, -128, -69, 93, -63, -66, -43, 127, -101, 121, -12, 106, -5, -76, -58, -37, -128, -128, -128, -66, -48, 68, -18, 73, -128, 96, -5, 119, -45, 127, 49, 69, -26, 55, -11, -128, 59, -91, -47, -118, -128, -95, -58, 127, -7, 23, -57, 26, -73, -36, -114, -59, 127, 127, 63, -45, 71, -12, -128, -127, 114, 119, -44, -97, 127, 87, 33, -128, -18, -90, 127, 42, 107, 18, 98, -39, -50, 8, 22, 123, -93, 36, -38, -13, -128, -128, -87, 29, 108, -128, -85, -107, 127, -100, 47, -106, 127, 15, 44, -28, 75, 103, 59, 73, -10, -31, 53, 79, -108, 58, -13, 27, -54, -78, -53, 26, -109, 97, 45, -70, -36, 37, -16, -102, 123, 79, 68, 5, -3, -101, -76, 39, 127, 64, -78, -100, -128, 26, -117, -53, -66, 52, 11, -68, -10, 34, 98, 106, 111, 17, 63, -91, -128, -128, -103, -96, 127, 8, 118, -128, -38, -57, 49, -101, 6, 11, 42, -18, -80, -73, 11, -86, -36, -91, -75, 107, 42, 127, 78, 43, 17, 65, 60, 75, -32, -113, -34, 23, -128, -128, -63, 127, 87, -128, -87, 127, 127, 60, -32, -66, -16, -98, -106, -108, 28, -86, 88, 109, 98, 127, 55, 118, 102, 127, -21, 26, -87, 112, -52, 59, -49, 109, -109, -118, 81, 73, 127, -17, 127, -1, 66, -112, -24, -101, -8, 75, 6, -38, -27, 112, -73, -80, -34, -102, -52, -65, 92, -34, -39, 48, -128, -128, 0, 21, -42, -108, 127, 49, 15, -79, -121, 21, -47, 16, -60, -81, -85, -29, -128, -79, 23, 34, -128, -76, -118, 91, -90, 74, -21, -28, -21, 127, 27, 1, 122, 127, -98, 79, 6, 112, 8, 127, -38, 28, -87, 43, -128, -50, -58, -128, -128, -128, -128, -111, -128, 74, -121, 48, -23, 96, 49, 58, 81, 68, -5, 127, 37, -76, 39, -34, 87, -87, -45, -90, -22, 121, -29, 87, 7, 127, 21, -119, 10, -49, -63, -76, 16, -81, -29, 114, -71, 45, -59, 127, 60, -53, -113, 114, -55, 121, -116, 22, -96, -45, 63, 52, 124, 55, 79, -52, -128, -88, 47, 6, -128, -63, 116, 127, 90, 95, 95, 73, 127, 24, 0, -112, 13, -85, 47, -75, -93, 127, 15, 70, -26, 53, 96, 17, 39, -128, -116, -49, -8, -98, 6, -34, 58, -70, -102, -57, 60, -95, 96, 127, 43, 54, -70, 74, -73, 127, 18, -31, -18, -32, -127, -90, -31, -59, -127, -124, 85, 39, 103, 8, 10, 113, -34, -58, -128, 68, -85, 28, -128, 8, -48, -26, -128, -80, -58, -31, -85, 102, -75, 44, 121, 75, -60, -128, -128, -63, -78, 42, -128, -59, -70, 103, 1, 124, 95, 33, 102, 50, -64, -85, 90, 54, 23, 127, 47, 100, -22, -2, -88, -96, 96, 114, 127, 127, 117, 70, -50, 127, 91, 52, 96, 74, 127, -75, 0, -97, 103, -85, 8, -103, -26, 8, 127, 93, 17, -49, 5, -97, 87, 28, 97, -11, -81, -48, 68, 6, -87, -128, -108, -48, -65, -79, -90, -101, -97, -26, -123, -118, -66, 60, 79, -47, 119, 52, 112, 29, -26, -128, -45, -76, -39, -128, -54, -65, 127, 29, -29, -80, -28, 11, 11, 97, 47, 86, -42, -58, 24, 27, -57, -64, -54, -33, -101, -114, -65, 8, 78, -68, 1, -68, -128, -58, 127, -24, -108, -124, 60, -33, -15, -128, -38, 12, -18, -48, -42, 13, -128, 95, -128, 32, -128, 45, -58, 74, -128, 79, 59, 127, -92, -128, -74, 64, 119, -29, -3, -112, -128, 21, -11, 39, 31, -47, 33, 11, 87, 116, -50, 81, -118, 66, 38, 127, 39, -6, -15, 116, 80, -119, 48, 119, 122, -10, -127, -107, -68, -66, 1, 71, 29, 52, 37, 100, 69, -128, 75, 74, 113, -128, 47, -54, 22, -76, 98, 32, 127, 34, -128, -128, 8, -128, -128, -128, -65, -50, 69, 45, 74, -93, 15, 27, -45, -111, -122, -80, -5, 23, 34, 3, -85, 64, 85, 127, 122, 28, -15, 74, 29, -113, 44, -18, -71, -32, -55, -70, -8, 101, -128, -32, -113, -3, -21, -128, -119, -103, 97, -123, -107, -98, 27, -106, -27, 36, 21, -36, 54, 97, -53, -128, -128, -97, -54, 23, -79, -26, -50, -34, 92, 11, -95, -102, -60, -128, -101, -91, 42, 98, 53, 63, -90, 26, -44, 121 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
