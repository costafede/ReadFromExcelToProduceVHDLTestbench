-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            41, 91, 16, 40, 45, 82, -48, 33, -62, -103, 107, -14, -119, 53     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( 39, 99, -116, 97, 18, 105, -80, 69, 61, 49, 36, -82, -17, -6, 95, -52, -37, 105, 70, 123, -11, -91, 104, 7, -31, -49, -19, -6, -65, -113, 45, 126, -96, 92, -44, -113, 82, 101, -30, -78, -107, -117, -40, -7, 41, -119, 112, -97, -4, -67, 10, 25, 58, -81, 32, -75, 3, -40, -123, 8, -8, 5, 114, 111, 72, 36, -39, 14, 12, 124, -49, -118, -124, 33, -20, -35, -37, -20, 37, -2, 122, 40, -120, -101, -36, 75, 66, 98, -95, 78, -4, 69, 49, 4, 51, -117, 74, -77, 20, 34, -6, 97, -34, -45, -94, 61, -101, -11, -89, 62, 55, -110, -25, -49, 42, 101, 31, 103, 91, -9, 22, -34, -53, 123, 30, -8, -107, -42, -72, 118, -59, 115, 5, -57, 125, 107, 80, -84, 81, 41, -10, 126, -102, 100, 17, 9, -100, 77, 9, 12, -53, 42, 78, 27, -109, 120, -38, -23, -107, -117, -33, -36, 71, 56, -90, 19, -7, -20, -63, -37, 89, -28, -7, 110, 69, 23, 26, 34, 96, 18, 60, 94, 8, -60, 106, 16, 47, 85, -14, -88, 24, 46, -121, 88, 72, 78, 49, 6, 34, -102, 31, 75, -128, -72, -17, -11, -32, -120, -33, -53, 106, 89, 8, 105, 37, -55, -23, 51, 83, -59, 66, -89, -18, 94, 77, -41, 47, -118, -90, 57, -103, 16, 82, 27, 16, -108, -54, 21, 98, -60, 84, 76, -19, 37, -126, 18, 98, 7, -125, -29, 69, 64, 125, -48, -21, 97, -71, -92, 62, -14, -14, -14, 80, 16, -48, 67, 100, -123, -89, -126, 50, -71, -30, -81, 112, -103, -127, 20, 98, -83, -79, 8, 54, -58, -28, -2, 21, -110, -92, 79, 59, 61, 8, -32, 119, 124, -3, -22, 27, 124, -66, 123, -95, 56, -73, -96, -52, -101, 106, 33, -104, -34, 103, -5, 22, 126, -52, 73, 40, 57, 81, -74, -79, -55, -127, -36, -91, 110, 88, 122, 36, 83, 2, -3, 41, 61, 47, -45, 92, -6, -86, -21, 54, -68, -104, 98, 0, -49, 119, 79, 100, -64, 96, 25, 29, 123, 83, -6, 48, 92, -38, -110, 56, -14, -14, -16, 123, -127, 111, 120, -95, -40, -4, -12, 106, 26, 51, 30, -39, 33, 28, 56, -21, 23, -98, -21, -34, -120, 52, -64, 111, -61, 105, 2, -116, -105, -53, 67, 122, -63, 83, -116, -102, -91, -95, 31, 80, 29, 21, -26, -102, 50, -97, -13, 104, 125, 65, -33, -10, 76, -106, 47, 30, -71, -4, 54, -80, 35, 87, 99, -20, 37, -112, 119, -98, 92, -78, -72, -49, -90, 72, -114, -123, 24, -107, 45, 80, 68, -70, 53, -60, 98, -107, 44, -94, -51, 95, 30, -2, -91, -96, -89, 28, 56, -125, 81, -108, -34, 75, -125, 48, -102, -119, -33, 68, 1, -80, 62, -104, 98, 66, -3, 119, -97, -121, 117, -34, 123, -5, -13, 2, 93, 101, 39, 63, 97, -116, -114, 119, -49, -106, 95, 78, 68, 113, -46, 118, 30, 11, -12, -43, -21, 83, 18, 125, 70, 78, 119, -119, 31, -110, -70, -97, 2, 4, -64, 88, -111, 70, 125, 109, 84, -81, -97, 119, -48, -36, 121, -99, -92, -77, -40, 91, -69, -56, -10, 81, -22, -123, 50, 28, -105, 99, 13, -117, -9, 107, -83, -120, 78, 13, -52, -60, -15, 4, 69, 101, 105, -95, -24, 117, -24, 79, -69, -42, -87, 81, -56, -64, -35, -68, -70, 123, 23, -14, -109, 11, 24, -106, 10, -8, 91, -114, 72, 71, 26, -76, 35, -63, -19, -94, 56, -98, 28, 41, -35, 66, 91, 113, -87, -125, -122, 99, 25, -34, 90, -21, 114, -53, 15, 51, -125, 47, -62, 42, 24, 126, 11, -62, -93, 9, 3, -128, 4, -5, -16, 10, -15, -72, -63, 73, 20, -118, 126, -86, 12, 44, -86, 61, -52, -98, 48, -122, 84, 58, 17, 69, -118, 113, -118, 117, 79, -32, 57, 12, 65, -54, 24, 38, 21, 84, -3, 75, 127, 67, 37, -119, 57, 38, -50, -36, -86, 93, -50, -98, 124, 62, 92, -65, -125, 40, 43, 125, 10, -12, 41, -107, -115, 0, 44, -28, 94, -106, -50, 15, -128, 63, -126, -96, 80, 103, 46, -47, -121, 77, 28, -110, -51, -26, 102, -89, 64, 124, 54, 27, 114, -94, -56, 104, 52, 49, 101, -123, -24, -7, -16, -36, -26, -114, 59, -46, -43, 9, -94, -119, 86, -70, -86, -64, -20, 19, 21, -72, 127, 31, -68, -67, -122, -58, -6, 100, 21, -124, -84, -106, -55, 15, -26, 123, 123, 77, 118, 51, 41, 13, -33, -43, -1, 48, -63, 10, -21, 71, -56, 49, -91, 93, 2, -65, 49, -13, 43, 99, 44, 44, -98, -57, -21, 56, -98, 17, 114, -104, -42, -66, 42, 121, -109, 118, -90, -101, 31, -65, -4, 100, -82, 24, 79, -7, -71, -101, 19, 99, -71, 99, 51, -65, 54, 124, 14, 104, 55, 124, 86, 60, 20, -46, -27, -71, 35, -95, 86, -73, -78, 74, -20, -6, 74, -127, 96, 67, -69, -78, -96, 10, 39, -110, -69, -62, -28, 1, -49, -94, -71, -16, -119, -72, 63, 113, 93, -1, 27, 27, 93, -23, 43, -34, -59, 46, 105, 63, 66, 124, -31, 59, 34, 37, 124, 126, -116, 25, -67, -80, 8, 48, 85, 94, -54, 16, -42, 28, 68, -68, -84, 115, -4, 14, 96, 123, -41, 20, -103, 48, 44, -60, -95, 34, 25, 46, -10, -15, -57, 99, 18, 71, 30, 22, 38, 73, -13, -105, -113, -5, -104, -87, -9, 97, 118, 24, -73, -11, 53, 47, -98, -122, -72, 110, -98, -60, 68, -96, -84, -104, -128, -88, -85, -57, 90, 69, 79, 125, -116, 90, 96, 5, 110, 78, -116, -126, -93, 125, -122, 125, -57, 49, -45, 11, -30, 53, -1, 18, -42, -39, 67, -35, 52, 21, 61, -66, -102, 106, -15, 116, -72, 90, 44, 31, -63, 34, 0, -38, 61, 95, -63, -36, 20, 86, -40, -12, 57, 24, -23, 109, -1, -105, 86, -47, 51, 32, -43, 40, -89, -100, 13, -119, -46, 115, 114, -23, 51, 21, 38, -38, 87, 23, -97, -102, -56, -19, -112, -105, 46, -103, 106, 116, 58, 73, 36, -87, 105, 45, -98, -105, 101, -128, 50, 29, -104, -120, 119, 16, 58, -55, -38, -82, -3, -74, -127, -12, -91, 68, 125, -38, -44, -86, -75, -61, 42, -98, 43, -35, 32, -87, -105, -128, 76, -127, -87, 0, -82, 24, 116, -114, 5, -50, -38, -109, -113, 62, 92, 62, -34, -99, 13, -61, 61, 1, 66, 109, -10, -34, -58, -116, -67, 104, 65, 77, 71, 22, 46, 6, -111, 105, -29, 63, -14, -106, 21, 119, -124, -21, -101, 121, 79, -11, 12, -50, -85, -55, -39, 60, -118, 41, -42, -77, -92, -50, 108, 30, 57, 77, -54, 36, -126, 28, -92, -34, -28, 117, 80, -22, -2, 109, 49, -106, -54, 101, 42, 30, -125, -56, -89, -8, 65, -39, 72, 81, -20, 55, -46, 30, 124, -77, -17, 32, 79, -60, -96, 14, -97, -15, 49, 33, -124, -85, 116, -115, 98, 80, 58, -108, 45, -40, 111, -18, -83, -8, 65, -17, -74, -90, 0, 7, 62, 125, 5, 13, 34, -124, -44, 126, 96, 99, 55, -108, -53, 8, -44, 19, -51, -14, 16, -63, -40, -91, 126, -53, 60, 67, 74, -43, 124, -119, -96, 125, 85, -6, 94, -10, 46, 93, -28, 113, -70, 1, 35, -2, -44, 34, -81, 10, -28, -7, -92, 7, 81, 34, -86, -14, 48, 31, 54, 8, -80, 64, -127, 61, -6, 14, 86, -116, -3, -66, -104, -101, -4, 106, 116, 2, -98, -8, -31, 91, -108, -27, -29, 17, 127, 96, 57, 28, 50, 6, 89, -91, 102, -54, 124, -55, 29, 49, -59, -115, 20, -28, 100, -49, 104, -122, -128, -54, 22, 72, -94, 124, 86, 78, -93, 28, -124, -75, 52, -51, 66, 104, 101, 12, 3, -74, 42, 0, 30, -50, -112, 2, 118, -2, -79, -63, 114, 62, 14, 55, -109, -35, 118, -70, 119, 108, -23, -20, -127, 85, 60, -2, -66, 119, -19, 15, -5, 32, -109, -69, 34, -10, -63, -65, -62, 45, 19, -50, 10, 85, 73, 58, -46, -125, -115, 41, 62, -65, 119, -46, -117, 77, 95, -96, -123, 45, 109, 21, -68, 97, -47, -100, -123, -67, -103, -30, 81, 42, 108, -16, 28, 24, -104, 27, 90, 61, -47, -16, 34, -7, -6, -25, -85, 83, -55, -92, -75, -98, -85, -24, 87, 34, -41, 67, 20, 95, -90, 59, -80, -57, -8, -126, -108, -77, 34, 115, -37, -118, -22, 119, -73, -108, -94, -60, 59, 36, 19, -54, 79, -28, 71, 106, -88, -73, 9, 29, 22, -117, -96, -57, -55, 11, -42, 76, -86, 111, -41, 120, -76, 33, -96, 37, 121, 89, 108, 88, 38, 120, 18, 43, 44, -113, 21, -20, 6, 57, -79, -3, -91, 59, -7, 18, -80, 62, -49, 28, 73, -93, -116, 22, 24, 10, -13, -114, -110, 24, 102, 123, -104, 68, -27, 82, -86, -39, -58, -39, -74, 71, 39, -26, -91, -75, -113, -19, 79, 39, -4, -4, 113, 22, -37, -62, -66, -43, -73, 48, 97, -110, 127, -76, -2, 49, 81, 126, -38, -86, -110, 93, 114, 52, 114, -93, -46, -6, 95, 58, -71, -44, 24, 33, 109, 59, 119, -34, -126, 68, -105, 103, 43, -95, 62, -106, 116, -35, -1, -124, 33, -107, -46, 67, 25, -34, -121, -33, -33, 66, -73, 103, 59, 118, 89, -38, 9, 125, -16, 17, -21, 82, -114, -5, 14, -12, 85, 91, -8, 2, 81, 11, -106, -96, 0, 103, 119, -96, 12, -77, 78, 81, -42, -52, -98, 56, -14, 26, 107, 105, -87, -50, 99, -121, 55, -19, 37, -68, -107, -43, 39, 48, -96, -39, 123, 54, -114, 10, 65, 91, -8, -104, -58, 41, -74, 86, 106, 80, 83, 108, -102, -8, -46, -2, -76, 97, 108, -86, 45, -86, -97, -58, -105, 19, -127, 116, -4, 29, 112, -120, -103, -45, 53, 16, 58, -80, -113, -76, 96, 60, 91, 125, -44, -99, 46, -115, -64, 21, 87, -61, 60, -5, 15, 67, -12, -4, 30, -51, 117, -112, -47, 118, 34, -87, -47, -98, 119, -12, 106, 59, 85, 104, -43, 13, 52, -49, 91, 35, -87, -83, -6, -124, -36, 66, -79, -95, -95, 38, 60, -30, 12, -96, 16, -1, 116, 24, -44, -31, -105, 99, -74, -63, 27, 29, -99, -128, 127, 48, -114, -16, 59, -70, -115, 111, -103, 103, 111, 63, -110, 71, 62, -18, 108, 11, -5, -16, 10, 3, -69, -74, 3, 113, 88, -25, 83, -68, 52, -72, 24, 98, 116, -124, -86, -65, -13, -17, -14, -30, 93, 14, -106, 23, 112, 89, 58, -121, 80, 15, -93, 61, 92, 71, 58, 77, -9, 84, 16, 14, -57, 53, -97, -113, -12, 6, 19, 126, -74, 94, -124, 116, -44, -54, 60, 115, -81, 59, -45, -122, 4, 20, 13, -80, 60, 37, 82, 15, -9, -117, 106, 50, -90, -89, 59, -104, 64, 50, 101, 67, -105, -18, 12, 1, 17, -118, -25, 81, 100, -91, -75, 77, 84, 118, -53, -87, -68, -67, -96, 119, 66, 117, 56, -120, 57, -25, -20, -118, -83, 0, -113, -88, 74, 119, 32, 31, 67, 107, 71, 114, -2, -76, 17, 70, 6, -23, 74, 115, 122, 59, 2, 113, -29, -67, -71, -35, 19, -41, -28, -58, 8, 38, -40, 30, -72, 4, 102, -30, -9, -71, 112, 54, 49, -102, -27, 6, -23, -23, 40, -42, -99, 70, -70, -48, -67, -98, 11, -101, 23, 75, -113, 119, 62, 8, 14, 54, -34, -120, -16, -52, 41, 8, 18, -117, 108, -29, 34, -94, 54, -117, -111, 76, -40, 81, -99, 106, -28, 110, 7, 48, -94, 14, 57, 103, -104, -1, 105, -27, -86, -82, 33, -1, -86, 113, -71, 30, 80, 32, 44, -114, 90, 35, -5, 67, 11, 66, 68, 27, -45, -5, 85, -31, 107, -70, 51, 121, 10, 41, -14, 66, 28, -44, 46, -99, 20, 92, 117, -14, -23, 14, 23, 57, -35, -114, 16, -77, 98, -32, 80, 24, -2, -91, 85, -45, 123, 99, 25, -56, -62, 35, -116, 79, -38, -88, 89, -94, 103, -118, -21, -112, -32, -18, -107, -76, 38, 126, 34, 84, -54, 62, -117, -117, 21, -1, 45, -103, 6, -119, -54, 84, 72, -47, -60, -46, -88, -65, 52, 86, -45, -21, 6, -32, 107, -112, 93, 22, 61, -104, 2, 125, 4, -112, -80, -50, -95, 89, -96, -79, -49, 3, 56, -40, -89, 65, 13, -119, -114, 97, 78, 20, -3, 83, 57, -63, 125, 110, 114, 92, 49, 105, -41, 95, -36, -112, 75, 89, -80, 69, 78, 51, 12, 120, -68, -122, -12, 51, 38, -37, -24, 119, 120, 82, -24, -35, -22, 8, 54, 106, 16, 113, 15, 123, -4, -93, -17, 26, 68, -57, -93, 78, 72, 88, -65, -109, 86, -73, -52, -83, -66, -76, 22, 37, 97, 43, 61, 52, 95, -89, -39, -24, -115, 45, 71, 41, 85, 126, -93, 70, -109, 111, 104, -98, -121, 122, 18, 18, -19, 22, 74, 25, 99, -65, 89, -127, 29, 42, -126, -4, 67, 116, 78, -103, 57, -6, -64, -103, 46, -80, 20, 84, -56, -47, 78, 5, 92, -46, 108, 63, 75, 56, -28, -108, -32, 95, 24, -109, -96, 75, -66, -68, 51, -52, 83, 84, 13, 55, 85, -64, 83, -29, -71, 4, -125, 107, -87, 58, -100, 31, -18, -81, -9, -99, -8, -76, -106, -66, 83, -50, -19, 119, 106, -122, -44, -25, -43, -93, -16, 4, -25, 114, 83, 70, -36, 17, -105, 87, 62, 14, -30, 72, 20, 3, -22, 117, 38, 87, -30, -43, -17, 97, -67, 95, 44, -23, -103, -45, -68, -9, 83, 18, -119, -62, -82, -110, -32, -66, -31, -56, -123, 9, -127, 115, -119, -120, 112, -18, 47, 58, -34, 88, 106, 4, 24, -99, -96, -45, 70, 80, 79, 63, -60, 54, -11, -104, 59, -36, 48, 123, -50, 47, -16, 127, -51, 115, 92, -36, -27, -97, -87, -109, -14, -34, 54, 110, 119, 96, -17, 100, 53, 59, 49, -112, -32, 118, -86, 9, -78, 8, -60, 54, 0, 74, 63, -72, -17, -41, 24, -62, 30, 64, 115, 75, -22, -10, 123, 101, 66, 108, 48, -110, -71, 43, -108, 4, 18, 64, -111, 35, -30, -106, -48, -80, -95, -1, 88, -34, 28, 114, -42, -61, -113, 46, 119, -72, -77, -8, 6, 20, 96, -122, -49, 73, -92, -8, -27, 30, -68, -45, -1, -51, -98, 76, -71, -62, -41, 88, -55, -79, 15, 11, -7, 107, -13, -128, 112, 115, -77, -96, -93, -66, 1, 31, -53, -108, 47, 5, -97, 34, -117, -98, 15, -37, -24, -110, 33, 26, 97, 18, -71, -12, -53, 65, 16, -102, 53, -27, 8, -18, 114, 51, -77, -74, 11, 34, -114, 87, -30, 110, -127, -88, 78, -83, 86, -106, 8, 20, 10, 31, -71, 30, 56, 34, -17, -21, 56, -127, -78, 116, 47, -95, -48, -97, -3, 121, -93, -98, 55, -29, 100, 92, -96, 52, 72, -52, -35, 88, -39, -25, -54, -102, -19, 88, 22, 92, -54, 5, 55, -117, -17, 76, -110, 1, 35, -34, 14, 42, -126, 89, 77, -101, 38, -13, 53, 123, 1, 96, -68, 78, 21, -31, 64, -27, 93, 126, 112, 56, 85, -111, -112, 4, -61, 90, 99, 24, -31, -87, 75, 41, 82, 99, -84, -39, 99, -96, 27, -102, -9, 3, 25, 87, 1, 59, -104, -3, 82, -106, -87, 53, -59, 87, -53, -49, -99, -100, 51, 87, -22, 40, 28, -29, 125, -50, -127, -112, -24, 58, 7, -97, -105, -124, -23, 110, 3, -1, 103, -76, 124, -12, 56, 81, 55, 115, 68, -98, -14, -57, 70, -16, 103, -54, -21, -84, -35, -35, -35, -44, -74, -47, -9, -30, -106, 7, 59, -62, 38, -89, 120, 101, 63, -102, 105, 115, 22, -123, -125, -60, -119, 90, -69, 102, 60, 108, -29, 0, -12, -103, 48, -97, -69, -91, 22, -11, -118, -15, -79, 71, -106, -57, 80, 15, 87, 111, 9, -42, 18, 43, 22, 109, 117, -117, -17, -12, -113, -54, 125, 52, -82, 107, 25, 53, -125, -75, 34, 40, 96, -89, -104, -84, 3, -92, -64, -87, 127, -22, -93, 45, -6, -18, -117, 117, -104, 44, 106, -115, 53, -56, -98, -4, 30, -5, 122, -96, 32, 12, -104, 47, 22, -112, 68, -93, 5, 40, -35, 24, 84, 79, 114, -10, 82, -108, 39, -99, 42, -100, -99, 12, -27, 44, -127, -85, 56, 61, 116, 74, 53, 109, 53, -126, -14, -23, 98, 42, -14, 32, 27, -57, 6, 35, 61, 87, -36, -77, -124, -73, -15, 47, 62, -30, -113, 77, 62, 80, 22, -100, 26, -12, 122, -105, -77, 42, 20, 122, 13, -81, -66, -78, -11, -108, -72, -35, -23, -88, 64, -51, -46, -94, 19, 72, -44, 84, -109, 70, -68, -2, 18, -28, -114, -97, -25, 86, -21, 78, 57, 100, 66, 125, 44, 20, 94, 110, 68, -109, 121, -88, -72, 23, -36, -57, 99, 61, -60, 92, -75, 30, -101, -91, -126, -122, 125, -89, 65, -63, 76, 88, 58, 33, -90, 89, -128, -117, 120, 99, 64, 60, -18, -4, 58, -118, 109, 58, -13, 16, -113, 53, 39, -49, 124, 78, -94, 25, 4, 75, 53, -82, -10, -124, -94, 60, 96, 34, -89, -93, 2, 6, -49, -32, 39, 78, 48, -122, 42, 44, 40, -41, 91, -29, 125, -50, -8, 89, -69, -73, -1, 73, 112, -71, -64, -46, -29, -27, -43, -80, -6, -22, -112, -40, -22, 81, 60, 17, -65, 113, -92, -102, -33, -102, -16, -45, 28, -59, -127, -67, 32, -20, -91, 93, -50, 36, -30, 57, -99, -80, -111, -110, 105, 123, 95, -111, 57, -115, -62, -85, 17, -25, -51, 45, 50, -108, -112, 39, -56, -13, -83, 75, 74, 65, 114, -32, 56, -40, -26, -48, -59, -36, -72, -71, -118, 21, 38, 112, -108, 123, -46, 80, 73, -72, -23, 80, -128, 64, -128, 76, -111, -17, -51, 108, -127, -72, 120, 95, 53, 91, 91, -29, -29, -2, 118, 43, 29, -10, 31, -84, 65, -34, 95, -127, -12, 107, 43, -21, -119, -55, 3, 38, 29, 53, 33, 0, 101, -77, 45, 39, -115, 21, -102, 108, 3, -39, 116, -75, 14, 42, 106, -58, -68, -112, -2, -67, -36, 19, -30, 24, 15, 78, -72, -24, 104, 60, 58, -16, -57, -27, -10, -16, -54, 109, 40, 126, -126, -13, -75, 91, 91, 107, -86, 7, 51, 7, -117, -96, 57, 103, 64, 97, -42, -80, 63, -77, 15, 53, -96, -96, 64, 83, -90, 80, -41, 71, -70, -71, -84, 93, -9, -24, -74, 117, -102, 4, 98, -93, 125, -71, 92, -77, 118, -47, -55, -31, -96, 102, -7, 3, 48, -108, -88, -47, 105, 101, 15, -72, 58, -50, -52, -77, -125, 18, -67, -95, 31, 108, -91, -28, -17, 95, -81, -35, -85, 69, 126, -126, -73, 60, 58, 38, -35, -30, 91, 127, -30, 90, 53, -38, 54, 36, -91, 55, 89, -11, -68, 110, 125, -127, 58, -90, 80, 102, -45, 103, -27, -109, -126, 86, -95, 12, 93, 34, 123, -88, -17, 92, -29, -54, 14, 82, 59, -42, -117, -102, -39, -29, 64, 95, 101, 48, -9, -30, 92, -108, -105, 110, -99, -91, -16, 69, -44, -91, -51, 33, 6, -103, 73, 31, -90, 73, 110, -66, 120, -110, 75, 81, -22, -9, -105, 38, -45, -60, -52, -83, 67, -80, 11, 127, 3, -84, 108, 119, 34, -56, 126, -52, 90, 51, -71, 51, -92, 120, 18, -57, 55, -98, 84, 81, -41, -108, -76, 58, 52, -26, 77, -3, 127, -53, 100, 20, 28, 18, 59, -87, -40, -23, -100, -48, -128, -9, 89, -6, 32, -50, -17, -52, -113, 83, -1, -1, 86, 35, -59, -93, -86, -82, -61, 19, -88, -61, -100, -33, -6, 102, 94, -115, 19, 108, 97, -102, 95, -7, 27, 40, -79, -38, 106, -22, -21, -114, -112, -32, -84, -46, 60, 54, 71, 55, -81, 99, 89, -46, 75, -15, 8, -64, -69, 100, 6, -35, -52, 93, 116, 118, 81, 20, -50, -3, -77, -73, -71, -100, -121, -75, 60, -53, -70, 69, 91, 10, -56, -15, 79, 17, 96, 98, -26, 19, 50, -122, -122, -30, 3, -31, -30, 109, -16, 125, 25, 108, -121, -128, -87, -102, -52, 90, 94, 3, -11, -101, -93, -122, 65, -122, -91, 41, 103, -26, -20, 125, -61, 24, -10, 109, 112, 113, -84, 93, -5, 48, -79, -84, 35, -113, 4, -109, 21, 16, -110, 36, -105, 73, -70, -53, 121, -44, 4, -82, 117, 86, 91, 0, 100, 5, 109, 97, -84, -14, 66, 111, -128, -90, 23, -58, 46, -7, 29, 84, -30, -124, 112, -39, -65, -66, -54, -36, -34, -40, -7, -123, -111, 103, -39, 106, -71, 41, 84, 64, -83, 64, 85, 46, -109, -77, -23, -63, -98, 82, -72, -10, 120, -82, 121, 103, 0, -29, -42, 64, -94, -15, 13, -94, -85, 106, -97, -97, 39, -115, -66, 12, -78, -76, 116, 96, -55, 114, -87, -70, -88, 93, -55, 108, 108, -97, -75, 45, -88, -128, 99, -71, 11, 116, 2, -114, 15, -112, 104, 94, -98, 19, -120, -48, -103, 59, -117, -125, -53, 121, -81, 98, 112, 78, -55, -34, 63, -86, -113, 90, -67, -81, 107, -54, 50, 119, -24, -121, -73, 82, -95, 100, -110, -92, -75, 80, -94, 29, -122, -75, 33, -45, 39, -83, 25, 23, 46, -127, 58, -81, 22, -81, -30, 32, 0, 38, -103, -88, 61, -51, 80, -94, 80, -76, -45, -62, 89, 76, -94, 76, -10, 77, 60, -29, 105, -75, 38, 11, -39, 119, 32, 98, -128, 22, -36, 66, 5, 111, 127, 59, -93, 35, -5, 82, 53, 122, -36, -26, -13, 2, -41, -109, -72, -113, -3, -105, 57, -61, -90, 12, -88, 41, -105, -78, -120, -21, -12, 90, -54, -121, 11, -115, -94, -76, -46, -57, 19, -39, 56, 41, 125, 77, 86, -36, -118, -108, -101, -112, 40, -68, -125, 39, -88, -11, -50, -87, -77, -34, -6, -51, 58, 40, 50, 62, 87, -117, 115, 70, 95, -104, -32, -12, 54, 17, -67, 35, -28, 113, -26, 8, -53, 33, 84, -22, 31, -70, -86, 105, -70, 80, -27, 76, -11, 48, -116, 77, -61, -113, 73, 27, -4, -33, -6, 66, 78, -67, 70, 84, 69, 35, 124, -79, 74, 26, -114, -27, 85, 43, 80, 36, -77, 102, -75, 29, 88, 119, 119, 98, -118, 116, -65, 86, -97, 55, 3, -35, 125, 124, 89, -2, 109, -65, 113, -80, 59, -76, 1, 110, -33, -60, -72, -47, -5, -3, -9, 85, 19, -11, 79, -111, 110, 32, 70, 34, -107, 85, 44, -25, -73, -16, 75, -59, -108, -84, 126, 77, 126, 116, 38, -1, 92, 55, 10, 48, 113, 10, 108, 70, 103, -29, -97, -103, -32, -108, -8, -48, -12, -17, 50, 94, 31, -25, -2, 74, -70, 28, 17, -4, -3, -29, 22, 126, -99, -17, 50, -82, -58, 81, 75, -128, -39, 0, -41, 12, 53, 28, 28, 125, 10, -33, -35, -65, 80, -41, 56, 97, 92, -8, 93, -29, 62, -59, -89, 26, 99, 121, -1, 68, 34, 10, 67, 15, 12, -12, -84, -102, 28, 41, -7, -33, 32, 119, 65, -14, -112, -28, 7, 34, 124, -86, 10, -34, 112, 41, 86, 96, -74, -105, 104, -75, 78, -78, -44, 115, -125, -100, 68, 94, 98, 40, 118, 21, -116, -79, 8, 124, -88, -39, 66, -68, 14, 46, -9, -59, -106, -69, 59, -82, 59, 98, -41, -51, -106, -103, 66, -115, -50, -59, -55, -26, 3, -43, -86, 54, 99, -65, -85, -32, 124, 24, -73, 11, 3, 108, 55, -57, -81, -39, 71, 49, -53, -38, 19, 85, -6, -48, 114, -66, -47, -29, 62, -28, -127, 72, 34, 61, 10, 42, -29, 45, 91, 79, -78, 0, 9, -46, 63, 104, -46, -10, 71, 47, 40, 83, -47, 57, -62, 21, 10, -95, -26, 27, 91, 59, -66, 40, 36, 33, 114, 125, -81, -124, 8, -60, 100, -36, 6, 68, -114, -71, 68, 87, -108, -33, -17, -86, -44, 45, -97, 99, 95, 65, 39, 114, 41, 56, -71, 102, -83, 82, -33, -102, -100, -37, 29, -53, 51, -3, 79, -77, 103, -17, -26, -5, -102, 57, 8, -26, 34, 106, -65, 5, 52, -78, 116, -66, -64, 45, -68, -85, -35, 83, 37, 88, 95, -5, 51, -89, -52, 90, -109, 3, -123, -56, -9, 31, -125, -99, 14, -32, 98, 28, 47, 11, -114, 53, 1, 57, 54, -72, 122, -53, 102, -7, -89, -27, 14, -76, 20, 83, 84, -58, -89, -78, 110, -28, -110, 123, -67, 61, -7, 27, -103, 24, 45, 76, -77, 40, 116, -103, -116, 75, -39, 97, -96, -65, 119, 124, 7, -33, -128, -74, 93, 95, 58, 16, 45, 0, -43, 105, -109, 34, -74, -106, 12, 2, -117, 122, -13, -106, 8, 74, -106, -3, 9, -30, -50, 27, -30, -117, -122, 9, -45, 64, 122, 67, 40, 85, -110, -126, 78, 30, -55, 117, 110, -15, 47, -26, 107, 109, 48, 101, 94, -79, -117, 28, -50, 74, 123, -128, 27, -107, 49, 63, 98, -124, -81, 46, 124, -106, -78, -77, -103, -117, 47, -36, 30, 93, -6, -89, -93, 46, 124, 96, -125, 39, -120, -91, -31, 111, -11, -31, -82, -87, 30, 42, 73, 87, -44, 65, -112, -56, 86, 36, 18, -106, -58, 26, 20, -27, 88, 57, -18, -86, 7, -106, 50, -7, -55, -13, 104, 98, 97, 36, -26, -19, 84, -19, -99, 113, -58, 29, -124, -1, -108, 90, -24, 6, 46, 40, 13, -112, 110, -57, 5, 96, -76, 19, 111, -78, -31, 98, -74, -2, -76, -53, -11, 12, 77, 95, -30, 36, -56, 1, -15, -90, -85, 101, -7, 76, 25, -67, 90, 101, -21, 3, -64, 40, 58, 1, 104, -3, -79, -34, 102, 40, 10, -86, -45, 100, -92, 104, 29, -74, -80, -7, 101, -77, 31, -76, -64, -32, 70, -108, -25, 34, -15, 4, 47, 43, -44, -100, -27, -75, -103, 119, -71, 25, 60, -77, 52, -21, -108, -82, 47, -62, 123, 95, 113, -32, 118, -90, 47, -50, -64, 91, 76, -91, 55, 121, -115, -11, 61, 101, -21, 89, 54, -57, 15, -59, -4, -98, -34, -95, 40, -64, -54, 99, -128, 82, -34, -14, 19, -127, -17, -111, -104, -103, -21, 56, 66, -64, -116, 91, -120, 64, -94, -40, -61, 50, -92, 70, -125, -13, -47, 100, -64, 27, 10, 87, -75, -72, -20, 94, 125, -4, -55, 89, -26, 15, 43, -20, 17, -49, -59, 46, 94, -127, -71, -98, -84, 122, -76, 96, -70, 118, -99, 53, 6, -121, -82, -75, 22, -85, -25, -119, -43, -86, 98, 115, 53, -108, -96, 37, 22, -27, -38, -118, -68, -41, -114, 37, -70, 85, -73, 9, 114, -101, -58, -114, -97, 91, -33, 51, 58, -32, 5, 90, -22, -83, 68, 110, -84, -96, -104, 7, -123, -103, 22, -42, -27, 40, -8, 8, 46, 14, -46, -23, 79, -122, 92, 34, 21, -58, 35, -12, -92, 76, -78, 62, -30, 89, -52, -118, -106, -95, -11, -45, -75, -63, 65, 92, -76, 18, -9, -38, -97, 91, 123, -16, 106, -10, 89, 126, -81, -125, 109, -80, -115, 63, 40, 91, 16, -35, 31, 12, 108, 61, 37, 19, 14, -33, -94, 31, -100, -101, -86, -72, 23, -40, -46, 6, -123, -100, 17, -62, 22, 10, 93, 87, -115, -10, 115, 114, -112, -102, -65, -120, -44, 28, 112, 56, -82, 22, -84, 124, -117, 19, -29, 120, -25, -107, -62, 13, -13, 126, -2, -93, -25, 55, -48, 101, -106, 123, -4, 12, 56, 119, 73, 93, -122, -73, 21, 75, 49, -87, 49, 116, 76, -32, -96, -109, -30, -93, -122, 67, -66, 57, 97, -27, 7, 127, 110, 121, -5, 118, 116, -127, -53, -50, -94, -100, -67, -79, 66, -88, 80, 16, -121, -79, -110, 68, -126, -97, -50, -28, 33, -103, -30, -60, -57, -119, -3, -101, -118, 75, 37, 91, 91, -87, -116, 32, 78, -2, -12, 86, 11, 114, -64, 68, -85, 22, -26, 64, -31, -72, 64, -45, -87, -83, -44, 55, 31, 21, -37, 86, -77, -58, 4, -9, -78, 68, 12, 5, -95, 50, -35, -15, -80, 56, 79, 27, -91, -30, 33, 120, -47, 101, 76, -80, 43, 55, 27, -3, 116, -76, -52, -124, 74, 125, 14, -85, 78, -39, 92, 47, -98, -38, 12, -36, -37, 125, 125, 58, -121, 34, 116, 30, -54, 31, 90, 70, 89, 87, 69, 17, 88, 1, 86, -19, 127, 111, 14, -30, -93, -114, -74, -105, 58, -74, 82, -102, -49, 78, -38, 91, 0, -24, -10, 0, 125, 110, -47, -97, 40, -10, 108, -101, -76, -2, 5, 57, 49, 80, 112, 91, 112, 66, 110, -99, -31, 52, -27, 12, 5, 1, -33, -70, 17, -52, -107, 7, -76, -28, -110, 70, 45, -89, -42, -55, -77, -2, 99, -7, 21, 8, 64, -92, -41, 95, -54, -102, -57, 113, -73, -71, 116, -68, -127, 119, -95, -72, -99, -36, -45, 67, -60, -128, -128, 36, 22, 5, -104, 95, -89, 45, -21, 78, 25, 9, 18, 123, 97, -46, 36, 69, -65, 49, 14, 77, 45, 21, 64, -11, -64, -113, 63, -73, -99, -10, 9, 35, 35, -24, -107, 98, -50, 51, 44, -103, -30, 26, -92, 58, 108, -61, 21, 52, 8, -28, 70, 124, -84, 8, -68, 104, -42, 55, -74, -34, 97, 74, -54, -98, -15, -92, 68, 118, 11, -111, 14, 6, 6, 58, 111, -8, 69, -118, 77, -76, -121, 12, 12, 107, 75, -31, -27, 10, 120, -6, 34, -123, 70, 85, -55, -109, -86, -17, 75, -14, -82, 41, -13, -38, -92, -106, -45, 27, 80, 15, -7, -103, -66, 108, 61, 77, 111, 106, 34, -78, -113, -91, -87, -62, -54, 25, 11, -2, 121, -58, 7, 29, -34, -127, 44, -51, 99, -51, 69, 71, 84, -29, -2, -60, -84, -125, -38, -59, 111, -64, -23, 88, -76, -46, 109, -101, -117, -61, -104, -127, -88, -86, -77, -30, 54, -124, -71, 15, 127, 36, 28, -101, 70, -89, -34, -32, -74, -64, 111, 86, 126, -108, -101, 119, -112, -13, 66, -78, -20, 27, 41, -100, -9, 52, -33, 90, 98, -40, -18, 5, -26, -17, -56, 127, -56, 4, 83, -122, -42, 32, -56, 42, -107, 29, -38, -88, -44, -44, -107, 47, -9, -101, 64, 81, 38, 108, 115, -84, -128, -63, -115, -93, -47, -47, -37, 101, 21, -78, 103, 64, 98, -7, -101, 93, 62, -23, -117, -76, -96, -83, 20, 65, 52, -87, -107, -113, 23, -73, 66, 52, -46, 15, -76, 4, -107, 111, -95, 49, 68, 23, -28, -47, -96, 31, -35, -35, 120, 66, 52, 37, 8, 69, 111, 55, -109, -105, 43, 62, 70, -9, -7, -46, -73, 112, 102, 2, 41, -49, 21, 63, -51, -57, 91, 35, 110, 99, 11, -116, -105, 99, -113, 50, 25, 66, 69, 62, -79, 28, 55, 82, 12, 111, -50, 3, 114, -70, -47, 90, 43, 109, -47, -20, -64, -67, 66, 14, -18, 35, -49, 116, 119, 86, -62, -87, 12, 13, -121, 21, 5, 89, 6, 82, -110, -101, -11, -84, -60, -43, -16, -17, 85, 5, 105, -19, 37, 15, -40, -109, -58, 122, -37, -97, 5, 102, 33, -112, 45, 37, -118, 15, 50, -105, -114, -48, -68, 33, 34, -79, 63, 63, 30, 117, -68, -95, 77, -38, 6, 18, -86, 83, -59, -20, 125, 64, 90, 55, -60, 109, 113, 5, 66, -82, -12, 4, -113, -13, 20, 36, -108, 126, 113, 0, -80, 34, -113, -29, 13, 37, 116, -30, -82, -38, -88, -107, -3, 8, -50, 8, -96, 121, 62, -110, 20, 63, -119, 33, 65, 121, 79, -71, 91, 83, 118, -64, -127, -13, -36, -21, -88, -12, 54, -33, 75, 83, -121, 60, -60, 110, 127, -119, 83, 87, -20, -33, -4, 100, -34, 114, -31, 118, 28, 91, 87, -33, 77, -54, -28, 15, -88, -46, -89, -56, 47, -7, -103, -47, -126, 43, -78, -1, 114, 14, 46, 84, 59, 62, -31, 66, -10, 12, -69, -51, 55, -80, 53, 18, 95, -47, 52, -40, -121, -21, 66, -92, -50, 70, 105, 116, 20, -5, 95, 23, -64, 28, 48, -80, -46, -34, -86, -87, -70, -10, -86, 87, -100, 71, 122, -5, 89, 57, 126, 96, -115, -77, 94, 33, -24, -27, -103, -2, 124, -74, -127, 45, 58, -106, -43, 29, -45, -100, 119, -106, 86, -122, 111, 40, 116, -110, 16, -11, 77, 102, -44, 43, -16, 72, -94, -22, -23, -70, 17, 38, -31, 45, -62, -4, 120, -50, -108, 57, 80, -44, -52, 23, 127, -119, 97, -47, 97, 122, 127, 30, 122, 117, 6, 96, 45, -120, -19, -67, 5, 30, 0, 92, 0, 31, 64, 111, -30, -49, -93, 109, 25, 124, -49, -83, -116, -79, 21, 124, -63, -103, -85, -55, -18, -25, 48, 88, -51, 51, -35, 11, -72, 85, 95, -56, -49, -33, -98, -2, -2, 22, 100, -45, -84, 27, 15, -9, 81, 77, -82, -9, 40, -59, -2, 60, -44, 36, -38, -11, 7, -57, 73, -23, -106, -109, -52, 103, 28, -74, 107, 54, -60, -99, 21, -56, 34, 20, -41, 61, 99, 46, 40, 30, -75, -101, 105, -79, -55, 70, 115, 90, 1, -119, 23, -94, -64, -41, 81, -3, -112, 26, -51, 112, -73, 8, -5, 9, -99, 123, 58, 34, 11, -76, -57, -124, -100, 39, 56, -33, -83, 110, 124, -5, 100, -69, -49, -92, 124, 79, 49, 37, 7, -78, 94, -65, 94, -43, 28, -74, -82, -121, -28, 88, -62, 7, 117, 115, 82, -41, -2, 40, 96, 51, 118, 17, -16, 0, 38, 84, -50, 74, -93, -100, 32, -105, -88, 81, 107, 11, -109, -67, -118, -124, 18, -37, 79, -48, 111, 104, -48, -53, -125, -90, 8, -111, -34, 80, -50, 47, 18, -114, -11, -37, -74, 59, -118, 111, -7, 48, 92, -59, -28, 27, 108, 106, 57, 121, 124, -100, 32, -102, 90, 67, -106, -89, -91, 113, 92, 106, 3, 38, -96, -19, 105, -47, 114, 81, -61, -62, -43, -127, -59, -6, 39, -7, 110, -72, 41, 21, -94, -43, -25, -45, 32, -8, -69, 66, 69, 121, 7, -127, 18, -8, 23, -56, -121, -18, 57, -93, 88, 60, 110, 87, -5, -112, -48, 22, 115, 52, 94, -73, -100, 83, -111, -110, -53, -44, 93, 88, -3, 31, 120, -44, 90, -72, -124, 86, 48, 5, 77, 124, 46, -110, -62, -43, 92, -42, -73, 47, -116, 85, -67, 94, -5, -119, 99, -95, -29, -79, 58, 115, -95, -102, 65, -63, 73, -81, 68, -73, 110, -111, 7, 9, -109, 18, 30, -2, 1, 69, -25, -75, -116, -68, -113, -55, 34, 62, -124, -44, -14, -53, -100, -119, -96, 85, 70, -122, 72, -58, 1, -13, 0, -122, -8, 111, -107, -72, 31, -128, -26, -10, -106, 67, -24, -103, -87, -22, 11, 93, 54, 84, 118, -91, -85, 93, 115, 39, 111, -99, 43, 19, 90, 4, 63, -40, 53, -50, 57, 17, 68, -67, 103, -85, 100, 6, 103, 45, 40, -115, 9, 91, 3, -49, 69, 117, -101, 14, 7, 86, 90, -3, 111, -45, -3, 74, 118, 52, -87, 91, -116, -81, -12, 74, 25, -95, 95, 48, 102, 59, 26, -38, 102, 15, 21, 117, -114, 52, 68, 20, 21, -75, -70, 71, -84, 92, -126, -93, 35, 8, 3, -99, 52, 112, -96, 69, 92, 88, 5, -43, -19, 119, -33, -121, -128, -64, 57, -120, -35, 72, 38, 30, 111, 101, -83, -100, -65, -103, 42, -23, 116, -43, -17, -98, -1, 76, 33, -35, -126, -32, -32, 17, -11, -47, 101, -15, -38, -21, 21, 7, -79, -66, -90, 121, 121, 49, 4, 41, -50, 36, -109, -62, 42, 37, -61, -100, 36, 38, -30, -77, -23, -67, -93, -80, -57, 82, -5, -31, -103, -65, 29, -108, 38, -113, 12, 78, -30, 99, -33, -24, -8, 39, -43, -100, 32, 36, -32, -85, -112, 44, -77, 113, -78, 49, -71, 127, 2, 110, 49, -106, 34, 92, -9, 46, -122, 68, -92, 77, 40, 107, -116, 102, -40, -79, 103, -105, 44, -45, -109, -51, -114, -63, 92, 6, 120, -80, -63, 15, 127, 45, -98, -92, -68, 66, -125, 44, 4, 12, 26, -57, -98, -38, -115, 43, -21, -27, 72, 66, -26, 3, 66, 32, -50, -84, -64, 30, 117, 124, 67, -105, -126, -109, -8, -93, -77, -96, -100, -1, 85, -62, -13, -59, -7, 120, 94, -62, 75, -31, -79, 47, 98, -98, -59, -9, -38, -78, 62, 126, 92, -2, 84, 49, 3, -31, 47, 88, 0, 76, 113, -58, 38, -28, -121, 52, -2, -24, 31, -117, 97, -111, -86, 5, -6, 50, -11, -24, 24, 72, 81, -72, 82, 87, -22, -75, 14, 84, -122, -5, -44, -67, -35, -68, 5, -7, 57, -70, -43, 104, -39, 23, -59, 89, -36, 11, -32, 70, 75, 10, 114, 120, 118, -79, -124, 76, -35, -67, -58, -38, 110, 1, 24, 95, 125, 26, 48, -31, -128, -24, 2, -19, -124, 6, -61, -5, 37, -11, -72, 117, -61, -53, 62, 98, -94, 50, 17, -88, -28, 114, 21, 96, 14, -5, -13, -6, 25, -16, 122, 100, 10, 116, -29, -3, 79, 0, -39, -90, 101, 120, -47, 10, 103, 2, -122, -116, 82, 108, -96, -98, -76, 119, -32, 56, -118, -47, 4, 76, 84, -8, 114, -114, 93, -39, 59, -78, 92, 119, 15, -67, -32, -107, -95, 23, 80, -18, -40, -50, 40, -36, 75, -4, -100, 54, 106, -111, -15, 24, -110, 48, -33, -13, -80, -31, 113, 79, 126, 52, 114, -40, -58, -18, -22, 100, 8, 84, 50, 22, -40, 73, 32, -113, 107, 30, 41, 50, 54, -107, 41, -70, -11, 68, -50, 80, -103, 43, 110, -99, 15, 42, 119, 11, -66, 7, -88, 58, 101, -85, -112, -108, -14, -84, -16, -48, -10, 85, -13, 88, 92, 108, 71, -128, -23, -64, 104, -71, -79, 23, -61, 15, 125, -117, 41, 66, -90, 28, -62, -24, 89, 106, 96, 19, -41, -34, 22, 60, 88, -64, -20, 94, 100, 111, -62, 68, 22, 21, 126, -123, 22, -127, -71, 11, 76, -119, 92, 81, -6, -63, 60, 42, -14, 12, 74, -72, -4, 24, -40, 69, -113, -123, -98, 81, -80, 103, -119, 127, 125, 87, -39, 103, 7, -3, 108, -63, 91, -112, 85, -88, -69, 24, 46, -50, 65, -54, 117, -14, 47, -17, 86, 97, 69, 64, 34, -41, -14, 51, 98, 44, 126, -97, 92, -35, -34, -118, -121, -18, -22, -124, -57, -108, -83, 78, -51, -78, 21, -112, 97, 121, 125, -80, 73, 47, -62, 60, -113, -84, -8, -28, 87, 83, 21, -36, -109, -12, -110, 31, 19, 16, -54, 115, 20, 124, 10, 18, -96, -66, 119, 40, 120, -128, 86, -28, -51, 9, -98, 119, -37, 43, 81, -74, -15, -53, 42, -97, 70, 92, 72, -60, 73, -8, -51, -23, 35, -88, -37, 120, -105, 81, -75, 108, 67, -17, -128, 109, 101, 59, 38, 24, -48, -16, 21, -30, -69, -83, 24, 118, 92, -114, 60, -11, -17, -65, 17, -46, 97, -82, 91, -74, 52, -9, -67, 31, -115, -37, -108, 48, 30, 28, -76, 15, 27, -107, 97, 91, 83, 37, 25, -123, -53, -105, 122, 21, 96, -22, -46, -13, -109, 21, -33, 62, 6, -92, 95, 49, 71, 49, 90, 99, 127, -64, -105, -128, 29, -41, 48, -25, -21, -20, -99, -109, 92, 4, -89, -59, -111, -109, -72, -85, 87, 49, -15, -123, 84, -32, 7, -38, 70, 86, -85, -9, 33, 54, -57, -56, -39, 48, -123, 126, 52, -96, 51, -104, -23, -95, 71, 27, -6, -97, 103, -124, 43, -42, 54, 15, -23, 115, 85, 39, -3, -76, 31, 121, 18, 65, 123, 4, 60, -40, 68, -1, 67, 11, -90, 23, -16, -73, -97, 24, -121, 96, 0, 55, 114, -117, 93, -62, -18, 79, -114, -63, -22, 45, 12, -60, 46, 86, 94, 71, 21, -30, -19, 95, -88, 125, -95, 15, -42, 89, 68, 63, 85, 48, 109, -109, -72, 43, 6, 127, -59, 7, 67, -118, -55, -78, 110, -77, -77, -33, 13, -105, 54, 40, -59, 75, -113, 42, -55, 16, 104, -55, -115, 60, -55, 40, -10, -128, -83, 117, -12, -69, -83, -88, 29, -19, 29, 70, -63, 63, -11, -16, -48, 59, 26, 72, 111, 72, 114, -19, 107, -90, 43, -111, -111, -26, -84, 23, 107, 29, 65, 105, -21, -75, 70, -81, -83, 125, 15, -92, 120, -125, -102, 95, -2, -46, -39, 89, 97, -119, 85, 16, -126, -92, -17, -97, 82, 104, 21, 117, 25, 91, 6, 38, -24, 48, 84, 35, 77, -93, -47, -105, 77, 62, -41, -99, -103, 68, 85, -37, -90, -65, 107, -109, -20, -124, 43, -52, -120, -116, 109, -81, -3, -115, -24, 40, -31, 55, 14, 25, 31, -107, 112, 46, -56, -61, -92, -103, 99, 43, -26, -38, 42, 9, -76, 62, 10, -11, 73, -12, -83, 19, -73, 5, -23, 83, 48, 10, -52, 10, -77, -99, -107, -10, 103, 62, 95, -16, 63, 45, -26, -113, -39, 47, 111, -16, 18, 5, -36, 104, -36, -17, -29, 27, 60, 125, 57, 20, -25, 110, 124, 19, -45, -69, -96, -78, -121, 66, -95, 120, 13, 106, -101, 78, -4, 77, -22, 50, -56, 57, -94, -21, -2, -90, 105, -74, 26, -6, 112, -79, -14, 20, 115, 38, 86, 27, -123, 87, 25, 45, 2, -85, 109, 33, 40, 125, 70, -67, 46, -65, 42, -4, 33, -1, 116, 29, -52, 20, 120, 10, -50, -44, -68, -115, -113, 3, -111, -1, -70, -52, -57, -28, -6, -34, 15, 0, -122, 58, 61, 116, -46, -81, -81, -118, -41, 30, 60, -97, -92, 78, -17, -50, -14, 78, 125, -14, 10, -75, 47, -60, 30, -128, 16, 34, 75, 37, -79, -15, -20, 24, -98, 69, -7, -44, 103, 31, -6, -89, 126, 25, 96, 72, 122, -101, -109, 52, -36, -88, -118, 35, 118, -127, -58, -47, -94, 42, 31, 73, 86, -103, 58, -64, -56, 22, -13, 16, 44, 35, -123, 96, -36, -4, 27, 15, -41, -86, -11, -41, 19, -37, -121, 69, 25, 87, -124, -17, -83, -95, -121, -8, 117, 36, 102, -37, 35, 105, -3, -18, -20, 40, -72, -96, -66, -86, -83, -90, -82, -40, 10, -48, 93, -70, -81, 3, 28, 62, 113, 48, 100, 87, 37, 82, -68, 106, 74, 10, 17, -19, -108, -32, -36, -120, 63, -116, -17, 65, -75, -29, 81, 83, -77, 52, -24, -43, 31, 45, 52, 108, 34, -70, 122, 118, -101, 18, -114, -50, -99, 2, 32, -103, -99, -127, -21, 44, -65, 83, -73, -105, 14, 96, -50, 115, 106, 101, 78, 115, 60, 56, 55, -106, -114, -52, -127, 80, 53, 95, -124, 45, -24, 23, 100, -18, -32, 89, -91, 74, -67, 21, 64, -98, -26, 70, -43, 69, 78, -54, -38, -121, 111, -30, 21, 3, -81, 11, 94, -119, 70, -60, 89, 13, 7, -20, -99, -73, -108, 4, 118, 118, 16, -13, 2, -47, -97, 24, 127, -115, 40, -109, 68, -85, 62, 42, -4, 19, 116, -4, -34, 81, -91, -39, -124, 86, 33, -98, -98, -83, 33, -29, -98, 62, -49, 14, -65, -44, -21, 72, -70, -81, 2, -25, 1, 35, 8, 15, -94, -99, -117, -89, 94, 3, -111, 30, 1, -21, 96, -119, 2, 17, 86, -107, -114, -84, 46, -95, -29, 91, -113, 61, -46, -21, -74, -75, -12, 49, 17, 4, -101, 14, -80, -1, 14, 77, -127, -107, -115, 66, 120, -126, -89, -123, -3, 47, 113, -87, -38, 108, 69, -19, -61, 6, -95, -83, -85, -30, -29, 29, 113, -45, 85, -105, -45, -83, 100, -23, -66, 52, 54, -16, 89, 93, 127, 17, -44, -63, -128, -110, 73, 12, 58, -58, 56, 49, 25, 114, -105, 7, -48, -106, -24, 9, -76, -24, 96, 122, 38, -49, 80, -12, -71, -12, -65, 113, -83, -106, -118, -101, -46, -68, -84, 71, -69, -8, -7, 93, -84, -77, 108, 36, 10, 35, 17, 36, 20, -40, -73, -18, -31, 80, 81, -104, 125, -34, 52, -34, 28, 5, -16, 22, 124, -70, 60, 36, 106, -42, -71, 78, -42, -113, -7, 86, -8, -102, 84, -46, -60, -28, 1, 82, -123, 42, -109, 111, 86, 118, -115, 20, 27, 66, 66, -128, 75, 53, -72, -114, 76, -48, 121, -8, -66, -44, 115, -86, 73, -74, -80, 72, -122, -73, -48, -35, 55, 64, -58, -34, 91, 52, -22, 30, -125, -32, -53, -46, -52, -18, -97, 75, 46, -13, 12, 66, -64, 36, -116, 98, -47, 25, 58, 57, 96, 7, -67, -101, 36, 95, 23, 10, -104, -110, -6, -54, 59, 70, -51, -98, -18, 62, -9, 65, -55, 105, -119, 6, -25, -41, -34, 24, 64, 105, 117, -37, 83, 78, -48, -11, 19, -62, -24, -77, -31, -6, 18, -39, -127, -2, 114, 108, 102, 117, -73, 42, -27, -12, -53, -38, 44, 40, 46, 0, -128, 84, -115, -109, 106, -40, -30, -127, 18, 2, 15, 9, 20, 82, 47, -41, -45, -123, 65, -100, -54, -13, -39, -88, 91, -49, -67, -63, -116, -74, -123, -97, 21, -26, 83, -123, 124, -4, -67, 59, -122, 78, 3, -118, 97, 39, 126, -28, 90, -60, -67, 68, -22, -17, -4, 57, 105, -89, -11, -68, 127, 49, 60, -47, -114, 107, 115, 84, -20, 36, 93, -90, 25, -28, -117, -90, 105, 33, 108, -57, 73, -82, -36, 56, 21, -54, -28, 78, 25, -44, -93, -77, -96, -114, -14, -99, -110, 111, -45, 7, -115, -7, -54, -77, -3, 111, 118, 4, -73, 49, 60, -31, -44, 43, -86, 86, -89, 48, -37, -70, 51, 34, -43, -113, 7, 122, 56, 31, -89, -38, 6, 60, 14, -105, 91, 49, 24, 44, -87, -99, 106, -37, 102, 72, -81, -107, -4, -116, -20, 46, 79, 73, -54, -100, -125, -75, 6, -99, 3, -35, 127, -109, -97, -38, -35, 37, -7, 28, -92, -79, 63, 88, 98, 87, -19, -102, -42, 41, 88, 46, -20, 29, 96, -86, -123, 70, -98, -77, -80, -126, 21, -16, 64, -20, 27, -16, -55, -55, -76, 117, 66, 7, -128, 18, -118, 18, -87, 29, -109, 3, -2, -29, -31, -28, -88, -18, 92, 34, 88, -73, 127, -120, -9, 84, -36, 76, -127, -125, 61, -107, -96, -49, -81, -108, 44, -19, -40, 117, -96, -42, 9, -68, -17, -98, 19, -69, 71, -70, 6, -68, 3, 81, -64, -59, 92, -32, 123, 2, -107, 125, 25, 25, -45, -56, 113, -13, 57, 7, -71, -32, 106, 9, 61, 111, 86, 18, 77, 85, -116, -106, 93, -124, 41, -83, 18, 87, 105, -2, -128, -58, -5, 82, 11, -49, -26, -126, -76, -93, 17, 74, -117, 26, 54, -1, 77, -118, -94, -12, -122, -54, -49, 115, -126, 118, -111, -49, -89, -13, 82, 47, -50, 50, 124, 65, 112, 19, -42, -26, -78, 80, -85, 51, -40, 58, -96, -109, 118, 12, 9, -100, 70, -124, -106, -75, 54, -100, 98, 77, 58, -46, 117, 81, -22, 75, -63, 37, 29, 118, 64, -3, 95, 47, -79, -57, -104, -75, -88, 15, 50, -57, 103, -13, -34, -43, 65, 51, 58, -49, -3, 48, -36, -8, -121, 9, 82, -26, -98, -7, 69, -58, 31, 27, 42, 3, 17, -22, 74, -34, 5, -72, -35, 3, 4, -53, 127, 23, -87, 125, 37, 74, 32, 86, 52, -65, 22, -88, 41, -10, 44, 119, 0, 62, 77, -33, 18, -9, -43, -87, -103, 15, 85, 126, 12, 33, 112, -106, -60, 121, 83, -19, -119, -16, -83, -103, 91, -59, -61, -77, 40, 49, -74, 126, 72, 101, 123, 55, 103, -126, -77, 95, 89, -41, 108, -58, 109, -119, 125, 113, -59, 123, -19, -16, -8, 65, -74, 47, -100, 58, 17, 23, -39, -85, -36, -126, -30, 75, 36, -40, -17, -30, -103, -63, -43, -86, -80, 114, -118, 113, -45, -102, 8, -114, -36, -94, 65, 47, -86, 61, -47, 74, 93, 77, -106, -32, 49, 75, 24, 10, -44, 106, -88, -73, 44, -118, 91, -124, 56, -83, -52, 24, -102, 110, -36, -7, -90, -22, 124, 29, -92, -121, 104, -37, -99, 111, -68, -55, -75, -61, 19, -95, -22, 1, 9, 109, 59, 32, 27, 104, -40, -106, 72, 72, 126, 9, 53, -114, -23, -25, -86, 62, -76, -121, 80, -92, 126, 10, 101, -47, 63, 17, 20, 22, -116, 24, 25, 119, 84, -19, -59, 18, 48, -79, 21, -85, -17, 65, 11, -73, 110, -78, 21, 72, 120, -88, 73, -12, -13, 5, -58, 105, 2, 45, -10, -43, -106, -64, 51, -35, -102, -2, 93, 95, 52, -78, -110, 59, 122, -3, 101, 109, -20, -28, 25, 70, -128, -66, -17, 29, 105, -24, 87, -24, 80, 93, 127, 54, 14, 72, 39, -124, 29, 47, 24, 115, 102, -48, 73, -8, 73, -128, -74, 2, 36, -70, 0, -122, -97, 83, 60, -73, -103, -70, -69, -12, 105, -31, -100, -86, -29, 103, 105, 123, -111, -60, -43, 20, -64, 97, 87, -96, 59, -19, -46, -3, -99, -96, -29, 127, -45, 52, 107, -71, 91, 9, -121, -44, -4, 23, 121, -62, 115, 23, 99, -85, 91, -11, 30, 51, 105, -98, -32, 106, -23, 76, 17, -29, -84, -103, -87, -94, -12, 67, -42, -122, 16, 25, 109, 107, 123, -126, 15, -20, 77, 97, 23, -17, 127, 93, -109, -93, -89, -89, -107, -52, -12, 28, 45, 43, -45, -38, 15, -83, -31, 15, -21, 35, 107, 119, 94, 29, -103, 125, -10, 90, 98, 80, 54, 120, 96, 71, 85, 27, -75, -71, -117, -23, -26, 42, 31, 64, 31, 1, -115, -14, -7, -44, -127, 42, -105, -127, -111, 127, -96, 72, -50, 117, 31, 101, 113, -37, -5, -52, 127, -57, -126, 63, 44, 38, 6, 101, 89, -42, -113, -30, 55, 94, 57, -27, 76, 58, 7, 19, -51, -45, -1, 75, 98, -27, 103, -80, -66, 70, 93, -77, -8, -92, 91, -69, 23, 64, -33, 40, 126, -65, 95, -90, -20, -38, 49, -98, 32, -31, -10, 63, -25, -119, -89, -121, -4, 50, -27, -112, 68, 126, 34, 102, -24, 50, -16, 28, 53, -98, 103, 108, -81, -127, 107, 60, 57, -56, -21, -84, -2, 29, -124, -108, -118, -23, 22, -123, -17, 56, -62, 73, -4, 104, -20, 69, 57, 44, 56, 114, 98, 34, -96, -109, 60, 47, -5, 49, -31, 0, -46, -105, -34, 33, -22, 33, 25, -101, 103, 22, -37, 4, 76, 26, 61, 26, -19, -91, -63, 38, -127, 28, -103, 59, 56, -34, -15, -98, 6, -5, -120, 54, 40, -35, 42, 10, -9, 121, -54, -23, -55, -75, -24, -96, -86, -115, -80, 98, 23, 1, 16, 1, 8, -128, -24, 18, 37, -96, -98, -45, 118, 103, 44, -82, 82, 105, -26, -32, -11, -29, 56, -15, 5, -62, -52, 35, 1, 86, 3, -42, 31, -33, 124, 71, -31, 72, -64, -105, 86, -43, -77, 66, 80, 94, 40, 99, -51, -28, -70, 87, -27, -19, -8, -46, 28, 45, -99, 26, 67, -78, -44, 37, -81, -63, 10, -17, 3, 20, 126, 92, -76, 112, 47, 73, -124, 29, -123, -107, 43, -33, -21, -48, -88, 34, 58, -69, 52, 72, -28, -71, -2, 39, 89, -78, -75, -63, -85, 103, -37, -46, 26, 47, -23, -74, 27, -88, -26, -4, 25, -128, 41, -19, 79, 58, 75, 96, 33, -75, 77, 126, -68, -66, 95, 98, 48, 0, -44, -68, 3, -99, -31, 106, -70, -55, -88, -64, 11, -124, -70, -80, 25, 65, -7, -124, -77, 10, -36, -62, -62, -27, 90, 112, -67, -121, 50, -102, -103, 12, -71, -10, -30, -92, -12, 87, 57, 78, 85, 89, 0, -80, 41, 60, -43, 40, 80, 94, 21, -114, -21, -124, 59, 13, -111, -87, 4, 91, 57, -4, 14, -11, -116, -57, -16, 118, 15, 20, -72, -18, -47, -2, -44, -114, 97, -89, 11, -4, 1, -94, -55, 21, 6, 52, 78, -86, 4, -18, -105, -84, -28, -28, -76, -64, -60, 104, -28, -73, 109, -39, -117, -107, 56, 9, 98, 64, -54, 95, 123, 45, -40, -51, -31, 122, 35, 29, -81, -99, 122, -35, 31, -53, -36, 126, 29, 115, 121, 16, 124, 70, 10, -47, -98, -14, 102, 55, 126, 66, -74, 69, 30, 9, -74, 2, -125, -4, -33, -66, -114, -75, 67, 64, 10, -78, -5, 15, 37, -8, 120, 85, -99, -95, 116, -44, -126, 79, 14, 20, 81, -49, 57, 4, 1, 24, -119, -51, 93, -21, 107, 44, 90, 110, 97, 2, 80, 13, -71, 0, -34, -44, -107, 64, -44, 89, -8, 113, -55, 90, 72, 26, 52, 48, -7, 49, 84, -48, 122, -112, 90, -27, 113, -98, 126, 67, 57, 44, 73, 91, -105, 88, -38, -53, -104, 113, -83, -60, -12, 65, 31, -40, 121, -87, 112, 116, -81, -23, 77, -78, 48, -68, -76, 86, 56, 91, -74, -3, -5, 1, 83, 14, -54, -50, 83, 111, -45, 44, -106, 32, -123, 57, 37, -72, -98, 70, -36, 15, -36, 96, -121, -101, 10, 6, -119, -103, -57, -16, 68, 84, 77, 11, 28, -44, -50, 81, 74, 86, 127, 112, -34, -54, -89, -94, -116, 127, -88, 15, -123, -31, 103, -48, -111, 98, -14, -57, -36, 94, 23, 63, -16, -109, -63, 56, 113, -120, -21, 37, -90, 81, -113, -19, 92, 17, -27, -118, -52, -113, 101, -40, 101, 91, 65, -117, 125, -1, -99, -53, -114, 71, 27, -8, -103, 76, -89, -6, 12, 57, 8, -101, -108, 74, 80, -9, -81, -41, 91, 60, -113, -125, 32, 62, -68, -108, 57, 65, -101, 14, -4, -30, -108, 105, -109, 70, -13, 59, 53, 57, 19, -35, 17, -24, 113, -65, 111, 122, 91, -91, -86, 60, -122, -121, 76, 57, -41, -123, 41, -81, -122, -66, -67, 104, -127, -125, 33, 58, 87, -39, 122, -82, -68, 113, -59, -12, -120, -24, -126, 92, 66, -126, 32, -120, 41, 36, -32, -105, -78, 26, -114, 5, -10, 31, 22, -58, -94, 43, -27, 34, -38, -8, 67, 15, 109, 78, -14, -11, 81, -66, 24, 17, 32, -38, 45, 80, 32, 96, 33, 16, -106, -125, -36, -119, 30, 79, 113, -46, -80, 28, -109, 23, 13, -92, 109, 24, -6, -36, 112, 125, 39, -114, -24, 111, 50, 7, -75, 0, 20, -57, -53, 28, 87, -126, 60, -29, 23, 61, -26, -123, 42, 80, -33, 97, 48, 48, -35, -7, -10, -118, -122, 74, 80, 100, -107, -14, -8, 54, 45, 51, -72, -110, 64, 4, -128, 5, 43, 15, 85, 20, -27, 101, 55, -85, -25, -2, 63, -74, 92, 46, -95, -41, 94, 120, -111, -49, -47, -78, 24, 86, 126, -93, 90, 83, 64, -99, -124, -100, -51, 98, -83, -85, -44, 54, 112, -33, -5, -28, 30, -82, -33, 56, 3, -60, 48, -93, -20, 21, -39, 94, -67, -95, 1, 124, 101, 53, -122, -25, -26, -99, -112, -80, -26, -15, -111, -49, -58, -113, 93, 57, 45, -14, -44, -73, -10, -55, 3, -122, 53, -54, 119, -95, -79, 31, -79, -14, 54, -89, -20, 74, -62, -71, -105, 20, -47, 24, -34, 46, -120, -16, 111, -20, 99, 113, -61, -14, -109, 122, -65, 100, -24, 39, -34, 87, 64, 70, 8, -23, -103, -78, 2, 36, 2, 35, 98, -118, -35, -114, 26, 110, -48, -90, 41, 48, 126, -39, -13, 92, 92, 83, 10, -67, 99, -47, -8, 8, -70, -17, -101, -7, -116, -37, 4, 66, -35, 10, 109, -102, 49, 81, 110, 39, 0, 6, -30, -17, -121, -51, 48, 76, -90, -78, -9, -30, 15, -89, 45, -89, 124, -57, -27, 71, -60, 30, 110, -29, -6, -50, 14, -29, 117, 51, -4, -42, -115, -89, 45, 57, -84, -58, -72, 118, 8, 125, -52, -121, -23, -15, -33, -74, 86, -120, -77, -122, -107, -99, -49, -96, 68, 71, 65, -36, 85, 119, -63, -48, 105, 49, 21, -84, 22, -53, -28, 68, -107, -103, -12, 43, 51, 79, 55, 112, 8, 101, -2, -126, 57, 10, -4, 59, 126, -101, 17, -25, -65, -24, -118, -84, 58, 52, 127, 3, 89, 27, -86, -124, -18, -88, 93, -63, 67, -77, -28, 27, -102, 113, -115, 8, -36, -54, 109, 48, -31, -50, 28, -79, -36, -124, 41, 95, -70, -53, -120, -13, 37, -25, 0, -79, -119, -43, 82, -78, -11, -72, 20, -78, 103, 74, 70, 51, 90, -110, -88, 92, -119, -53, 88, -7, -80, -125, -71, 109, -38, 69, 77, -29, -110, 72, -26, 122, -82, 48, 37, -16, 46, 84, -17, 127, -68, 68, -40, 75, 61, -80, -84, -3, -25, -6, 53, 18, -101, 83, -48, 121, 76, 81, 6, 76, -106, 109, -84, -61, 54, -106, 28, 113, 11, 27, -47, 118, 62, 28, 99, -88, 3, 52, 45, -35, 60, 25, -104, -15, 116, 21, -91, -112, 78, -95, -46, 88, 61, -116, -39, -10, 103, 66, 4, 118, 81, -62, 51, -14, -29, 59, -122, 7, 44, -57, -91, -116, -108, -108, -123, -127, 101, 75, -10, 26, -56, -34, -18, -43, -42, -57, 74, -23, -63, -75, -80, -80, -32, -71, 13, -69, 104, 53, -68, -35, -118, 52, 96, -117, -128, 41, 65, -55, 90, -62, 80, -56, -1, 109, -36, -27, 95, 68, 85, -91, -45, -56, 77, -46, 32, -66, -113, 27, 23, -22, 49, -8, -9, -16, 9, 8, 112, 92, -53, 21, -102, 37, -41, 69, -19, 88, 106, 62, -122, 74, -14, 63, 100, 121, 105, -14, 9, -5, 64, 103, 99, 75, -21, 70, 53, 54, -86, -114, -94, 89, 72, 101, -66, 111, 86, 60, -126, 108, 23, 15, -54, -25, 36, -46, -57, 37, 25, -103, -125, 3, -40, 22, -43, -57, -44, -115, 55, 15, 68, -41, 91, -94, 123, -108, 59, 57, -75, -90, 10, 23, -69, -80, 38, 81, 58, 57, -78, -112, -48, 58, -122, -96, -9, 9, 54, -52, 116, 67, -113, -80, 34, 89, 99, 103, 115, -110, -96, -1, 96, -8, 60, 50, 79, -77, -28, 12, -101, -53, 117, 48, 108, 52, 113, -90, -100, -66, -48, 0, 85, 125, 5, -99, 17, 99, 84, -18, -66, -20, 99, 112, 44, -9, 25, -105, 5, -10, 98, 107, -92, 49, -27, -110, -93, -68, -117, -41, 114, -22, 101, 55, 61, -76, -5, -28, 8, -23, 57, -30, 62, 16, 78, 22, 12, 78, -47, -116, -81, 100, -75, -81, 74, -87, 98, 93, -119, 123, -86, -20, -17, -8, -9, -123, 12, -24, -33, -43, 79, 43, -86, -86, -10, 103, 2, 67, 75, 26, 17, 113, 23, -90, 55, 64, -120, 81, 75, 10, -126, -7, -83, 8, 105, -81, -104, -52, -119, -105, 86, 61, 74, -43, 15, -2, 24, 41, -64, -63, 7, 116, -36, -34, 118, -92, -57, 92, -91, -17, -20, 4, 73, -106, -38, 78, -39, 116, 19, 100, 38, -51, -70, -53, 61, -95, 92, 100, -32, 112, -97, 87, -7, 31, 46, 95, -27, 46, 12, -103, 92, -2, 19, 9, -100, 32, -120, -72, 15, -73, -71, 42, -88, -41, -126, -70, -64, 99, -123, 124, -19, -6, 62, 12, -120, -118, 110, -53, 118, 86, -69, -117, -73, -110, -44, 86, -118, -9, -76, -68, -95, 101, 108, 10, 53, -80, 91, 11, -99, 30, 97, 44, -73, -69, 108, -63, -110, -55, 102, -24, -99, -60, 103, -22, 108, 53, 79, -83, 77, -52, -124, -80, -4, -63, -83, -81, -49, -114, 104, -22, -21, 67, -127, -20, 57, 9, -97, 81, -68, -110, -79, -66, 106, 60, 117, 83, -70, 57, -7, 112, -26, -92, -3, 14, -35, 0, 88, -125, -79, 6, 47, 19, 51, -109, 91, -93, -122, 93, -77, 95, 87, 112, -52, -118, 76, 6, -36, 36, 31, 29, -20, 29, -127, -27, -1, 55, -93, -120, 24, 30, -112, 67, -106, 47, -71, 45, 72, -101, 15, -115, 45, 33, -5, -42, 66, -66, 94, 35, 93, -33, 30, 120, 27, -85, 26, 91, -94, 31, -116, 43, 8, 66, 55, 18, 73, -117, -41, -76, 19, 36, -23, -98, -11, 127, 83, -125, -80, 45, 27, -104, 47, 16, -99, -121, -97, -90, -31, 8, 54, -98, 12, 16, 46, 86, 101, -10, 53, -6, 15, -118, -118, -78, -100, 115, 95, -5, -64, 83, 0, 0, -6, 76, 71, -44, -120, -82, -29, 81, 2, -121, 104, 22, -29, 2, 104, 40, 19, -92, -121, -23, 68, 0, 0, 122, 60, 88, 51, 74, -84, -92, -11, -22, -55, -15, -4, 114, 14, -46, 44, 59, -41, -101, 19, -70, 30, 84, -73, -68, 27, -26, -84, -122, 123, 63, 63, -86, -13, 76, 59, -103, -58, -121, -100, -100, 114, 74, 125, -13, -79, 112, 78, 44, 113, 9, 113, 90, 26, 72, -124, 88, -43, -122, 73, 88, 27, 37, 60, -114, 50, -115, 103, -106, 57, -41, 93, 25, 74, -123, -4, 32, -3, -53, -68, 108, 4, 106, 61, 123, -4, -117, 127, -53, 64, -14, 113, -48, 103, -24, -73, 95, 27, 16, -110, -11, 12, 60, 7, -38, -108, 111, 48, 94, -25, 21, 106, -43, 44, 5, 36, 4, 31, 63, 15, 125, -15, -27, 64, -106, 121, 63, 65, 15, 79, -103, -120, 96, -41, 30, -92, 46, 11, 118, 26, 110, -118, 86, -50, 47, 113, 64, 102, 73, 49, 118, -115, 17, -4, 51, -63, 98, -84, 30, 30, -73, 63, -108, 51, 17, -116, -123, 36, -23, 37, -59, -126, -41, 20, 63, -12, -113, -17, 65, -66, -53, 47, 106, -81, 30, 43, -97, 33, 36, -17, 53, 32, -96, 59, -128, 36, -62, 27, 115, -21, -70, -5, -85, -79, -49, -77, -67, -31, 16, -52, -34, -113, 8, -114, -3, -74, -69, 122, 116, -111, -89, 89, -89, 123, 76, -127, -19, -97, 71, 60, -119, 87, -83, 70, 125, -75, -46, -75, 89, -29, 48, -119, -80, -69, 127, 27, -12, -46, -77, -25, 123, -21, 21, -64, -85, -6, -23, -87, 50, 7, 116, -111, -41, -76, 57, 69, 102, -24, -46, 70, -50, 121, 43, -118, -34, -115, 126, 26, -78, 82, -3, -104, 93, 68, 127, 98, -19, 35, 69, -76, -14, -17, -26, -67, -66, 47, 105, -127, 102, 49, 85, -17, 52, -124, -109, -73, -125, 57, -3, 68, -16, -64, -71, 123, 105, -78, -8, 25, -86, 29, 22, 92, 41, -63, 23, 104, 10, 32, 24, -76, 33, 106, -50, -43, 83, 99, 57, -109, 65, -70, 119, 30, 17, 86, 5, 13, -22, 104, -34, -23, 63, 27, 116, -3, 104, 41, 39, -45, -87, -37, -108, 1, -21, -15, 94, -94, -58, -72, 44, -108, -70, -74, 45, -31, -52, 77, 0, -45, -9, 52, -124, -103, 31, 120, 96, 6, -4, 106, 43, -128, -99, 67, 24, 43, -6, -98, 36, 37, 57, -99, -65, 10, 51, -104, 86, 115, 19, -101, -10, 73, 58, -15, 15, 102, -77, -105, 120, -29, -93, -119, 93, 58, 24, -43, 66, -11, -91, -100, 62, 82, -109, -20, -71, -26, -60, 30, 5, 9, -75, -32, 86, 45, 28, 44, -21, 51, 3, -35, -11, 102, 90, -36, -38, -22, -102, 24, 29, 33, 73, 61, 112, -102, 104, -7, -63, -65, 3, -9, -48, 117, 55, -50, 84, -92, 32, -127, -66, 68, -44, 127, -38, 33, 2, -67, -43, -93, -21, 33, -111, -46, 46, -58, 109, -11, 96, -22, -10, -65, -44, 2, 93, 68, -13, 10, -104, -69, 63, 29, 69, 24, 21, -70, 7, 36, -45, -100, 112, -73, -115, -76, 32, 13, -124, -5, -110, -37, -121, -29, -35, -17, -52, -102, 103, -63, -76, -33, 124, 95, 16, -42, -65, -124, 29, 104, -75, -84, -44, -44, -14, 33, -45, 107, -41, -59, 57, 77, -86, 2, 64, -106, -17, -39, -44, -54, -16, -119, -108, 76, 113, -122, 73, -62, -99, -33, -54, -102, -32, -48, -126, 9, -122, -30, -62, 56, 34, -59, -110, -47, -62, 28, 83, 4, 72, 57, 89, -94, 24, 100, -38, 22, -28, -22, 17, 65, -68, -11, 57, -73, -10, -112, 105, -34, 30, 59, -32, -45, -90, 52, -60, 19, 9, -31, -80, 55, 94, -1, 85, 127, -105, -35, 107, 78, -81, 114, 118, -127, 36, -64, 64, 114, -117, 6, 36, -67, 4, 79, -13, 115, 43, -95, 4, -1, 12, 9, 87, 69, 98, -11, 92, 83, 4, -6, -37, 10, -19, 60, -114, 92, -88, 108, 125, -14, -46, 95, -29, -43, -103, -35, 107, 126, 63, 4, 117, 16, 71, -43, -60, -60, 22, -12, 2, 45, -91, 113, -68, 119, -17, 114, 60, 7, 77, -24, -92, -28, -108, 78, -21, -45, -41, -7, -91, 81, -46, -1, -126, -66, 97, 93, 40, -85, -26, 123, -103, 97, -35, 70, 25, 42, 91, 36, -57, -9, -114, -124, 51, -106, 54, -3, -45, -43, 46, 30, -26, 78, -92, -58, 43, -102, 93, -87, 110, 122, -34, 12, 104, -121, -85, -44, 75, 76, 9, -74, -128, 54, -34, -70, 76, -14, 85, -1, 11, 127, -29, -13, 36, -28, -44, 16, -29, 66, 89, -56, -125, -20, -24, -16, -54, -61, 99, -99, -64, -12, -57, -26, 69, -124, 108, -51, -127, -11, 93, 36, -123, -20, -33, -55, 118, 3, -72, 10, 43, -93, -110, -72, -47, 21, -79, -28, 86, 89, 75, 15, -73, 52, -31, -29, 75, -89, 65, -76, -29, 39, 44, 20, -110, -36, 98, -64, -4, 21, 117, 13, -21, -19, 120, 52, -5, 43, 45, -2, 100, -121, 66, 80, 29, 103, -42, 105, -107, -55, -125, 72, 12, -125, 59, 6, -14, 1, -128, -51, -113, 112, 125, -106, -96, -39, -47, -102, -121, 103, -5, 23, 103, 18, -13, -127, -121, -79, 82, 20, -16, -8, 52, -38, -19, 39, 58, -11, -27, 123, -20, 26, -125, -62, 28, -112, -19, -39, 91, -49, 50, 60, -62, -118, 96, -101, -55, 14, -59, 60, -40, -73, -52, 60, 31, -41, 45, 16, 113, 74, -84, 111, 106, 112, -65, -91, -76, 100, -8, 69, -67, 19, -1, -40, -55, -42, 83, 120, -27, 89, 17, -55, -5, 40, -43, 34, 2, -37, 16, 17, -76, -8, 119, 68, -14, -26, 114, -21, 42, -66, -42, 39, -100, 88, -105, -102, -70, 122, 55, -75, 95, -84, 55, -18, 76, 100, 85, 25, 111, -33, 57, 61, -44, 53, -51, -113, -49, 75, 57, -13, 55, 3, -42, -22, -15, 81, 104, 27, 64, 27, -119, -41, 33, 67, -61, -74, -81, 56, 6, 85, -74, -118, -50, 88, 94, -126, 14, -34, -66, -69, 27, -19, -23, 34, -90, 112, 123, 19, 81, -113, 116, 83, 106, -30, -83, 63, -107, -34, 72, -32, 125, -52, -22, -110, -77, -76, -82, -122, -116, -72, -106, -65, 121, 117, -80, -106, 45, 70, 44, -6, -90, -22, 78, 38, -70, -115, 100, -48, -64, 58, 46, -75, 42, -18, -109, -124, 4, -123, -54, 52, -74, 74, -80, -60, -82, -25, -66, -94, -78, 3, 66, 54, -24, 59, 59, 7, -34, 122, -93, -77, -109, -82, -51, 123, 20, -128, 62, 47, 9, 73, 52, -92, 12, 80, -80, 73, 49, 79, -94, -101, -8, 77, -104, -66, 20, -68, -24, -60, 57, -101, -24, 62, -11, 66, -115, 127, 87, 29, -53, -24, -42, -116, -119, -116, 83, -40, 10, 40, -77, 31, -87, -46, 65, 11, 71, 82, -38, -58, -56, -75, 6, -79, 103, 123, -101, -14, 50, -15, 47, 98, -27, -87, -76, -2, -4, 31, -99, -28, -28, -82, -10, -15, 42, -122, 104, 126, -119, -124, 119, -85, 73, -98, 14, -85, -36, -64, -110, 40, 70, 53, 108, 91, -20, 79, -59, -12, 40, -5, -90, -46, 2, 36, 39, -48, 116, -55, -28, 55, -98, 12, -9, -117, 114, -25, 109, -64, -99, -12, 11, 117, -113, 46, 38, -109, 94, -36, 12, 106, 105, -71, -74, 69, 87, -55, 83, 0, -72, -88, -45, 113, 7, 14, -106, -12, 55, -13, 48, 103, -44, 43, 109, 38, -120, -115, -102, -37, 73, 28, 54, 73, 48, 49, -118, -95, -3, 13, -20, 0, 97, -83, -20, 90, -71, 62, 18, 34, 9, 85, -43, -58, 107, -115, -68, -10, -52, -52, 100, -5, 20, -73, -85, -18, 110, -113, 85, -96, 47, -114, 56, -90, -71, 78, -4, 9, -101, -75, -128, 116, 62, -116, 42, -127, -82, 95, -20, 99, 2, -29, 110, 3, 17, -97, -93, 48, -74, 14, -59, 20, 59, 127, -124, 55, 64, 93, 78, -12, 64, 89, 36, 40, 109, -52, 86, -22, 41, 44, -112, -53, -3, -57, -35, 87, -62, 10, -97, 112, 40, -12, -20, 63, 95, 26, 96, 20, -7, 41, 60, -52, -121, 9, 28, -3, 113, 102, -8, 102, 114, -115, 83, 109, 89, -78, 104, 71, -8, 107, 52, -34, -64, 79, 107, 46, -89, 4, 77, 67, 103, 121, 54, 67, -67, -58, 1, -37, 8, 52, -77, 10, -80, -117, 32, 41, -44, 31, 68, 32, -15, 23, 44, 20, -16, 90, -45, 54, 121, 11, 98, -83, -24, -6, -28, -125, 121, -105, -57, 102, -89, 30, -58, -98, -85, 95, 29, 22, -117, 14, -61, -9, 46, -79, -88, -88, -95, 72, -80, 58, -121, 127, -40, -66, 59, -49, -69, 56, -100, 79, 58, 89, -61, -92, -68, -66, -31, 89, 105, 21, -95, -95, 105, -84, -99, 74, -85, 5, -22, 117, 9, 1, 73, -91, 111, 119, 10, 14, -99, 81, 4, 86, -44, -16, 67, 109, -94, -94, -94, 52, 40, 105, -40, 126, 90, -7, 73, 6, -102, -117, 17, 108, 91, 81, 32, 82, 15, 125, 17, -6, 126, 35, 59, -35, 19, 19, 5, 64, -26, 0, 3, -107, -124, -81, 19, 60, 35, -86, -76, -103, 121, 7, -64, -8, -7, -60, -38, 3, -29, 18, 63, 99, 67, -66, 111, -64, -23, -77, 14, -43, -80, -52, 36, 73, 88, 10, 36, 96, -60, -80, -88, 90, -69, -76, 37, 8, 40, 121, -68, 46, 38, -114, -10, -92, 120, -6, -25, 13, 10, 31, -23, 45, 79, 52, 42, -71, 12, -125, -55, 126, -15, 125, -2, -94, 76, 54, -124, 7, 63, 59, -114, -29, -66, 69, 96, -118, 106, -102, -29, -6, 27, -92, 42, -67, -109, -127, 24, -114, -48, 79, 20, -95, -34, -126, -82, 45, -89, 95, -28, 84, 43, 97, -71, 6, -14, -101, -63, 30, 45, -102, -87, 114, -117, -119, -67, -27, -112, -11, 22, -98, 4, -109, 96, -112, -55, -64, -23, 33, -128, -19, -77, 0, 65, 6, -51, 37, 18, -52, -110, 100, 122, -125, -87, 73, -124, 78, 74, 97, -101, 112, -76, -63, 85, 111, -120, 63, -74, 33, -122, -109, 45, 56, -117, -11, -100, -42, -19, 39, 117, -42, 62, 51, -93, 74, 8, -28, -86, 43, 55, 51, -68, 63, 36, 45, 59, -113, 106, 73, -68, -61, 61, -121, -5, -2, 48, -112, 70, -23, -37, -25, -109, 26, -30, -120, 70, 120, 82, -31, -118, 115, 40, 77, 123, -97, -78, -115, 117, 0, 81, -97, -65, 94, -56, 95, 77, 18, -34, 21, -120, -5, -52, 80, 32, 110, 50, -50, -35, -39, 41, 115, -65, 13, 69, 32, -22, -104, 96, 51, -64, 4, -73, 91, -32, -76, -116, -66, -107, -84, 82, -8, -42, 42, 119, -125, 108, 126, 117, -116, 102, -128, -77, -1, 53, -32, 6, 1, 25, -48, -5, 25, -12, -31, 80, -49, -29, -56, 123, 111, 6, 106, -60, -128, -112, -4, -18, -10, 10, -115, -58, -14, -97, -59, 4, 4, -115, -2, 77, 86, 67, 88, -1, 97, -24, -14, 10, -5, -25, 120, 118, -96, 56, 75, 29, 117, -116, 116, 17, -116, -110, 73, 114, 2, 60, 21, 57, -48, 59, 26, -1, -90, -97, -93, -87, -117, 77, -5, -115, 71, 125, -10, 59, -120, 85, -60, -91, 0, 124, -10, -46, -89, -104, -17, 14, -99, -128, -87, -68, -91, -37, 70, 42, 61, -72, -25, -58, -83, 105, 55, 10, -113, -7, 60, -83, -20, 125, -120, -102, 97, -7, 65, 72, -106, -87, 102, 114, -49, 11, 17, 50, 32, 15, -1, -110, -82, 124, -46, 104, 49, 61, 72, 19, 86, 24, -93, -21, -96, -54, 107, 87, 61, 85, 116, 9, 59, -68, -79, -99, 101, -95, 100, -17, -13, -55, 63, 113, 66, -38, -109, -125, -72, 42, -5, 33, 36, 82, 31, -51, -12, -118, 113, 76, -122, -17, -71, 37, -25, -61, 13, -70, 82, 89, -73, 72, -112, -58, -111, 120, -17, -58, -104, 124, 121, 110, 23, -106, -57, -17, 83, -13, 10, -53, -128, -3, 76, 83, -92, 87, 30, -39, -57, 45, 93, -81, -34, 47, 121, -86, 1, -6, 47, -2, 5, -60, -101, 28, 114, -3, 92, -103, 5, 63, -101, 69, -45, 52, -86, 113, 20, -14, -29, 97, -61, -103, -30, -82, 38, 103, 61, -28, -76, -14, 73, -127, -22, -24, -55, -77, 28, 69, 31, 13, -4, 52, -34, -27, 8, 102, -31, 38, 69, -62, 17, -7, -86, -10, 70, -96, -80, 105, 40, -25, 105, 114, 119, -10, 69, -101, -16, 2, -49, 92, 121, 70, -24, -73, -46, -37, -13, 127, -39, -25, 117, 5, -23, 109, 105, 96, -110, 105, -49, -53, 44, 115, -32, -57, -49, 120, 71, 57, 87, -67, -41, 103, -20, 17, 123, 107, 95, -108, -103, -4, -124, -127, 15, 50, -23, -32, 61, -126, -42, 31, 77, -67, 78, 19, 58, 109, -123, 85, 10, -120, -83, -17, -63, 11, -46, 117, -40, 44, 68, 70, -58, -102, 61, -24, 55, -58, 86, -14, 105, -29, -109, 37, -16, -120, -105, -59, -102, -123, 92, 127, -103, -90, -128, -28, 10, -102, -67, 113, 20, -19, -121, 1, -68, 91, 88, 100, -114, 73, 82, 104, -114, 8, 98, 79, -96, -99, -85, 55, -40, -73, 23, 107, 28, -123, 67, 112, -57, 108, -6, -32, 8, -45, 111, 79, 28, -26, -85, -20, -79, 102, -36, 126, 47, 97, -41, 69, -31, 51, -76, -77, -70, 85, -115, 11, 73, 92, 65, 95, -118, -62, -2, -20, -15, 97, 19, -71, 29, 8, -122, -12, 117, -27, 3, -114, 86, 87, -89, -84, -6, 27, 60, 73, -63, -62, -125, -16, 22, -124, -2, -88, 13, -128, 88, -79, 82, 45, 109, -63, -24, -76, 120, -110, -25, 15, -20, -46, 64, 90, -12, 78, -103, -98, -78, 76, 127, -23, -1, 71, -77, 111, -93, -41, -61, -37, -88, -114, 115, 70, -36, -91, -125, 26, -108, -60, -116, -34, 74, 115, -126, -105, 15, -66, -111, 42, -65, 124, -51, -107, -86, -60, 23, -24, 40, -42, 47, 110, 27, -71, -51, -88, 110, 121, 57, 98, -107, 89, -44, -11, -68, 17, -12, -72, 79, -44, 14, -44, 7, -93, -54, -29, 62, 38, 93, -59, -91, 106, -10, -125, 3, -44, -85, 121, 126, -97, -6, 5, -97, 127, 63, 36, 1, -75, 47, -27, 97, -90, -80, -115, -69, 50, -77, -91, 36, 58, 112, 85, 31, -45, 41, 104, 86, 13, 33, 58, 1, 122, -86, -40, 76, -26, 41, 69, -12, -92, 70, 86, 11, -93, -122, -86, 51, 22, 125, 37, 85, -92, 21, 19, -116, -92, 68, 99, -97, 28, -17, -110, 21, 72, 114, -34, -80, 106, -73, 78, -17, 10, 0, -90, 116, -114, 89, -100, -21, -1, -24, -46, 109, -84, -59, -74, -80, 29, 74, 4, -73, -26, 83, 58, -51, -117, -38, 59, -75, -68, -22, -3, 99, 59, -104, 10, 69, 105, -124, 101, 62, -75, 54, -53, 122, -120, -50, -94, 115, 30, 25, -58, -18, -69, -74, -1, -117, -106, 97, -16, -24, 25, -103, -67, 103, 103, 97, -72, 33, 108, -43, 30, -86, 50, -83, 13, -82, 26, 19, 90, 32, -53, -59, -99, 53, 71, 13, 43, 117, -45, 1, 58, -73, 71, -49, 15, -97, 127, 16, -69, -44, 63, 47, -110, -44, -1, -107, 118, 99, 62, -122, 93, -18, 90, -65, 43, -86, 89, 34, 54, -127, -81, 119, 100, 77, 123, -5, -65, -82, -36, 47, 103, -123, 92, 98, -38, -64, 0, 41, -44, 11, 102, -108, 60, -56, 64, 51, 39, 85, 0, -20, -95, 7, -5, -92, 29, -109, 90, -10, 106, 8, -34, 19, 18, 75, -65, -14, 119, -126, -95, -40, -2, 106, 20, 87, 72, -65, 8, 65, -79, -94, -51, -84, -75, 43, 10, 109, -102, -110, -96, 109, 23, -77, 91, -53, -60, -64, 59, 79, -9, 124, 42, 109, -73, -111, 68, -119, -10, -43, 109, 21, 117, 109, -26, 36, -17, 35, 53, -23, -11, -29, 20, 87, -86, -112, 78, -96, 12, -7, 23, 4, -67, 95, -76, 12, -100, -3, 110, -22, 85, 23, -115, -45, -21, 102, 3, 43, -51, 76, 123, 117, 10, 37, 67, 33, 57, -29, 30, -46, -51, -111, -105, -115, 4, 45, -55, -54, 90, 114, -87, 85, -10, 114, -75, -27, 19, -32, -27, -97, 28, -58, -39, -103, 15, 31, -16, -99, -5, -105, -28, 92, 109, 67, -109, -6, -4, -81, 112, -18, 72, -123, 116, 124, -22, 86, -19, -22, -88, 54, 89, 58, -5, -74, -13, -14, 108, -101, 97, -44, 66, -85, 122, 46, 39, -17, 113, -44, -2, -73, 19, 54, 9, 80, 13, 116, 34, 78, 44, -99, 29, 127, 101, 89, 52, -88, 1, 23, -40, 13, 43, -94, -114, 63, -106, 30, 35, -98, -28, -86, 57, -22, 64, -123, -101, -20, 30, 80, -80, 81, -69, 85, 110, -91, 60, -127, -119, 32, -42, -97, -109, 95, -54, -8, -18, 7, -40, -100, 65, 108, 76, -99, 89, 35, -114, 43, 72, 12, 5, 62, 107, 19, 3, 10, -99, -35, -113, -51, 81, -19, 108, 27, -62, 26, 17, 64, -61, 19, -99, -72, 3, 50, -8, -37, 104, -103, 100, 13, 36, -74, 41, 16, 109, -48, 44, -11, 85, -80, -27, -51, 82, 12, -45, -92, 61, -24, -72, -10, 76, -36, -80, 49, 91, -82, 104, 74, 16, 104, -47, 17, 77, -29, -32, 19, -55, 120, 119, -81, 115, -78, -84, -39, 21, 110, -101, 90, -79, 21, 68, -14, -42, -59, -122, 106, 53, 59, -87, -29, 67, 48, -32, 105, 111, 14, 62, -12, -124, 91, 55, 83, 42, -41, -20, 55, 125, 66, -63, -118, 7, -110, -39, -53, 12, 126, -111, 5, 76, -116, 116, 5, -60, -96, -13, -58, 84, 63, 20, 38, -79, 54, 42, -16, -69, 27, -78, -104, -24, -36, -110, 3, -108, -97, -78, -36, -75, -94, 44, -101, 110, 90, 115, 99, 43, 15, 46, 79, -12, 86, -105, -17, 78, 55, -115, 68, -78, -81, 89, -14, 110, -118, -47, -12, 30, 20, -45, 54, 37, -50, -20, 39, -67, 68, -13, -21, -41, -48, -106, 98, 78, -104, 49, -69, 14, -68, 123, 75, 60, 112, 101, 27, -35, -54, -98, 124, 21, -58, -85, 12, -83, 28, -77, 28, -117, -122, -93, -88, 109, 39, 48, 23, 74, -46, 43, -98, -53, 88, -102, -61, 29, 25, 94, -15, -85, -82, -71, 21, 66, 37, -66, -53, 51, -121, -76, -47, -1, -83, 23, -6, -46, -1, 96, 12, -50, -48, 119, -74, -78, 68, -77, -110, 86, -96, -58, 1, -82, -57, -5, 69, 107, 104, 41, 43, -80, -28, 17, -26, -86, -119, 112, -72, -56, 68, 71, 14, 4, 80, -42, 108, -119, -92, 84, -63, -25, 87, 109, 99, 53, 120, -37, -71, -35, -24, 62, 19, 1, -79, 118, 54, 1, 1, -114, 19, -35, 24, 65, -71, -5, 6, 107, -67, 8, 9, 122, 11, -74, -26, -84, -75, 23, -50, -1, 51, -99, -67, 41, -100, -74, -59, 89, -16, -10, 48, 17, 62, -14, -126, -14, 30, -54, 62, -32, -102, -103, -69, 110, -5, -41, 75, -49, 53, -1, 89, -52, 62, -22, -60, -13, -8, -127, 16, -88, 15, -107, -25, -68, -70, 75, 16, 87, 60, 99, 40, 111, 0, -84, -101, 121, 3, 59, 74, 10, 45, 107, -93, 15, 81, 70, 23, -56, 65, 109, 123, 115, 120, -96, -88, 68, -49, 64, 36, -28, -23, -34, -50, -75, -50, -95, 121, 100, -54, 90, 23, 98, 120, 31, -42, -43, 109, -88, 24, -42, -66, 22, -95, -118, 56, 30, 91, 47, -44, 106, 77, -75, -24, -85, 19, -22, -61, 49, -104, 19, -99, -76, 8, -83, -76, 11, 18, 98, 100, 65, -25, 75, 103, -36, -87, 86, 105, -92, 87, -9, -29, 93, 16, 15, -60, 104, -119, 2, -40, -9, -110, 118, -61, -26, -79, -37, -2, -120, -55, 0, 120, -88, -67, 103, -18, -124, 69, -105, -112, 3, 79, 102, -58, -83, 0, -44, -80, 89, 36, 93, 85, -54, -56, -46, -33, -25, 66, -97, -110, -18, 94, 13, 38, -24, 12, 33, -122, -50, 4, -104, 15, -12, 77, 15, -53, -28, -46, -111, 18, 67, 116, -116, -40, -84, -106, 112, -73, -124, 118, 90, 82, -107, -38, 72, -85, 101, -34, 57, 33, 97, -127, -90, -48, 83, 13, 82, 58, -59, -99, -64, 29, 68, -65, 21, 106, 5, 2, -97, -125, -72, 27, -126, -8, 77, -38, 15, 96, 39, 95, -100, 38, 96, 9, -23, -34, 43, 22, -15, 34, 79, -34, 32, 69, -114, 45, -62, 99, 115, 10, -7, -73, 123, 29, -86, 97, 83, -91, 106, -54, 37, 14, 1, 39, 35, -51, -27, 19, 115, -11, -50, 115, -41, 78, 94, 15, -80, 105, 58, 114, 43, 92, -42, -66, 72, -74, -59, 125, 6, 72, -115, 23, 97, 65, 122, -26, -60, 121, -68, 20, -115, 71, 112, -114, -36, -78, 27, -74, 93, 0, 80, -36, 19, -20, 111, -66, -109, 61, -94, -90, -25, -124, 116, -14, -17, -19, -27, 67, -70, 14, -7, -85, 64, -23, -62, 107, 101, 95, 31, 4, -3, 37, 76, -19, 123, -44, 74, -105, 80, 14, 54, -50, -1, -37, -88, -21, 79, -120, 115, -46, -110, -54, 94, -13, -62, 101, -2, 32, -86, 3, -108, 34, -13, -127, -84, 112, 116, 55, -53, 50, -5, -81, -3, -102, -50, -48, 126, 113, -118, -95, 23, 19, -43, -45, -28, 95, -20, 70, 75, -112, -40, -22, 37, -68, -36, -47, 118, 51, -16, 30, -42, -3, 74, 28, -95, 2, -127, -43, 106, -27, -95, 127, -104, -25, 87, -32, -7, 87, 84, -89, -28, -114, 79, 43, 94, -3, -106, -90, -28, -41, 83, -107, -8, 23, -16, 64, 93, 41, -116, -23, 77, 16, -6, -25, 119, 16, -2, -53, -34, -29, 27, 66, -37, 4, -24, 109, 61, 57, -102, -126, 60, 86, 28, -119, -39, 19, -32, 21, -22, -120, -48, 126, 1, 105, 4, 61, -7, -88, -17, 69, 93, 79, -24, -93, -92, 91, 24, 111, -112, 2, 60, 89, -44, 74, 21, -121, 3, -42, 28, 31, 16, -56, -29, 65, 5, -43, 75, 84, -59, -8, -100, 44, -58, -19, 35, 36, -16, 125, -66, -23, 97, -15, -83, 119, -59, -116, 25, -6, 124, -20, -78, -74, 68, 87, -124, -92, 37, 119, 19, 114, -120, 87, 61, -14, -46, -10, 95, -47, -61, 58, 27, 96, 6, 77, -78, -81, 11, -121, 44, 42, -27, -75, -54, 33, -59, 43, 103, 25, 114, 32, -89, 48, -9, 27, 90, -82, -46, -106, -29, 12, 21, -79, -117, -37, -41, 43, -63, 36, 20, 35, -37, 42, -24, 28, 69, -77, -42, -119, 67, 9, -62, -114, -46, 93, -85, -28, 72, -124, -36, 88, 73, 53, -48, 115, -22, 68, 78, 117, 43, -62, -32, 40, -98, -15, 42, -53, 73, 77, 34, 33, -35, -72, 14, -120, -56, 53, -78, -98, -12, -30, 60, -30, 96, -124, -70, 120, 13, -105, -127, 32, -107, -32, -82, -64, 115, -103, -122, -76, -96, -7, 6, 59, -20, -111, 58, -85, 64, 115, -67, -113, 8, 90, 39, -109, -103, 103, -26, 69, -110, 17, 95, -108, -93, 49, 40, -71, -35, -87, -27, 5, 112, 120, -78, 95, -7, 13, 94, -14, 66, 33, -69, 6, -34, -76, 73, -11, 114, 7, -77, -114, -24, -8, 87, 19, -35, 97, 117, 20, -87, 35, 28, -112, 118, 72, -98, 66, -120, -84, 41, -38, -101, 111, 58, 92, -47, -118, 30, -75, -5, -69, -115, -9, -67, -70, -80, 112, 48, 2, -20, -102, -29, -113, 23, 16, -30, 90, -111, 1, 105, 72, -95, -77, 2, -56, -118, -123, 49, 106, -77, -51, 94, -108, -117, 30, 75, -26, -13, 5, -47, -83, -39, 46, 114, -17, 57, -25, 68, 36, 11, -99, -70, 80, -72, -107, 65, -89, 59, -49, 92, 46, 119, 87, 16, 123, -30, 73, 47, 74, 112, -113, -66, 13, 100, -119, -124, 85, -59, -116, -44, -44, 106, -38, 41, 54, 46, 14, -37, -17, 108, -55, 1, 88, 126, -66, 96, 125, -82, -48, -58, -73, -62, -78, -108, 84, 1, 7, 93, -83, -15, -117, 28, 30, -52, -43, -36, -7, 61, -30, -12, 79, 27, -98, -115, 23, -25, -13, -27, -34, -24, -23, -23, 66, -6, -1, -30, -53, 46, -91, 121, -97, -66, 25, -91, -49, -1, 86, -71, 23, 11, -43, -84, -125, 12, -121, 69, -26, 71, -34, 16, -48, -75, -3, 6, -69, -60, 121, -63, -110, 99, 15, 118, -123, 34, -94, 42, -30, -46, -85, 52, -62, 83, -14, 8, -8, 97, -40, -75, 0, -118, 10, 98, 106, 78, 21, 88, 45, 13, 19, -77, -95, 72, 79, 3, 107, -29, -83, -102, -55, -128, 115, -75, 111, 125, -42, -89, -7, 123, 124, -115, -12, -97, 63, -79, -53, 57, 111, 30, -125, -85, -16, 11, -125, 127, 12, -126, -108, -35, 93, 30, 13, -98, 1, 57, -106, -31, 82, -15, 81, -125, -73, -55, 25, 31, 32, 75, 78, 117, -39, -79, -86, -124, -7, -36, -111, -52, -126, 112, 23, -16, -63, 115, -5, -54, 38, -68, 104, -113, 102, -65, -105, 102, -52, 116, 104, -15, 1, 11, -84, -37, -24, 103, 124, 21, -41, 73, 79, -122, 85, -114, -23, -92, -84, -69, -33, 11, -104, 82, 92, -1, -28, 7, -102, -113, -31, -6, 61, 37, -14, 27, -76, -119, 22, 35, -19, 5, -12, 87, 101, 51, 92, -48, -26, -94, 46, -87, 103, 64, -9, 107, 35, 31, -50, 57, 58, -128, -8, 19, 90, -1, -49, 90, 113, -4, 44, 46, 23, 112, 94, 7, -54, 46, 64, 4, 101, 96, 17, 41, 67, -45, -128, -85, 96, 84, -32, -6, -119, -48, -71, -11, 19, 87, 73, 44, 14, -29, 19, 79, -115, 76, 43, 121, 24, 125, -46, -80, -109, 32, 107, -78, 6, -61, 80, -44, 0, -29, 83, -28, -87, -91, -20, 71, 15, 56, -17, -114, -46, 10, -61, -71, -61, -111, -99, -91, 4, 66, 127, 47, -96, 39, 58, -64, -127, 20, 56, 127, 77, 78, 97, -69, -115, -72, 51, -82, 83, -71, -94, 73, 65, -45, 7, 50, 116, -39, -51, -65, -18, -48, -59, -69, -88, 90, -14, -111, 24, -43, 74, 76, -7, 60, 87, -33, -89, -121, -60, 15, 60, 102, -99, -28, 100, 6, 53, 117, -107, 92, 96, -62, 60, -125, 86, -90, 117, -97, 88, -14, 46, 83, -112, -112, 13, 122, -58, 96, 78, -38, -40, -77, 119, 24, 78, 43, 40, 7, 41, 49, 62, -127, 59, -73, -60, -28, 110, -119, 33, 101, 57, -47, 32, -71, -54, -65, -93, 110, 50, -29, 20, 16, 16, 56, 86, -123, -106, 17, 61, -42, -67, -23, -122, -35, 0, -81, -27, 64, 30, 97, -3, -62, 118, 127, -37, 111, -124, -84, 81, 21, 95, 43, -18, 23, 14, -120, 108, -125, 125, -115, -56, -117, 98, 84, -2, 22, -84, -1, 24, 19, -7, 116, 20, 96, -84, 108, -55, -34, 73, 34, -104, -43, 2, 7, 25, -23, -101, 97, 4, -26, -8, -127, -74, 81, 35, 53, 66, -67, 70, -54, -16, 37, 67, -45, 7, -49, 116, -45, 48, -83, 18, -14, 109, 89, -64, 62, 63, -39, -114, 105, -126, 67, -73, -18, 54, -108, 94, 66, -121, -92, 37, -5, 57, 59, -4, -58, -34, -28, -47, -86, 75, 5, -32, 104, 21, -121, -124, 113, -110, 67, 121, 18, -78, -27, 89, 60, 99, -4, 12, -87, 67, 68, 23, 105, -34, 124, 68, 126, 11, 89, -64, 115, -118, 83, -113, 39, -21, -77, -37, 73, -58, 85, -56, -17, -48, 8, 13, -109, 109, 114, -10, 89, 21, -44, 30, 113, -101, 72, -100, -65, -83, 47, 42, -26, 20, 37, 119, -107, -95, 41, -5, 37, -120, -95, -110, 126, -103, 119, -57, -90, -5, -44, 123, 110, -44, -41, -15, -42, -118, 60, 71, -8, -65, 22, -10, 57, 6, 71, 41, -83, -24, 54, -79, -60, 45, -83, 77, 33, 31, -109, -92, 10, -27, 95, 55, -103, -75, -111, 27, 31, 83, 51, 48, -23, -43, 69, 41, 116, -95, 15, 6, -22, -111, 39, 76, -125, -93, 50, -105, 14, -101, 108, -112, 8, 38, 106, 2, -90, -99, 78, -70, 39, 104, 7, 35, -107, -50, 37, -53, -41, 51, -18, 101, -115, -87, -5, -45, 4, 59, -96, -14, -126, -109, -49, -119, 28, 103, -17, 120, 25, 4, 52, 17, -85, -48, 99, 86, 60, -42, -63, -118, -76, 72, 96, 36, -95, 94, -13, -57, 47, 109, 37, 86, -40, -91, -101, -23, -2, 42, 30, 84, -74, -78, 91, 43, -85, 64, -77, -31, -91, 88, -29, -104, -23, -14, 113, 125, -88, 107, -62, -119, 26, 106, -63, -93, -18, -6, -62, -54, -82, -21, -51, 19, 21, 90, 95, 54, 12, -112, -25, 65, -37, -13, 62, -88, 15, 82, 8, 124, -40, 75, -124, 76, -41, 31, -49, 15, 44, 48, 37, -113, 100, -117, -25, 15, 72, -25, -39, -47, 15, -21, -118, -67, 41, 93, -16, 29, 69, -26, 87, -18, -47, 11, 117, -95, -69, -41, 67, 79, 34, 6, 102, 12, 36, -62, -23, 95, -41, -57, -74, 70, -30, -65, 78, -13, 37, -117, -112, 11, 75, -77, -15, -65, -75, -17, -19, -126, 29, -83, -40, -90, 55, -13, -90, -28, 11, 92, 115, -95, 81, -100, -41, 80, -110, 119, 98, 25, 78, -18, 46, 30, 12, -9, 109, 43, 93, 120, -45, 58, -115, 82, -15, 61, -106, 43, 127, -92, 111, -128, 120, 12, 68, -112, -8, 74, 102, -96, -98, 21, 125, 126, 114, 8, 83, 3, -5, -20, -4, -53, -73, -79, -101, 30, -125, -57, -91, 94, 94, 33, -72, 97, -117, 28, 24, 21, 20, -65, -19, -95, 62, -127, 37, 96, -53, 93, 41, 66, -68, 34, 11, -32, 120, 46, -98, -76, 112, 120, 83, 92, -101, 25, 55, -94, -128, -102, 104, 16, -74, -115, -11, 6, 100, -1, 120, 44, -114, -15, 116, -28, -29, 30, -78, -119, 37, 87, 32, -47, -57, 47, 51, 31, -36, 5, -93, -87, 57, 106, 26, 25, -28, -42, -55, -41, -80, 44, 24, 42, 83, 126, 96, 91, -103, -13, -90, -43, 42, 47, -104, -73, 88, -30, 58, 28, -10, 109, -53, 70, 69, 4, -116, 65, -118, -104, 89, 55, 79, -51, -10, 14, -50, -100, 4, -10, -62, -108, 75, 68, 70, 102, 31, -60, -65, 6, 105, -30, 127, 96, 119, 108, 82, 75, -56, 30, 99, -27, 28, -18, -117, 48, -5, -60, -39, 76, 85, 114, 88, 22, 69, -13, -81, 5, 63, 20, 126, -116, -125, 17, -16, -46, -86, -80, -80, 9, 15, 71, 83, -47, 61, -74, -117, -79, 107, 25, 62, -126, -104, -8, -78, 11, -102, 23, 95, -32, -112, -33, 34, -127, 25, -96, 46, 110, 63, 13, 59, 67, 10, -110, 61, 77, -102, -79, -58, 61, -25, -89, 90, 57, -122, -71, -90, 69, -63, -12, 94, -115, -70, -20, -36, 72, -20, -120, -19, 80, -96, -1, 28, 106, -108, -53, 44, 53, 20, -80, 10, 27, -87, 52, -26, -72, -43, 95, -113, 79, 108, 48, -78, -7, -68, -50, -5, -54, 56, -72, 97, 70, 94, 4, 12, -100, 31, 32, 86, 91, 102, -42, 14, 113, -14, 47, 61, -40, -16, -40, 55, 98, -94, -91, 61, 88, 124, -52, 116, -114, -9, -126, 122, 74, 118, -51, 123, -92, 113, -69, 24, -15, 48, 20, -71, 65, -84, 45, 88, -7, 57, 82, 67, 82, -53, -28, 90, 50, 14, 67, 68, 27, 70, 58, 82, -27, -13, -36, -52, 101, 74, -3, 126, 74, -40, -108, 79, 57, 98, 71, -16, -19, 67, -77, 9, 76, 34, 70, -20, 65, -114, -38, -75, -83, 68, -12, -10, -107, 17, 53, 71, -109, -6, -7, -47, -54, 47, 22, 77, 3, 3, -48, 18, 26, 103, 73, 20, 34, -13, 39, 33, 39, 30, 42, 44, -19, 6, 74, 1, -86, -128, 117, 103, -13, 71, -119, -97, -33, 0, -14, -20, -9, -29, 40, 34, -29, -32, -128, -62, 36, -28, 65, -74, -92, -48, 94, -79, -42, -50, 58, 108, -37, -128, 3, -16, 119, -90, 43, -10, -28, 38, 76, -17, 116, -31, 56, 118, 126, 12, 4, -1, 32, 81, 30, 30, -84, -10, 19, -51, 16, -105, 112, -51, -5, 4, 92, -112, -94, 1, -59, -127, -126, -76, -88, 92, 62, -100, 24, -78, -115, -67, 24, -91, 32, 43, 6, 96, 37, 12, 95, -43, -3, -52, 126, 5, -106, -19, -76, 5, 101, -52, -19, -120, 43, -123, -17, 63, -122, -45, -116, 37, -106, -91, -112, -6, -47, 114, 79, 76, 28, -100, 8, 40, -100, -99, -48, -83, -30, -11, 92, -43, 1, 76, 71, -84, -58, -102, -109, -79, -84, -34, 44, -44, 4, -42, 18, -94, -94, 57, -11, 51, 51, -66, 104, 53, -88, 105, 16, 84, -12, 99, 61, -80, -84, -127, -84, -95, -10, 50, -118, -44, -12, 124, -4, -3, -9, -22, 58, 3, 32, -17, -120, 6, -52, -28, -113, -53, -25, -98, 85, 115, 107, 104, 112, -118, 16, 41, 70, -87, -96, 33, 54, 5, -54, -101, 61, -5, 69, -69, 102, 37, 3, -7, 35, -49, -89, 127, 115, -24, -15, -16, -37, 47, -13, 93, 31, 115, 32, -8, -110, -56, 93, 51, -38, 107, 110, -106, 10, 68, 86, 84, -65, -65, 125, 37, -94, 21, 7, 38, -24, -6, -109, 110, -22, 28, -30, 103, 53, 56, 35, -47, -29, -1, -1, -114, 88, -20, -2, -63, -59, 39, 72, -61, 34, 31, -8, 98, 51, 116, 85, -22, -95, -43, -64, -105, 1, -53, -124, -98, -120, -128, -75, -37, -79, -124, 125, 107, 93, -44, -4, -73, 0, 124, -31, -40, 76, -45, 122, -62, 98, -21, -40, -3, -67, 71, 9, -52, -102, 80, -120, -105, -90, -93, 62, -83, 76, -76, 21, -115, -44, 35, -126, -86, -9, 12, -124, 52, -102, 42, 83, -79, -72, 93, 5, 107, -92, 11, -45, 96, -74, -30, 9, -87, -35, 68, -104, -20, 112, -91, -125, 39, -12, 42, -64, -24, 60, 53, -82, 70, 127, 17, -37, 45, -125, 109, -89, 71, 24, -9, 51, -1, -6, 106, 120, 57, -109, -70, -95, -108, -83, -106, 43, -99, 109, 123, 93, -90, 54, -32, 99, 66, -121, 73, 102, 25, 39, -77, -53, -87, 43, -5, -126, -116, 76, -114, 0, -54, -125, -15, 47, -48, -13, 100, -91, -79, -66, -25, 106, -40, 90, -83, 18, -94, 18, -55, 62, -119, -85, 24, 18, -26, 94, -36, 59, 16, 47, -5, 2, -91, 78, 9, 105, 77, 28, 10, 120, 33, 34, 22, 67, -59, -2, -119, 32, 110, 18, -121, 20, 10, -47, 63, 117, -43, 69, -37, 25, 34, 43, 101, -60, -115, -80, 114, -71, 96, 24, -73, 18, -4, 52, -11, 73, -16, 76, 7, 23, -61, -57, 93, 49, 59, -73, -25, -11, -122, 113, 52, 26, -14, -25, -89, -102, 72, 80, -98, -11, -62, -5, -94, 80, -69, -7, -109, 92, 19, -36, -100, -89, -26, -56, 90, 90, -67, 121, -67, -35, 39, -109, -59, -47, -15, 42, -50, -40, 68, 102, -106, 68, -61, -121, -108, 60, 118, 109, -113, 92, 12, 94, -111, -105, -28, 5, 90, -126, 30, 84, -40, 96, -40, -32, 71, 81, 75, 62, 88, 63, -121, 87, -88, -40, 83, 27, 25, 120, -103, 46, -92, 5, 71, 101, -59, 115, 13, 97, 1, 80, 87, 38, 47, 79, 111, 123, 14, 23, 124, 81, 107, -68, 83, 27, -77, -77, -42, -123, -6, -43, 28, -52, -71, -85, -80, 45, 0, -116, 51, 3, -30, 104, -75, 81, 12, 106, 51, 19, 95, 57, -29, 51, 70, 28, 86, -6, 113, 10, -112, -100, -60, -101, 51, 94, -36, -47, -108, -27, 16, 114, 104, 94, -66, 57, 40, -32, -70, 114, 107, 17, 66, 74, -121, 48, 11, -74, 110, -125, 2, -57, -54, -111, 88, 65, -1, -31, -1, -63, 69, -91, -32, 95, -101, -6, -111, 48, -48, -104, 110, 3, 95, -39, -119, -72, 6, -119, 23, -2, 21, 51, 63, -4, 93, -28, 71, 103, -119, -27, -98, 44, -81, 35, -16, -48, -7, 14, -52, 77, -87, -16, 46, -114, -98, 49, -91, 24, -125, -64, 42, 17, -4, 97, 34, 114, 72, -88, 75, -34, -36, -80, -63, 91, -16, 55, -29, -20, 58, -82, -38, -61, -4, 117, 96, 29, -8, -47, 68, -70, 78, -41, 82, -113, -59, -16, -51, 99, 44, 121, -128, 0, 24, 95, -49, 63, 12, -49, 83, 27, 30, 98, -97, -1, -11, -22, -65, 85, 97, -24, -45, 104, 124, -55, 64, -17, -42, 26, 56, -118, -18, -84, 30, -108, 67, 1, 99, -46, 16, -100, 75, -4, -15, 1, 40, -87, -64, 65, -84, -119, 45, -36, -26, -66, 59, 71, 103, -111, 112, 53, 113, -14, 20, -72, -56, 118, -63, -26, 45, -34, 111, -78, 40, -79, 0, 61, 113, -46, -107, 41, -72, 3, 55, -65, 54, 51, -11, 44, -126, -2, -117, -110, -52, 114, -72, -116, -58, 69, -94, -15, -2, 123, 73, 23, -70, 96, -108, -55, -39, 106, 68, 118, 61, -94, -55, -45, 62, 84, -82, 105, 6, -84, -49, 24, 106, -106, 95, 19, -95, -65, -20, 58, -119, -22, 64, 92, 56, -118, -50, 60, -13, 5, -96, -1, -21, -53, -91, -83, 68, 37, 75, 102, -80, 85, 16, 78, -35, 1, -63, -85, -7, 76, -121, 80, 10, 118, 67, -19, -5, 95, 36, 73, 30, -89, -115, 74, -39, -29, -118, -51, -112, -110, -13, 109, 92, -78, -125, 61, -32, 85, 18, 41, -90, 27, 91, 55, -114, 113, 0, 66, -5, -6, -52, 1, -121, -2, -43, -90, -66, 29, 36, -110, 28, 116, -127, -100, -76, -6, -7, 24, -77, 14, 114, 54, 101, 58, -29, -18, -17, 122, 22, -28, -83, 90, -26, -62, -106, -60, 4, -77, 31, 102, 34, -90, -105, 50, -12, 32, -66, 72, -77, 22, -53, 91, -82, -76, 5, 18, 64, 74, 124, -125, -1, -75, -78, -28, 39, -86, 57, 15, -115, -73, 73, 121, -111, -121, -127, 23, 125, -10, 13, 98, -101, 39, -37, -73, 58, -23, -123, 76, -116, 88, -48, 107, 124, -22, -1, -90, -34, -113, -110, -121, -53, 64, 14, 9, -126, 89, 26, -109, 44, 105, 120, 117, -59, 43, -126, 13, 55, 73, 126, -7, -5, 58, -109, 110, -4, -26, -15, -72, 79, 40, 65, -99, -9, 98, 59, -73, -89, -63, -110, 53, -44, 56, -48, -68, 59, -51, 56, -54, -81, -120, 54, -109, -105, 73, 54, 100, -10, -29, -103, 46, 109, 53, -24, 42, 32, 65, -45, -86, 57, 122, 98, -37, -117, 9, -36, 4, -69, -56, 28, -78, 3, 40, 81, -96, -109, 27, 62, -104, -58, -65, 68, 31, -85, 61, -24, -41, 19, 118, 79, 65, 68, 16, 74, -38, -18, 101, -68, 85, -113, -54, -126, -106, 121, 18, -51, 92, -79, 12, 12, -120, 124, 33, -50, -78, 80, 6, 43, 109, 122, 75, 70, -51, -110, -30, -122, 73, -72, -20, 4, -50, -1, -21, -34, 84, -67, 30, -28, -127, -128, -116, -2, -18, -1, -23, -123, -35, -69, -51, 38, 115, 123, 61, -4, 40, 100, 60, -49, 0, 7, -37, -47, 109, 82, 26, 24, -96, -74, -113, 100, -64, -19, 74, -24, 118, -66, -110, 77, -79, 8, -42, -28, 106, -5, 0, 81, -121, -29, 21, -121, -77, -56, -128, -77, -128, 125, -40, 22, 108, 41, -46, 16, 1, 69, -42, -89, -31, -31, -41, -14, 34, 118, 78, -49, -36, -89, -14, 26, -95, 70, -118, 2, 52, 10, -116, 61, 9, -61, -80, 82, 57, 67, -18, 64, 14, -23, -106, 112, 124, 121, 18, 112, 81, 66, 2, 18, -49, 19, -8, 14, -69, -7, 16, -78, -121, 59, 74, 55, -91, 53, 71, -46, 49, 121, -91, 125, -82, 106, -41, -20, 80, 112, -51, 107, -56, 74, 39, 75, 113, 89, -54, 15, -16, -3, 118, 105, -33, -5, 44, -37, 105, -39, 96, -45, 49, 37, -14, -45, 113, -71, 41, -45, 59, 66, 41, -117, 55, 0, 51, 16, 107, -2, -119, -27, 114, 59, -19, -33, 117, -65, 52, 83, -94, -62, -99, -6, -96, 117, 85, 2, 34, -124, 97, 49, -119, -100, 71, -42, -29, 68, -128, -42, 108, -128, -92, -29, -46, -30, 37, -69, -10, -41, -47, -15, 59, 78, -44, 26, -58, 78, -69, 124, 69, 105, -69, 24, -24, -18, 79, 113, 50, -113, -13, -75, 92, -21, 89, 17, -40, 20, 73, 41, -53, -111, -117, 126, -33, 104, 25, -69, 14, -38, 83, 111, 88, -94, 7, 111, -58, -37, 64, -34, 59, 90, 45, -108, 29, -107, 16, 48, -84, -76, 1, 35, 65, 16, -11, -86, 65, 41, -124, -75, -91, -19, 17, 40, 81, -53, 40, 0, 121, -46, 121, -97, -37, 58, 70, 51, -67, 123, 75, 78, 6, 50, -33, -54, -106, 105, 21, -59, -24, 67, -58, 34, -19, -54, 33, 92, -104, -39, 127, 48, -83, -25, 66, -126, -58, 35, -72, 39, 6, 90, -96, 110, -37, 55, -16, -115, 63, -92, 87, 31, -124, 80, -44, 22, 99, 63, 24, 53, -10, 122, -33, -103, -8, -119, 67, -20, -63, -3, 120, 63, -36, -86, -47, -83, -110, -46, -28, 118, 25, -13, 19, 37, -58, -55, 48, 125, 34, 42, 83, -117, 39, -96, 78, -23, -70, 84, -91, 88, 3, -98, -123, -106, -125, 71, 71, -8, -115, 21, -109, -115, -54, 100, -44, -44, -114, 93, -114, -42, 1, -77, -16, -94, 65, 39, -101, 14, 12, -36, -92, 91, -71, 80, 119, -42, 86, -126, -44, 110, -16, 85, 49, 125, -44, 60, -60, 78, -27, 79, -74, 3, -43, 7, 60, -73, 117, -42, 109, 66, 68, 41, 70, -45, -66, -21, 4, 38, -52, 68, -104, -71, 6, -22, 78, -33, -74, 77, 123, -94, 37, 121, -128, -37, 127, -102, -103, -37, -95, -78, -28, -119, 1, -22, 19, -34, 123, 94, 84, -30, 28, -55, 2, -110, -17, 13, 41, -19, -62, -72, -42, 126, 120, -57, 19, 121, 82, 63, 115, 35, -11, 71, -63, 109, -36, -33, -124, 122, 47, -36, 14, -122, -96, 89, 118, -69, -80, -64, -43, -35, -70, -32, -86, 24, 12, -91, 5, 100, -62, 75, 86, -22, 74, 43, 6, -125, 48, 4, 117, 57, 19, 28, -15, 43, 99, -116, 37, -66, -41, -82, 20, -50, 24, -93, -11, -63, 41, -16, 9, 81, 118, -82, -88, 59, 101, -15, 90, 104, -6, -74, 39, -29, -83, -24, -31, -71, -12, -68, 125, 112, 77, 17, -105, 4, -127, 63, 60, 56, 57, -53, -47, 72, 105, -110, -121, 64, -100, -99, 79, -100, 30, 12, -76, -25, -48, 110, -94, -61, -76, -60, 100, 63, 86, 104, -104, -88, -89, 82, -65, 30, 34, 31, -120, -126, 76, 62, 56, 3, -59, 42, -31, -43, -24, -98, -32, -25, -83, -66, 26, -96, -76, 73, -70, 25, -101, -94, -66, -110, -61, 28, -22, 118, -72, 120, -14, 33, -49, 60, -58, -120, 44, 57, -65, -23, 120, -91, 27, -46, -76, -94, -20, -10, 48, 101, -59, 55, 93, 119, -70, -122, -6, -28, 35, 98, 123, 41, -100, -73, 22, -77, -82, -60, -31, -70, 43, 53, 77, -106, 88, 82, 88, 52, -30, 113, -50, -123, 43, -9, -116, -26, 122, -75, 114, 52, 44, -54, 40, -112, -49, -12, 116, -82, 81, 126, 66, 126, 123, 124, -66, 33, 8, -5, -37, 31, -27, 14, -98, -73, 69, 75, -110, -100, 113, -68, 46, -25, -49, 3, -120, 84, -71, 25, -50, -93, 100, 49, -17, -23, -21, 72, -1, 45, 55, -112, -107, 82, -105, -45, 106, 23, 52, -128, -35, 15, 103, 124, 20, 62, -30, 49, 52, -94, -84, 94, -73, -127, 53, 54, 73, -31, 17, 46, 61, -63, 29, -84, -53, 17, -104, 25, 6, 14, 28, -57, -120, 70, 93, 105, 36, 118, -70, 32, -84, 123, 53, -71, -112, -87, 105, 61, 37, 70, 126, 55, -78, 30, -60, 72, -103, -48, -66, 30, -1, -116, -1, 2, 71, -8, -91, 90, 83, 114, 12, 53, 82, 26, 27, 98, -102, -109, -93, 54, 65, 89, -90, 49, -73, 73, -38, 102, 108, -86, 24, -123, -2, -89, -54, -41, 8, 104, -86, 66, 104, -95, -58, -84, 1, 62, 64, -93, 125, -119, 65, -46, -90, 106, 64, 50, 36, 96, -96, -59, 39, 2, 77, -22, 43, -118, 18, 119, 96, 14, 115, -62, -61, -70, 74, 83, 2, -123, 44, 3, -119, 8, -43, -4, 72, -50, -111, 68, 1, -44, 2, -18, 65, 75, -99, -99, 102, -110, -8, -20, -116, 21, -83, 118, -97, -71, 74, -85, 98, 42, 60, -5, 122, -123, 101, -94, -55, 41, 25, -13, 64, -115, 71, 118, -10, -121, 127, -96, 43, -70, -100, -126, 29, -11, -125, -82, 117, -63, 122, -40, 121, -18, 69, 52, 92, 71, -89, -35, -120, 54, -54, -79, -84, 64, 60, -106, -126, -24, 123, 37, 18, 46, -101, 79, 47, 54, 54, -96, 64, -39, -28, -100, 27, -8, -85, 117, 55, 93, -19, -46, -61, -42, -96, 118, -86, -31, -23, 108, -10, 36, 4, -123, 12, -60, -6, 39, -109, 90, 12, -42, 108, -19, -68, -9, -44, 74, -110, 53, 116, 16, -17, -116, 61, 24, 93, 116, 74, 74, 53, 67, -83, -89, -32, -8, -113, 15, -25, 77, 58, 93, -103, 75, 119, -125, -19, -86, 103, -73, -40, -26, -70, -109, -110, 50, 109, -87, -37, 105, 31, -126, 93, -25, 2, 84, -103, -80, -128, -120, 55, -127, 96, -68, -16, 92, 71, 29, 98, 77, 55, 125, 24, -90, -23, -119, -97, 52, -38, 50, -127, -12, 8, 46, 82, -69, 95, -109, -18, 58, 10, -36, 72, -60, 59, -40, -90, 103, 27, -38, 79, 116, 16, -31, -102, -82, -106, -23, -123, 47, 4, -4, 70, 15, 71, 31, 53, -39, -90, -89, 77, 99, -33, -43, -15, 125, -20, -14, 99, 9, 67, -123, -119, -12, -82, 84, 105, -40, -5, -62, -67, -120, -107, -21, 80, 106, -60, -65, 61, 36, -72, 69, 126, -121, 39, 46, -34, 73, -65, 75, 46, 21, 17, -106, 124, 25, -6, 81, 65, 83, -116, -79, -72, -107, 35, 38, -62, 76, -52, -75, -87, 40, 38, 77, 71, 14, -86, 127, 86, 116, -104, 16, -39, 93, 70, -62, -7, -51, 98, 30, 73, 77, -22, 82, 99, 8, -108, 7, 19, 62, 44, -68, 1, 30, 54, -90, -21, -2, 113, -54, 66, -114, -71, -116, -55, -19, -85, 39, 92, 82, 102, -58, 4, 96, 49, -46, -117, -38, 79, 5, -22, 26, 102, -64, -78, -59, -25, 83, 42, -41, -120, -26, 61, -9, -46, 113, -2, -1, -113, -23, -53, 66, -2, -102, -115, 39, 30, -84, 91, 86, 50, 6, -78, 25, 99, 82, 56, -107, 53, 119, 111, 108, -78, 51, -75, 123, -118, 43, 86, -77, -36, 45, -34, 84, 90, 68, -127, 101, 112, 77, -125, 81, 57, 25, 116, -25, -11, -8, 54, -51, -126, 74, 10, 118, 1, 125, -77, -40, 11, 114, -65, 23, 89, -42, 8, -126, -94, -91, -60, -47, 43, -41, 100, -90, -75, -121, -68, -115, 37, 37, 127, 66, -46, 96, -28, 105, -82, -52, 109, -71, 78, 44, 0, -62, -28, 48, -65, -31, 105, 111, 57, 44, 35, -7, 126, 119, 20, 96, 51, -85, 96, -106, -29, -35, 116, -113, -56, 111, 108, 91, 46, -75, -17, 27, -72, -98, 22, 20, -103, -20, -110, -86, -127, -46, 24, -62, -110, 40, 81, 96, -64, 19, 18, -14, -113, 7, -61, 46, -112, -81, -77, 83, 68, 21, -18, -70, 29, 34, 98, -108, -118, 18, 56, 69, -59, -25, -10, -119, -64, -104, 37, 80, 10, 73, -104, 7, 120, -94, 8, -84, -89, 120, -8, -1, 30, -79, -74, 78, -36, 123, 83, -95, -108, -98, 55, -38, 59, -122, -21, 83, -58, -94, 16, 60, -50, -42, -20, 36, -113, 63, 94, 125, -26, 21, 61, -56, 62, -7, 45, 93, 100, -48, -16, -32, 121, 23, 120, -37, 55, -82, -93, 72, -4, -56, -21, -13, -61, -55, -116, -62, -123, -43, 67, 7, -41, 18, -14, 126, 63, 79, -35, -115, 92, -79, -100, -53, -9, -106, -11, 49, 30, -3, 87, -24, 113, 110, 11, -64, -103, 78, -80, -2, 59, 73, -108, -18, 25, -87, 7, 19, 10, 6, -112, -116, -24, 57, 56, -71, -118, -69, -18, -107, 56, 16, -43, -57, 98, -111, -123, 19, 56, 96, -102, 70, -94, -13, -19, -122, -74, 104, 64, -24, -110, 72, -54, -28, -84, 17, 97, 89, 75, 85, -59, 13, 84, -9, -15, 100, 100, 5, 8, -18, 14, 2, 58, -16, -73, 69, 75, 21, 70, -118, 65, -89, 108, 68, -69, -63, -18, -82, -128, -81, 26, 67, -99, -12, 126, -91, 117, 50, 93, 5, -20, 41, 58, 121, -35, -115, -99, 31, 107, -3, -121, 90, -19, -32, 36, -89, 117, -102, 93, -62, -19, 4, -30, 10, 4, -49, -48, 40, -64, 42, -5, 14, 125, -90, -27, 52, 42, -95, -69, 97, 17, 110, -96, -112, -21, -117, -91, 26, 22, 25, -19, -35, -79, 65, -68, -57, 70, -18, 20, 126, -60, -58, 78, -72, 99, 39, 41, -60, 10, 101, -119, 118, -21, 97, 4, 27, -14, -43, -60, -86, -5, 8, 60, 118, 56, -123, -1, 88, 73, 6, 23, -67, 111, -26, 12, 114, -14, 8, -44, 84, 126, -33, 41, -107, 10, -125, -112, -63, -17, 8, 113, 44, -4, -48, -86, 56, -49, -27, -105, -23, 47, 38, 9, 124, -113, -97, -111, -8, 72, 101, 6, -53, -78, 88, -47, -124, 27, -65, 34, -75, -80, 69, 22, -45, -3, 84, 29, -71, -29, -14, -105, 4, -96, 48, 2, 103, 74, -103, 96, 35, -114, 43, 98, 47, -115, -10, 44, -27, -98, 50, -77, 91, -109, -87, 97, 72, -93, 114, -2, 96, 125, -108, -20, -66, -24, -31, -110, -81, -35, 49, 24, -10, 52, 78, -115, -29, -33, -82, -9, -46, 38, 105, 59, 101, 9, -80, -123, -77, 117, 46, 120, 66, 22, -5, 15, -53, 112, -1, -111, 36, 122, 84, 69, 96, -30, -60, -32, 53, -37, 101, -33, 72, -27, 113, 121, -15, 37, 105, 95, 93, -73, 78, 92, 66, 109, -2, -115, -74, -57, 66, -52, 18, -67, -117, 103, 49, 73, 118, -29, 81, 125, 77, 67, -127, 54, -29, -88, -81, -69, 48, -40, -59, 5, -103, -39, 27, 81, -30, -59, -49, 66, 36, -17, 121, -92, -39, 49, -46, -108, -52, -63, -52, 48, -52, 107, 10, 39, 80, 121, -88, -39, 40, 6, -123, 25, 66, -56, 84, 33, 60, -96, -125, -95, -16, 107, -101, 8, 125, 4, -59, 85, -113, 101, 44, -81, 127, -128, 60, 112, 66, 59, 91, 90, -116, 87, -80, 61, -119, -99, -41, 115, -43, 111, -83, -60, 122, 14, 13, -82, 18, -91, -110, 114, -57, -23, -111, -104, -58, -70, 42, -31, 63, -17, -106, -69, 94, -113, -39, -72, 103, -108, -61, -100, -60, 69, 56, 63, -49, -24, -45, -79, -82, 97, -44, 68, 37, -91, 37, 34, -79, -49, -48, -79, 28, -114, -111, -54, 86, 122, -128, 55, 16, 27, -20, 11, -21, 69, -110, -78, -74, -23, -27, -8, -105, 119, -121, 39, -48, 50, -15, -10, 0, 42, 123, -24, -33, 13, 39, -90, -31, 82, 85, 14, 15, -42, 45, -51, 20, -41, -105, 102, 4, 55, -84, -25, 38, 34, 120, 60, 47, -122, -29, -112, 62, -55, -2, -1, 101, -59, -52, -7, -8, -93, -102, 116, -26, -111, -21, -11, 110, -124, -20, 26, 105, 75, 42, 98, 46, 118, 41, -97, 46, 71, -113, -24, -12, -43, 30, 50, -16, 89, -54, -40, 122, 114, 104, -123, -117, -114, 13, -75, 126, -40, 67, -75, -1, 54, -80, -82, -114, -56, -32, 127, -83, -34, -54, -104, 20, -49, -29, 105, 76, 33, -76, -123, -19, 73, -66, -101, -78, 16, -52, 9, -127, 25, -37, -117, 127, 89, 17, 94, 113, 65, 97, 117, 99, -52, -78, 15, 116, 28, 59, -48, 122, 17, -46, 124, 86, 48, -93, -73, -38, 91, 103, -62, -42, 0, -63, -7, -94, 19, -92, -15, 98, 44, -56, -6, -86, 76, -103, 124, 119, 68, 93, -93, 48, -37, -12, 28, 37, 54, 40, 59, -110, -25, 8, 8, -77, 24, -80, 12, -11, 4, 1, 80, -113, -53, -110, 76, 86, -119, -94, -35, 94, 50, 112, -13, 4, 101, 83, -63, -74, -17, -71, -118, 74, 85, 31, 6, -56, -87, -77, -103, 68, -27, 43, 127, -53, 96, -62, 71, 49, -4, -40, -63, 125, 13, 70, -117, -100, -108, 96, -117, -50, 89, -84, 118, -53, -109, -64, -90, -42, -80, 70, 53, 71, -3, -113, -17, -37, -122, 40, -124, 38, 41, -70, -30, 125, -114, 10, -105, 123, 84, -99, 114, -13, 32, 109, 104, 83, -37, -87, -62, -105, 91, 127, 71, -5, 11, 67, 121, -88, 117, 32, -65, -98, 90, -106, -31, 24, -8, -4, -6, -27, -1, -61, -17, -127, 114, -35, 1, 6, -64, -98, 126, -16, 52, 82, 57, 51, -100, -25, 5, 45, 95, 71, 40, -84, 77, 44, -76, -52, -33, -121, -88, -70, -105, 48, 67, 39, -12, -34, 39, 20, 12, 49, 65, -14, -107, -1, -116, -104, -86, 70, -6, -82, -62, 79, 68, -85, 19, -61, 4, 8, -111, 20, -74, -83, 34, 123, 126, 73, -68, 32, 74, 44, 107, 87, -60, 20, -73, -51, -80, 88, 86, 32, 24, 30, -76, 125, 24, 56, 105, 7, 60, -81, -38, 53, -69, -83, 51, 6, -114, -122, -114, 27, 68, -99, -105, -95, -64, -3, -48, -78, 87, -37, 34, 49, 120, -115, 82, 0, -49, -86, 25, -62, 6, 43, 9, 120, 31, 84, 118, -75, -111, -14, 66, -61, 94, 3, -33, -26, 113, 64, -6, -100, -122, -6, -71, -91, -96, -26, -25, -125, -55, 94, -16, -44, 70, -16, 90, 69, 125, 125, 9, 50, 37, -113, -13, -96, 35, 85, 19, -44, -60, 16, 87, -4, 48, 52, -67, 111, 15, -119, -47, 25, 106, 37, 8, 52, -23, 120, 46, 51, 10, 96, -27, 111, -111, -97, -2, 113, 106, 50, -80, 106, -91, 92, -52, -13, -3, -103, -42, 41, 95, -31, 80, -22, -27, 20, 36, -5, 87, -24, -43, 9, -61, -40, 64, -96, 82, 5, 42, -89, 23, 17, -33, 111, 88, -128, -95, -15, 109, 47, 7, 4, -127, -63, -86, 78, -87, 14, 54, 81, 110, 25, 77, 27, -111, 105, 81, 86, 81, -123, 53, -121, -106, 29, 111, 74, -66, -19, 119, -40, -70, 68, -21, -39, -33, 49, 85, 15, -13, 9, -24, -105, -86, -48, -116, 127, -13, 67, 15, -33, -104, 34, 122, -26, 7, -99, 99, -25, -73, 52, -6, -47, 91, -1, -28, 67, 22, -128, -109, -20, -75, 54, 105, -34, 84, -5, 111, 110, -41, 95, 27, 73, 116, 9, -58, -5, 61, -80, 70, 59, 122, 44, -90, -121, 33, 53, -96, 1, 57, -31, -11, 73, -97, -68, -113, -47, -110, -85, -100, 6, 127, -4, 71, 84, -21, -7, -8, 36, 67, 119, -38, -95, -122, -84, -110, -89, 0, -51, 52, 46, -63, -88, -32, 47, -40, -24, 55, 80, 118, 67, 77, -61, 53, 83, 45, -17, 23, -72, -119, 87, -55, 82, 78, -96, -86, 73, 0, 33, -108, -121, 62, 5, 41, -92, 17, 94, 112, -14, -84, 77, 25, 94, -101, -8, -59, -43, -31, -60, 25, -115, -35, 70, -23, -57, 83, -74, -52, -54, 125, -124, 1, 77, -70, -81, -31, -72, -115, -63, 126, -86, -49, 46, -115, 9, -95, -61, -86, -104, 98, -49, 3, -61, -68, -90, 67, -118, -74, 116, -33, -22, 36, -109, -50, 44, -87, -58, 94, -81, 95, 123, -123, -68, 70, -17, 110, -47, 47, -105, -52, -12, 0, 118, 43, 110, -92, 104, -16, -56, 10, -103, 38, 16, -78, 112, -17, 29, -2, 95, -15, 14, -9, -3, 19, 115, 83, -80, -68, 13, -50, -125, -2, -109, 35, -56, 37, -44, 82, -117, 38, 36, 103, -43, 5, -74, 86, 92, -14, 37, -57, 56, 94, 7, 96, -45, -97, -87, 10, 80, 116, 74, -96, -8, 81, 52, -51, -92, -120, -23, 50, -45, 127, 66, -25, 14, -78, -29, -106, -58, -1, -126, 100, -74, 85, 3, -106, -20, -28, 7, -49, 112, 51, -38, -92, -60, -38, -58, -9, 24, -21, 82, -83, 121, 19, 86, -113, 79, 127, -80, 108, 49, -66, -7, 46, -2, -17, -89, -109, -13, -88, -34, 41, 53, 30, -8, -82, -67, -113, 51, -98, 65, -117, 25, -106, 94, 118, -22, 43, 30, -49, 126, 58, -86, -13, -117, 84, 64, 72, 56, -104, -102, 60, 40, 43, 20, -63, 13, -14, -82, -36, 34, 41, 49, -41, -97, -33, -67, 55, -108, -1, 67, 26, -28, -111, -62, 113, 118, -123, 23, 84, -3, 72, 18, -125, 124, 99, -54, 85, -81, -112, 114, -51, -68, -106, -73, -15, -111, -124, 121, 122, 97, 37, -81, -42, -59, 109, 31, 90, 127, 4, -25, 60, -37, -80, 61, -92, -28, 114, 4, -107, -94, -115, -28, -39, 23, -98, -18, -27, -121, 68, 36, 87, 24, -69, 3, 93, 78, 120, 100, -80, 116, -76, -119, 23, -27, 82, -94, -46, 16, 14, 24, 36, -120, -9, 84, -70, -36, 123, 19, 46, 73, 2, 94, -57, 97, -37, 42, -98, 91, -47, -41, -85, 109, -80, -83, -31, 58, 65, 125, -62, -56, -103, 103, 44, -79, 80, 125, 94, -89, 109, 112, 37, -29, -6, -89, 12, -16, 104, -49, -119, -37, -33, 111, -6, -3, 111, -18, 33, -63, -99, -38, 39, 29, 83, 13, 103, 114, 68, -41, 117, -12, -100, 32, 121, -43, 101, -76, -50, -96, 97, 61, 68, 78, -86, -43, -23, 53, 11, -74, 97, -101, -72, 44, 27, -106, 27, -107, 70, 98, 64, -54, 58, 58, 83, 1, 53, -52, 6, -25, -30, -5, -42, 78, -96, -98, -78, -90, 108, 25, -102, -75, 42, 52, 126, -36, 80, 126, 24, -105, -97, 78, -113, 81, 93, -35, 47, 115, -86, -79, 104, 78, 61, -38, 52, 39, 82, 76, -44, 57, 66, -99, 68, -111, -48, 112, 66, -19, -102, -126, -80, -102, -28, 103, -95, 104, -88, 75, 106, -52, 28, -53, -44, -125, -15, -104, 99, 62, 106, 56, 93, 59, -15, -121, -101, 114, -97, -107, -90, 61, 63, 93, 76, -29, -51, 11, -121, 43, -128, 54, 108, -47, -75, 56, 71, -121, -6, -10, 43, -114, 85, -103, -62, -25, 80, -63, 121, 127, -37, 112, -7, 86, -122, -112, 14, -41, -9, 63, -23, 48, -86, -45, 69, 31, 4, 119, 96, -117, 109, -82, 100, 122, 65, 44, 9, 74, 100, 13, 69, -59, 53, 87, 74, 18, -119, -57, -36, -111, 96, 6, -118, -37, -10, -61, -116, 94, 77, -116, -35, 24, 41, 67, -63, -49, 29, 7, -125, -23, -42, -102, 29, 52, -90, -102, -4, -115, 118, -34, 90, -123, -71, 108, -103, -115, 69, -44, -20, 59, 80, 29, 41, -108, -125, -9, -73, 85, -94, 28, -4, -32, 26, 87, -20, -128, -127, 30, 52, 8, 63, -58, 1, -66, -29, 83, 109, -125, -5, -44, -110, 46, -96, 7, -61, 97, -73, -69, -105, -73, -94, -103, -124, 116, -12, 22, -55, -69, 73, -15, -6, -38, -65, 108, -61, -25, 115, 81, -109, -90, 108, -72, -75, -127, 119, -114, -116, 82, 50, -42, -118, 95, 49, -76, 124, 48, -70, -111, -55, -49, 71, 79, 71, -120, 75, -126, -10, -85, 112, -4, 112, -96, -113, -101, 125, -100, 113, 55, 79, 22, 13, 35, -46, 107, -90, 50, 38, -97, -100, 29, 70, 125, 6, -110, 108, 102, -91, -30, 73, 93, 119, -8, 114, -48, -63, 103, 46, 59, -72, 90, -70, 127, 12, -43, 16, -41, 25, -28, -110, 85, -63, 32, 114, 82, -36, 68, -22, -28, -34, 9, -94, -6, -104, -7, -41, 93, 26, 45, -4, 21, -104, -79, -32, -86, 59, 92, -80, 49, 115, -106, 26, 115, -26, 72, -105, -123, -61, -89, -39, 46, -48, -46, 96, 75, 69, 93, -81, 104, 95, -26, -89, 13, 1, 39, -94, 21, 97, 86, -10, 115, -126, -100, -79, -8, -14, 48, -73, -12, -128, 76, -125, -116, -32, 113, -120, 86, -86, 20, -19, 17, 86, 109, 76, 37, 87, -106, 93, 97, -113, -54, -84, 61, 6, -20, 58, -111, -8, 103, 112, 49, 66, 58, 110, -102, 68, 94, 9, 49, -50, -48, -75, -56, 103, -108, 20, 34, 108, 39, 14, -112, 73, 55, 68, 57, -117, -65, 53, -72, 106, -4, -57, -12, -14, 90, -50, -94, -64, 12, 73, 121, -87, 30, 53, -38, -94, -8, -61, 116, 125, -32, -11, -33, -52, -101, -2, 43, 58, 21, -106, 25, 55, 118, -87, -113, 77, -92, 63, 17, 127, -80, 15, -44, 16, 107, -34, 38, -15, -108, 26, -12, 45, 109, 94, 103, -91, -81, -57, -38, -70, 34, 9, -120, -19, -25, 76, -55, 9, 114, 81, -61, 52, 14, 104, -15, 32, 11, -20, -9, 119, -98, -66, -31, -96, -12, -24, 21, -58, 98, 106, -5, -74, -55, 71, 17, 43, -73, -25, 100, 22, -79, -1, -10, 127, 76, 58, -123, 58, -44, 61, 85, -24, 86, -120, -70, -112, 117, 8, 23, 81, 45, -29, 124, 99, 20, -35, -32, -61, 95, 74, -23, -47, -39, 71, 109, 13, 66, -18, -29, 70, 59, -20, 63, 121, -91, 34, 82, -126, -41, -34, 105, -107, -95, 85, -22, -88, -124, 24, 60, -54, -6, -48, 108, 2, 55, 49, 59, 74, 126, -53, 25, 88, -127, 69, 32, 7, 92, 54, -26, 85, 105, 93, 56, -29, 93, 47, -35, 29, 29, -85, -55, 20, 40, -84, 66, -50, -76, 64, -63, -19, -103, 85, 103, 116, 78, -78, 75, -53, 99, 37, -127, -25, 109, 35, 58, 4, 32, 44, -1, -79, -15, -9, 24, 35, -55, -18, -114, -34, -28, -111, 34, 59, 22, -58, -88, -127, -82, 84, -81, -36, 64, -86, 92, -31, 54, 57, -54, -96, 112, 76, 39, 31, -121, 73, 52, -115, -63, 52, 58, -82, 35, -119, 61, 76, -46, 97, 76, 23, -91, -77, 68, 66, 80, -28, 42, -83, -110, -94, -65, -99, -98, -2, 78, 54, 108, -106, 99, 82, 75, 50, -117, -36, -51, 119, 70, -29, 15, -49, -38, 32, 27, 86, 75, -5, -52, 27, 49, 46, 9, 12, 53, 12, -87, 64, 37, 110, 16, -122, 75, 123, -122, 92, -38, -26, 109, 35, -88, 35, 116, -59, 7, 120, -116, 103, -91, 16, 21, 121, -118, 117, 92, 101, 100, 114, 16, -77, -69, -66, -53, 30, 99, -7, 7, -123, -11, 17, 16, 69, -6, 125, -39, -13, 63, -79, 82, 43, -114, 26, 5, -70, -40, -120, 39, 109, 8, -11, -59, -30, 3, -89, -107, -54, -84, 11, 46, 41, -14, 85, 1, 116, 108, 43, -94, -6, 88, 63, -107, 93, 82, -70, -94, -92, 73, -50, 112, 55, -3, -26, -114, -79, 32, -56, 111, -90, 0, -82, 25, -86, -12, 43, 92, 51, 23, 84, 105, -2, -59, -100, 3, 107, 50, 5, 2, -74, 3, 111, -7, 52, 90, 32, 81, -80, 47, -51, 40, 124, -76, 56, -23, -70, -17, 49, -69, 12, 45, 70, 53, -3, 74, -11, -4, -7, 91, 126, -98, -89, -68, -3, -57, -79, -5, -21, 60, -105, 40, 4, 47, 121, -82, 117, 83, 73, 64, -126, 121, 67, 77, 4, 7, 33, -87, 21, 78, -30, 97, -51, 103, -39, -97, -55, -70, -33, -58, 60, -3, 42, 112, -41, -9, -16, 9, -31, -5, -29, 84, -120, -24, -121, 42, 20, -78, -73, -118, 47, 115, -105, -40, -82, 47, -93, 50, -114, 81, -107, 25, 1, -13, -118, 68, -1, -29, 100, -112, -71, -119, 80, 88, 90, -31, 80, -68, 75, -7, -85, 86, 7, 9, -88, 56, 2, -64, -1, -6, -73, -5, -91, 46, 44, -91, -49, -37, 42, -50, 121, -88, -40, -8, 58, 33, 90, -51, 67, 64, 34, -43, -39, 63, -106, -119, 78, -60, 101, -78, -33, -71, -72, 127, -82, 82, -68, 4, 117, 41, -65, 97, -110, 35, -25, -5, 95, 56, -72, -37, -39, 85, -108, 16, -96, 99, -8, -52, -92, -49, -13, -27, 7, -75, 25, -80, -58, -112, 50, -45, 112, -120, -55, 50, 29, 13, -108, 99, -119, -17, -115, -31, -9, -128, 87, 42, -90, 82, -34, -37, 43, 87, 55, -124, -48, 67, 83, -112, 10, -128, 15, -41, 52, -117, -122, 21, 60, -125, 82, 20, 64, 0, -58, 56, 109, -97, -101, -41, -67, 35, -64, -58, -81, -41, -62, 124, 15, 10, -123, -14, 63, -96, 25, -128, -33, -117, -84, -49, -85, -68, -113, 68, 58, -73, -28, 60, -100, -79, -65, -98, -38, -74, -53, -101, -100, 107, 31, 53, -63, 12, 39, -98, -109, 40, -78, -117, 126, -80, 66, -36, -64, 25, -15, 86, -16, 116, -19, -40, -104, 95, 45, -23, -98, 107, -75, 96, -76, -55, 61, 115, -3, -1, -89, 124, 51, -74, 18, -31, -81, -105, 58, -100, -126, -123, -118, -24, -42, 38, -120, -37, -121, -4, 62, 36, 111, -117, -24, 103, 40, -39, 119, 112, -127, -111, -58, -120, 46, 82, -126, -40, -89, -117, -9, 80, 75, -70, -89, 108, -75, -25, 70, -86, 79, -27, -61, 113, 96, 29, -45, -77, -73, 78, -31, -106, 92, 25, -29, 18, -56, -112, 87, 114, 103, 51, -86, -18, -109, 101, -9, 69, 6, -95, -1, 109, -37, 83, 117, -77, -32, 64, 16, 46, 108, -115, -10, 104, -127, -21, -35, 2, 30, -56, -38, -119, 2, 88, -12, 16, -12, -52, 89, 29, -34, -87, 120, -65, -51, 12, -4, -25, 0, 40, 21, -54, -85, -74, -58, 9, -91, -100, 52, 92, -111, -107, -29, 119, -15, 65, -87, 5, -45, -73, 55, -126, 35, 42, 8, -125, -123, 59, 76, 117, 72, 23, -73, 60, 96, -56, -92, 52, -15, 124, 92, -111, -88, 82, 117, 112, -31, -59, -59, -104, 87, -100, -100, 95, -11, 45, -112, -76, 2, -80, 114, 88, 114, -46, 103, 92, 48, -64, 21, 63, -27, 79, -47, 100, 57, -118, -27, 103, 96, -2, -100, -100, 71, 127, -80, 76, 10, -3, -77, -84, 126, 2, -68, -122, -27, 123, 4, -19, -31, 78, 111, 33, 37, -112, -33, 44, -22, 104, -23, -101, 76, 115, 32, 24, 40, -122, -18, 85, -1, -115, 96, 11, 118, -39, -44, -97, 87, 92, -44, -65, -60, -105, -52, -68, -84, -95, 57, -123, 67, 57, -127, -37, 95, 60, -56, 42, 43, 9, -46, -85, 55, 32, 74, 68, -116, 25, 54, -40, 0, -63, 3, 46, -83, -128, 40, 9, -24, -15, -45, 1, 104, 39, -58, -8, 52, -121, -36, -68, 19, -39, -117, -92, -75, 1, 20, -18, 14, -39, 23, 62, 107, -92, -123, -59, -82, 106, -4, 79, -127, -48, 39, -17, -81, -95, -27, -73, 67, 3, -67, -122, -16, -126, 94, -103, 83, -88, 59, 89, -76, -91, -83, -109, 47, -49, 121, -30, -83, -78, 7, 101, -84, 3, -114, 76, 59, -105, 75, -32, 47, -114, -59, 38, -39, 12, -24, -14, 15, 75, -10, -93, 116, -89, -47, -92, -37, -80, 120, 110, -80, 85, 16, 108, -33, 39, 5, -56, 24, -69, -64, -61, -47, 83, 31, 41, -12, -81, 65, -53, 70, 103, -36, -68, -7, 26, 123, 30, 91, -45, -52, 60, 39, -49, 121, 2, 76, 81, -85, 60, 16, 113, -34, -122, 77, -23, 75, 8, 90, 75, 31, -37, -64, -45, -124, -121, 33, -90, 3, 80, -72, 60, 23, 20, -5, -21, -47, -36, -120, 90, 117, -95, 93, 126, -126, -73, 81, -103, 46, 76, 105, -29, -88, -125, 31, 114, -85, 87, -125, 33, 57, 39, 49, -104, -47, -32, 4, 67, -18, 53, 73, 57, 95, 45, 28, 39, 74, 34, 30, 38, -17, 72, -97, 108, -42, 45, 5, -123, -1, -102, -124, -62, 9, 75, -127, 62, 29, -13, 28, -36, 34, 38, -87, 81, -20, -13, -19, 126, 103, 80, 53, 48, 78, 57, -118, 115, 74, -4, -40, 4, 62, 111, -49, 75, 36, 117, -4, 7, 25, -34, 23, 7, 112, -111, 10, -85, -42, -97, 93, -17, 28, 58, 113, -44, -111, -100, 30, 120, -2, -12, -17, 88, 24, -102, 114, 29, 39, -15, 38, 119, -126, 108, -31, -122, -117, 45, 104, 30, -118, 53, 118, 106, -43, 56, 58, 114, -113, 44, -102, 32, 22, 66, 33, 122, -118, 72, 101, -63, 76, -25, -26, -2, -45, -45, 101, 84, -56, -124, 115, -16, 19, -93, -116, 83, -123, 76, 4, 7, 1, 110, 31, -48, -18, 112, 80, 89, 42, 45, 42, -100, -8, -9, 59, -124, 108, -116, 109, 61, -16, 74, -30, -29, -82, -58, -60, 17, 70, -110, -47, -43, 120, 99, 32, 41, -16, 125, -102, -128, 68, 101, 99, -65, 111, -93, -99, 113, -48, -9, 67, 123, -30, -97, -5, 76, -97, -33, -99, -43, -102, 57, -22, -126, 88, -88, 48, -113, -75, 12, -39, 68, 31, -108, 100, -68, -21, 84, -38, 24, -89, 69, -108, 44, -126, -10, 68, -61, 38, 21, -13, 24, 67, 88, 49, 94, 112, -94, -97, -45, -21, -59, 66, 9, 121, -122, 19, -2, -9, 6, 107, -110, 127, -126, -83, 52, 111, 28, 4, -94, -69, -24, -96, 51, 54, 81, -39, 116, 38, -99, 51, -124, -19, -114, -125, -70, -51, -74, -105, 110, 76, 63, -102, -47, 37, 62, -55, -57, 73, 66, 59, -4, -64, -98, 6, -89, 19, -10, -117, -11, 124, -82, -59, 80, -45, -7, 124, -70, 49, 21, 45, -36, 38, 55, -94, -104, 54, 6, 31, 81, 118, 11, -100, -1, 83, -18, 66, -66, -26, 24, 53, -33, -104, -54, 35, 112, 95, 62, -102, 99, 84, -50, -37, 119, -68, -19, -55, 2, -125, -42, -118, 7, 55, 67, 59, -113, 64, 86, -66, 100, 51, -76, 101, 34, 9, 119, 55, -20, -61, 103, -80, -112, -27, -21, -7, -15, 104, -59, 116, 59, 124, 79, -122, -19, -29, 126, -118, -126, -29, 113, -37, 69, -34, -46, -28, -10, 72, 80, -112, 119, 60, 8, 43, 115, 44, -92, -19, 98, 72, -7, 94, 13, 60, 27, -30, -35, -118, -21, 3, 30, 113, 0, -83, 77, -52, 105, -71, -20, 127, 16, -6, -93, 94, 54, -127, 44, -66, 37, -109, -32, 69, -82, -71, -127, -85, 89, 4, 25, -128, -65, -47, -59, 10, 67, -99, 11, 64, -118, 45, 6, -50, -96, 67, 111, -36, -108, -67, 30, 27, 77, 54, 23, 27, 35, 49, -71, -64, 87, -109, -32, 91, -107, -94, 84, -47, 12, 61, 8, 17, -124, -41, 99, 34, -100, -69, -117, -76, -5, 89, 32, -25, -26, 56, -16, 30, -27, -3, 15, -127, -94, 8, -86, -85, -52, -42, -2, 11, 110, -66, -75, -96, -74, 26, -86, 59, -3, 68, -7, -26, 23, -44, -113, 113, -89, 90, 75, -8, -100, -50, -118, -35, -33, -124, -23, 116, 104, -96, 80, 103, -71, 26, 40, 80, -54, 24, -110, 116, 118, 10, -104, -48, 98, -107, 113, -70, 17, 6, 58, -103, 77, 46, -107, 120, -57, 112, -127, 51, 114, -110, -74, -58, -74, 112, 41, -91, 67, -80, -24, 61, -95, 51, 47, 111, 12, 62, 80, -62, -57, 1, -62, -110, 56, 61, -33, 14, -25, 112, -45, -42, 94, -108, 26, -9, 20, -102, -112, -17, -56, 71, -91, -109, -4, -123, 6, 58, 2, -60, 92, -5, 92, -106, 117, 93, -109, -64, -121, 19, 42, 124, 77, -87, 67, -53, 44, 9, 118, 38, 40, 97, 68, 16, 94, -40, 101, -61, 55, -61, -107, 30, -71, -61, 64, 11, -49, 63, -104, 94, 75, -4, -14, 79, 103, -123, 69, -5, 81, -19, -67, 92, 4, -95, -11, -124, -71, -24, -51, 114, -86, 102, 110, 68, 38, 83, 120, 116, 17, 93, 20, -67, 99, -115, -88, 52, 44, -122, 38, 35, 115, 94, 118, -110, -34, 108, -35, -52, -32, -5, -103, 58, 105, -14, -115 );
    signal scenario_output : scenario_type :=( -128, 127, 127, 127, -128, 127, 127, 127, 116, 127, 127, 39, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -42, -128, 127, -128, -128, -128, -128, 127, -128, -107, 127, 127, -128, 127, -34, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -106, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 12, -128, -44, 127, -128, 127, -128, 127, 127, 127, -34, 127, 127, -5, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -117, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 65, 127, 127, 106, 127, 127, -128, -128, -128, 17, -128, -128, -128, -128, 11, -122, 127, 127, 127, 127, -37, 127, 127, -128, 127, -57, 127, -78, 127, -128, 127, 47, -128, -128, -128, -128, -128, 127, -128, -128, -60, -128, 127, -128, 127, 127, 127, 90, -45, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -123, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -53, -111, 127, 127, 127, 127, 127, 127, 127, 49, 127, -36, 127, -128, 60, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 102, 127, 127, -6, -128, 127, -128, -128, -32, 127, -128, -27, 127, 127, -10, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -106, 127, 127, 127, 127, 127, 127, 127, -90, 127, -128, -36, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -109, -128, 127, -18, -12, -128, -128, -128, -128, -128, -128, 127, -76, 118, -128, -128, -128, 127, 127, 127, 127, 127, -22, -85, 52, 127, -128, 127, -128, -128, 127, 127, -33, 127, 96, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 44, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -107, -128, -128, -128, -128, -128, -128, 127, -128, -128, -31, -128, 127, -50, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -100, 127, 127, 127, 127, 127, 127, 127, 127, -128, -42, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -43, 127, -128, -128, -80, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -117, 127, -128, -128, 107, -128, -36, 127, 127, 127, 127, 127, 127, 86, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 27, -128, -128, 127, -1, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 18, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -43, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -92, -128, -128, 75, -7, -128, 102, 69, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -81, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 111, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 85, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -114, -128, -103, 127, 127, -128, -128, -112, 127, -128, 21, 127, 127, 127, 127, 127, 88, 127, 127, 87, 127, 127, 127, -39, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -102, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -81, 127, 127, 127, 127, 127, 127, 127, 65, 48, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 121, -128, 127, 127, 127, 127, 127, 98, 127, -128, 127, -128, -128, 127, 65, -128, -128, 127, -78, -128, 127, -53, 127, -128, 108, -128, -128, -48, -128, 127, 127, -128, -128, 102, 127, -128, 0, 127, 127, -109, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -26, -128, 47, -128, -128, -128, 127, -128, -74, -73, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 85, -128, 127, 127, 127, 127, 127, 127, 127, 39, -49, -128, 127, 127, -128, 127, 127, 127, 127, 123, 127, -128, -68, -128, 97, 127, -58, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 44, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 100, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 34, 127, -36, 74, 13, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 3, -128, 127, 75, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -68, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -47, -128, -128, -128, -128, -128, -128, -128, -128, 109, 127, 127, 127, 127, 127, 127, 5, -128, 127, -128, -128, -128, 127, -128, 127, 127, -93, -128, 127, -128, -87, -128, -128, -128, -128, -128, -128, 127, -128, -128, -81, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -48, -128, -128, -128, 127, -128, -128, -128, 49, -1, -128, -3, 127, -128, -128, -128, 127, 127, 127, 127, 87, -128, -128, -128, 15, 127, 127, 127, 127, 127, -13, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 96, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 112, 127, 127, -128, -128, 127, 127, -128, -128, 68, -128, -128, -128, -128, -121, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -114, -128, -128, -128, 127, -128, -128, 127, -128, -128, 38, 127, -128, 127, 127, 127, -128, 22, -128, 127, -128, -128, -128, -112, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -13, 127, -113, 127, 113, -128, -60, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -50, 127, -128, 113, -128, -128, -128, 28, -128, -128, 49, 127, -128, -128, 127, 127, -24, 127, 66, 127, -128, 106, -128, 127, -128, 29, -128, -128, -128, -128, -128, -128, 127, 29, -128, 127, 127, 127, -128, -128, -128, 127, -18, 127, 127, 127, 127, 127, 127, 10, 127, -123, 127, -128, 127, 15, 127, -128, -128, -128, 43, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 5, 127, -128, -128, -128, 127, -91, -128, -128, 127, 127, 23, 127, 127, 23, 127, 117, 69, 127, 127, -128, 26, 127, 102, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -71, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -90, -128, -128, -128, -128, -38, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 102, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, 106, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -106, -128, 127, -128, 127, -128, 127, -128, 127, 111, 127, 127, 127, 127, 127, 127, 127, 127, 127, 58, -48, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -80, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -106, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 47, 127, 127, 127, -128, 76, -128, -128, -128, 39, -128, 127, 80, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 22, 127, -32, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -24, 109, -128, 127, -128, 28, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 100, 127, -128, -86, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -81, 127, 127, -128, 127, 127, 127, -119, 127, -128, -128, 127, -128, -128, 112, 127, 81, 21, 127, 55, -128, -128, 127, -128, -128, -128, -59, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 87, 127, -128, 127, 127, 23, -100, 127, -128, -128, -128, -128, -128, -128, -128, 127, 50, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -52, -128, -128, 127, -128, 12, 127, 127, 113, 127, 127, 127, 127, 127, -128, -128, 24, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 92, -128, -128, -128, -128, -128, -128, -16, -128, -128, -128, -128, 127, -128, 127, -109, 127, -128, -66, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -96, -128, 49, -128, 2, 75, 127, -128, 127, 127, 127, 127, 127, 127, -80, 127, 79, -128, -128, -128, 127, 127, -18, 127, 127, 127, -128, 127, 71, 127, -128, -128, -128, 93, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 10, 127, 127, -32, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -107, -128, 76, -50, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -39, -128, 127, -128, -128, 127, 127, 127, 6, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 95, 127, -128, -128, 127, 127, 127, -103, 127, -128, -128, -128, -128, -26, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -59, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 88, -128, -128, -128, -128, -128, -128, -128, -128, -128, 91, 127, 127, -128, -128, 127, 127, 127, -128, 127, 71, 10, -128, -85, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -93, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 97, -128, 127, -96, 127, -128, 127, -128, -128, -128, -102, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -97, 127, -76, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -102, 127, 127, 127, 127, 127, 127, 127, 127, 127, -111, 70, 100, 127, -71, 127, 127, 127, 127, -102, -128, -128, -128, 15, -128, 127, -93, 127, -128, 127, -111, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -52, 127, -128, 127, -128, -81, -128, -128, -128, -128, 127, -78, 127, 127, 127, -128, -128, -128, -2, -128, -128, -34, -128, -128, -128, 127, -128, -128, 34, -128, -128, -128, 97, -128, -128, 127, 127, 127, -128, 127, 24, 127, -128, 127, 127, 127, -128, -128, -59, -128, -128, -128, -128, -128, 118, -128, -128, -128, 71, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 16, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 95, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -6, 127, 38, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -85, -128, -128, -54, 127, 127, 127, 127, 127, 18, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -98, -128, 127, 127, 127, 32, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -75, -71, 127, 54, -128, -128, 127, -128, -128, -128, 88, -47, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -37, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 106, -128, -128, -128, -128, -26, 127, 127, 127, 127, -49, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 26, 127, -128, 127, 127, 127, -128, 7, -128, -128, -128, -26, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 37, -128, 127, 127, 127, 127, 127, -128, -128, 22, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 109, -128, -128, -128, -128, -128, -3, 127, 127, 127, 127, 127, 127, 127, 127, 3, 127, -28, -128, -128, 127, -128, 127, -128, 127, 127, 127, -75, 58, 127, -128, -128, 63, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -91, 127, -128, -128, -128, 127, -128, 88, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -73, 127, -128, 127, -128, -128, 127, 45, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 7, -128, -128, -128, -128, -128, -128, -128, -128, 13, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 36, 113, 127, -128, -128, -128, 127, 113, -128, 127, 127, 79, -128, 127, 127, -128, -128, -128, 127, -128, -90, -128, 95, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -6, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -75, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -69, -127, 127, 21, 127, 127, 47, -128, 127, -128, -128, -128, 127, -128, 127, -128, 34, 127, 44, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -18, 127, 127, 127, 127, 127, 127, 127, 24, -128, -128, -128, -31, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -86, 127, 127, -128, 127, 127, -116, -128, -128, -12, -128, -128, 76, -128, -128, -128, -49, -128, -128, 127, 127, 127, 127, -128, -128, -123, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 81, -128, -128, -128, -128, -128, -128, -128, -128, -128, -31, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 122, -128, 127, 17, 127, 127, 29, -128, -128, -128, -128, -128, -128, -128, -128, -128, -100, -128, -128, -128, 127, 36, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 38, -128, 127, -127, -128, -128, -128, -29, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 7, -128, 127, -128, -91, -50, -128, 127, -128, 127, -128, 127, 6, 127, -128, 127, -128, -128, -128, -68, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 116, -128, 127, 127, 127, 127, -23, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -95, 127, 127, 127, 127, -128, -128, -128, 127, 127, 81, 127, -128, -106, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 39, -128, -128, -36, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -26, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -47, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 87, 127, 127, 127, 127, -128, -128, -128, 127, 79, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 10, -38, 6, 127, 127, -124, 127, 127, -22, 80, -66, -128, -128, -128, 127, -128, -128, -128, 127, -119, -128, -128, 5, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -87, 127, -128, -128, -128, -128, -128, -128, -128, -128, 21, -128, 127, -128, 127, 54, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -78, 93, -128, 127, -128, -128, -128, -128, -128, 111, 127, -128, 127, 116, -91, -128, -128, -128, -128, -128, 127, -128, -128, -103, -128, -128, -128, 127, 66, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -8, 127, -128, 127, -128, -128, -128, 127, -128, 33, -128, 127, -128, -128, -114, 127, 57, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -123, 127, -128, 127, -128, 127, 127, 127, -128, -128, -22, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 26, 127, 127, -49, 127, -128, -128, -128, 64, -128, -128, -128, -128, -128, -128, 127, -128, 27, 127, 127, 127, 127, 127, 78, 57, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 33, 127, -1, 127, 127, 127, 127, 121, -128, -128, -31, -128, -55, 127, -128, -128, 127, 127, -128, 38, -128, 127, -128, -128, -128, 127, -128, -128, -58, 127, 60, -128, 127, -128, 127, -128, 127, -128, -121, -128, -128, -27, -128, 127, -128, -128, 127, -7, 98, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 43, -59, 127, 127, -128, 127, 127, -128, -31, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -31, 127, 127, 127, 127, 127, -128, -128, -106, -58, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 124, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 100, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -21, 74, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 101, 127, 127, 8, 127, 127, 127, 24, 127, -122, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 5, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -29, 127, -128, 100, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 85, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 107, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -60, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 123, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 11, -128, -128, -128, -128, 10, -128, -23, 85, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -10, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 93, 127, 127, -128, -128, 39, 58, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -33, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -101, -128, -128, -128, -128, -128, -90, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -3, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 6, -128, -128, -128, -128, -128, 127, -128, -78, -128, 127, -128, -5, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 52, -128, -128, -128, -128, -128, 127, -118, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -101, -128, 76, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 8, -128, 66, 127, 127, 52, 127, 127, 127, 127, -111, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -5, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -122, -45, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 53, 127, 127, 127, 101, 127, 127, 127, -128, 127, 107, 127, -128, -128, 24, 127, 127, -128, 127, -128, 127, 127, 127, 49, -70, -128, 34, -128, -10, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 90, 127, 127, 127, 127, 127, 11, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 69, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -24, 127, -128, -128, 0, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -92, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 124, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 111, 127, 127, 127, 127, 127, -5, -15, 69, 127, -128, 11, 127, 127, -128, -128, 127, 127, -128, 0, 127, -128, -128, 127, -11, -128, -23, 127, 127, 127, 127, 127, 48, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 42, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -49, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 42, -88, 109, -128, 127, -55, 127, -49, 127, 127, 127, -128, 127, 127, -101, -128, 127, -101, -79, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -65, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -80, -128, -128, 127, 127, 127, 127, -128, 127, 127, -66, -128, -128, 127, 127, -109, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -91, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 45, 127, -128, -128, -128, -54, 127, 76, -86, 127, 127, 127, 127, 127, 127, -128, 127, 44, -128, -128, 127, 44, 127, -128, -44, 127, -128, -128, 29, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -33, 127, -128, 113, -128, -128, -128, -128, -128, -128, 127, -128, 127, 95, 127, -128, -42, -128, -128, -128, -128, 127, 91, -7, 127, 127, 127, -128, -6, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -108, 127, 127, -128, 127, -128, 127, 34, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 33, 80, 127, 93, -118, 91, -128, -57, 127, -6, 127, 127, 127, 127, 127, -128, 114, -128, -128, -128, -128, -128, -128, 70, -128, -128, 127, -128, -128, -128, 127, -128, -112, -128, -128, -128, -128, -128, -128, 8, 127, 127, 127, 127, -128, 108, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -17, -128, 100, -18, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -21, -128, -128, 127, -128, -128, -128, -128, -128, -128, 16, 127, 127, 127, 1, 13, -128, 127, -128, -128, -32, -95, 34, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 78, -128, 127, -128, 127, -128, 97, -128, 127, 127, -128, 127, -28, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -7, -128, -128, -111, 127, 127, 127, 127, 127, -128, -128, -128, 57, -128, 32, -75, 127, 127, 127, 127, -108, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -85, -128, 127, 127, -128, -11, 71, 127, -128, 127, 127, -128, -128, -128, 43, -128, 127, -128, -128, -128, 127, -128, 127, 127, -90, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 63, -128, -128, 18, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -74, 127, 127, -128, 127, 127, -128, 127, 127, 127, 27, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 116, -128, 127, -128, -81, -128, -65, -128, 127, -128, 114, -128, 127, -128, -128, -128, 127, 127, 127, 0, 127, 127, 127, -33, 127, 6, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -75, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -91, 127, -128, 11, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -18, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -73, 127, 127, -128, 127, 127, -128, -128, -128, 58, -128, -128, -128, -128, -128, -128, 114, -128, 127, 127, -128, -128, 127, -128, 53, 100, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -86, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 28, -8, 127, 127, -128, -128, -128, -128, -128, -128, 69, -70, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -36, -34, -128, -128, 127, -128, -43, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 2, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 85, -128, -128, -128, -128, -128, -128, -128, -128, -114, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -15, 86, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 48, 127, -128, 127, -128, 127, -128, -128, -45, 127, -128, -128, -128, -128, -128, -128, -128, 127, -60, -128, -128, 127, -128, -128, 93, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, 71, 127, 127, -128, 127, 127, 127, 24, 127, 127, -128, 127, 127, -50, -128, 127, 70, 127, -128, 127, 127, 127, -3, 127, -128, 127, -100, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -101, -128, 127, -97, -50, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -12, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -73, -128, -128, -128, -128, -128, -128, 18, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 1, 127, -128, -128, 127, -128, -128, -79, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 18, 127, 127, 127, 127, 127, 127, 102, -128, 127, -128, -128, -128, 71, -128, -128, 18, -128, 127, -96, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 32, -16, 127, -128, 127, -128, 127, 42, 127, -128, -128, 127, -128, -128, -7, 127, -128, 127, 127, 44, -128, 127, 127, 127, 12, 127, -128, -128, -128, 127, 75, 50, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -101, 127, -128, -128, -128, -128, -128, -128, -128, -28, -128, -128, 127, 127, 127, 127, 127, 127, 127, 29, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 57, 127, 127, -128, -128, -128, -128, -128, -128, -128, 1, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -27, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 114, -103, 127, 127, -74, 127, 127, -128, -128, 127, -128, 34, 127, 127, -128, -128, 63, -128, -128, 102, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -18, -128, 127, 127, 127, 76, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -44, 123, -128, 127, -128, 127, -128, 127, -128, 111, -128, -128, -128, -128, -112, 127, 127, 127, 127, 127, 127, 127, -13, -128, 127, 127, -111, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -7, -128, 127, -128, -128, -128, 127, 11, 127, 127, 127, 127, 127, 10, 127, 127, 127, 127, 127, -128, 127, 127, 127, -5, 127, -128, 0, -128, -114, -128, -128, 127, 127, 127, 127, 75, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -47, -49, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 2, 127, 127, -128, -128, 31, 23, -128, -57, 38, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -52, -128, -128, 127, 76, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 85, 7, 90, -128, -128, -128, -128, -128, -112, 127, 97, 80, 90, 127, 127, 127, 127, 127, 127, -128, 127, 127, -64, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -123, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -78, -102, -128, -128, -128, 127, -128, 127, 27, -128, -128, 127, -128, -128, -86, 127, 127, 127, 127, 127, 127, 108, 114, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -34, 127, 127, -128, -128, -127, -128, 127, -128, -128, -128, 127, -128, -128, 100, -42, -128, 0, -128, 111, -128, 127, -128, 127, -128, 127, 74, 127, 127, 127, 127, 127, 127, -128, 39, -128, -128, -128, -106, -128, -128, -128, 127, 127, 127, -128, -50, 127, -128, -128, 127, 127, -128, 127, -8, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -97, -128, -102, 127, 127, 127, 127, 127, 127, 127, -128, 127, -22, 127, -128, 127, -128, -128, -128, -118, -128, -128, -128, -128, -128, -128, -128, 127, -27, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, 12, 121, -128, 17, 127, -128, -29, 127, 98, -70, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 5, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -6, -48, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -12, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 108, 127, 127, 127, 127, 127, -59, 127, -128, 127, -128, -87, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -18, 127, -122, -128, -128, -128, -128, -128, 127, -128, -128, -70, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -16, -13, -128, -128, -128, -128, -128, 127, -128, 127, 36, 127, -93, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -64, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, -95, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 69, -128, -128, -128, 16, -128, -128, 127, 127, 127, 127, 106, 127, 127, 127, -52, 127, 127, 127, 127, -128, -128, -128, -128, -128, -100, 127, 127, 127, 127, 127, 92, 32, -128, 127, -128, -118, 127, 127, -23, 64, 107, 127, -128, -128, -128, -128, -111, -128, 127, -128, 34, -128, 29, -128, -128, 127, -17, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -1, -128, -24, 79, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 64, 127, 127, 127, -6, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -68, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -60, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 68, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 116, -128, 127, -128, -109, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 33, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -117, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -122, -128, 127, -106, -128, -128, -128, 127, 127, 127, 91, 127, 127, 127, -128, -128, -128, 127, -128, -128, 33, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -15, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 123, -128, -128, -123, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -111, 97, -128, -128, -128, 127, -128, 86, -128, -128, -128, -128, -128, -128, -128, 127, 112, 32, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 18, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 108, 127, -124, 127, 127, 127, -128, 127, -128, -128, -119, 119, -128, -128, 127, 127, 127, 127, 127, 127, 57, 127, 127, 127, 127, 127, 127, 127, 127, -24, -128, 27, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -7, 55, 127, 127, -96, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 22, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 58, -128, 42, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 10, -128, 127, 45, -128, -128, 127, -128, -2, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -90, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 48, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -81, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -66, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -53, -128, -128, -15, -128, -128, 119, 127, 127, 127, 127, 127, 127, 70, 127, 127, -106, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -117, 127, -76, 127, -128, 64, -128, 92, 38, -128, 127, 127, 127, -128, 127, 127, -66, 127, 127, 119, 81, 121, -70, -128, -128, -128, -128, -128, -128, -128, -128, 10, 127, 127, 127, 127, 127, 127, -34, 127, -128, -128, -128, 98, -128, 127, -128, -128, 127, 127, -128, -128, 75, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -95, -128, 127, -128, -86, 127, 127, -128, 127, 127, 127, -128, 127, 123, -128, 97, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 21, -128, 127, -128, -78, -47, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 11, -37, 45, -128, -128, -128, 44, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 6, 127, -128, -128, 127, -128, 68, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -73, 127, -128, 127, 127, 127, -6, 127, 127, 127, 127, -59, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -116, -128, 37, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -58, -128, 127, -128, 127, -128, 127, -45, -128, -128, -128, 123, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 87, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 36, -68, -128, 127, 127, -21, -128, 127, 127, -128, -128, -128, 127, -128, 80, 127, 127, -128, 127, -109, -128, 127, -128, -3, -128, 127, -128, -1, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 108, 127, -59, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 102, 127, -128, 76, -128, -128, 127, -128, -128, 21, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -39, 127, 127, 127, 127, 127, 127, 127, 127, 109, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -106, -112, -128, -128, 127, -128, 127, -128, 127, -128, 53, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -102, 121, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 64, 127, 127, -128, -128, 127, -128, 59, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 57, -128, -128, -128, -128, -24, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, 48, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 112, -128, -128, -128, 68, 127, 127, -93, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -60, 127, 127, -2, 127, -128, -128, -128, -128, -128, 127, 13, 127, -128, 127, -128, -128, -128, -128, -128, -114, 127, 127, 127, 127, 127, -128, -128, 102, 127, -128, 127, 127, 127, 127, 127, 85, -128, 127, 117, 127, 127, 127, 127, 127, 127, 127, 127, 127, -97, -128, -128, -128, -128, -66, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -1, -128, -128, -128, -128, 113, -128, 127, -128, 127, -73, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 124, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 111, -128, 5, -128, 127, -128, 13, 79, 127, 127, -128, 42, -128, -44, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 106, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 102, 85, -128, 127, -128, -75, 127, -128, 127, 81, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 118, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -16, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -98, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 24, 127, -128, -128, -128, -128, -128, -128, -128, -128, -1, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 32, 49, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 118, 127, -128, 127, -102, 127, 127, 127, -128, 127, -128, 111, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -47, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, -33, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -91, -128, 127, -128, -128, -128, 17, -128, -128, 127, 58, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 122, -128, -128, -128, 127, -128, -128, -128, 75, -128, -128, -128, -128, -34, -128, 97, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 97, -50, 127, -128, 127, -128, 127, -128, -128, -128, 127, 3, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -38, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -42, 127, 127, 127, 127, -128, -128, -128, -28, 127, -128, 127, 127, 127, -128, 127, -128, 127, -112, 127, 74, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 39, -128, -109, -128, 127, -128, 127, -128, 127, 127, 127, -54, -128, 127, 127, 127, -128, 127, -114, 127, -128, 127, -128, 127, -128, 0, -128, 127, -128, -128, -128, -128, -128, -128, -88, -128, -128, 127, 127, -128, 127, -53, -128, -128, -128, -128, -128, -128, -128, -128, 65, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -7, -128, -128, -128, -128, -128, -128, -128, -6, -128, -117, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -86, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 74, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, -42, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -57, 127, -128, 97, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -76, 127, -128, -128, 127, 127, -128, -11, -128, 127, -102, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 37, 0, -128, -128, 127, -47, 127, -128, 127, -79, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 33, 127, 127, 108, -128, 127, -128, 113, -128, 127, -128, 74, -128, 127, -128, -128, -86, 127, 127, -17, -88, 127, 65, 127, -128, -128, 127, 127, 127, -118, 127, -128, 127, 31, 117, 127, 127, -128, 127, -128, -128, -128, 127, 39, 75, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 111, -128, -128, -44, -128, -128, -128, 127, 127, 127, 127, 127, 123, 127, 127, -47, 64, 127, 127, 127, -128, 75, -128, -128, -128, -128, -128, -128, -128, -128, 127, -109, 111, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -87, -128, -128, -128, -118, -128, -128, -128, -128, -3, 127, 127, -66, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -39, -128, -128, 127, -128, -128, -128, -128, 28, -128, 65, -128, 127, -128, -128, -128, 127, 127, 127, 42, 127, 127, 127, 127, -128, 127, 127, 127, 127, -53, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 63, -128, -80, 113, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 93, -128, 127, 127, 127, 127, 127, 127, 127, 102, 127, -128, -3, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 97, -128, -128, 60, 127, -128, 127, 127, 127, 127, 127, 127, 58, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 8, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -101, -91, -59, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 15, 127, -128, 22, -128, -128, -128, 127, 127, -122, 127, 127, 127, 123, 127, 127, 127, 127, -12, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 74, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -12, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -47, -128, 127, -128, -128, -128, -128, -117, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 43, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 8, 31, 127, 127, 127, 127, 127, -128, 127, 127, 127, 64, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 43, -128, 127, -128, 127, 127, 127, 8, -128, -39, 53, 127, 127, 127, 127, 127, 127, -128, -128, -128, -103, -128, 127, -128, 127, 127, 127, -95, 127, -128, 127, 127, 127, -128, 114, 127, 119, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 86, -37, 127, 127, -102, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -31, 64, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -97, -57, 127, 127, -28, 127, 69, 127, -128, -22, 127, 57, -22, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 103, -96, -74, -128, 127, 127, 127, -128, 127, 127, 127, -97, 127, -128, 57, 127, 127, 0, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -48, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -48, -11, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -23, -128, -128, -128, -128, -128, 127, 127, 127, -128, 2, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 32, -128, 127, 127, 127, -128, 113, 127, 127, 27, 127, 127, 127, 127, 127, 127, 12, -128, 127, 127, 88, 127, 127, 127, -101, 127, -128, -128, -128, 127, -128, 16, -128, 127, -128, 127, 127, 127, -3, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -7, 127, 127, 127, 127, 127, 127, 127, 127, -17, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -38, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -12, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 2, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 6, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -107, -128, -128, -128, 127, -128, 127, -128, -128, 2, -128, -128, -128, 113, -106, -128, 127, 127, 127, 127, 106, -128, 48, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -1, -128, 39, -128, -128, -128, -76, 127, 0, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 102, -128, -128, 127, 12, -128, 112, -128, -128, -128, -114, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 6, -128, -128, 127, 127, -128, 114, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 88, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -15, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -47, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 124, 127, 127, 127, 127, 127, 127, 127, 127, -37, -128, 127, 127, 127, 22, 127, -128, -122, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 44, 76, 101, -128, -128, -128, -128, -128, -128, -128, -38, -128, -128, 59, 127, -128, -128, 127, -128, -128, 96, 127, 127, 127, 127, 21, 127, 127, 127, 127, 127, -128, 87, 127, 0, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -73, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -47, -128, 127, 127, 127, 127, -112, -128, -128, 86, 55, -6, 127, 127, 127, 127, 127, 127, 127, 127, -98, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 13, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -10, 127, -74, -128, 127, 127, -90, 127, 66, 127, -128, 127, -128, -81, -128, 127, -123, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -79, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -93, -128, -3, 127, -128, -128, 127, 127, 127, 53, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -121, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 71, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 52, 127, 127, -128, -128, 127, 127, -128, -128, 80, 127, -128, -128, 127, 127, -128, 127, -128, 47, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 109, 127, -128, -128, 122, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 11, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 64, 10, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -8, 127, -109, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -63, 127, -128, 127, -128, -3, 127, -128, -69, 127, 127, -18, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 75, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -1, -108, -128, -15, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 75, -128, -44, 127, 127, -128, -128, -128, 127, -128, -59, -128, -128, -128, -12, -128, -128, -128, -128, 127, 127, 127, -122, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -86, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 87, -128, -128, -128, -128, 97, 75, -128, -128, -13, -128, -128, -128, 127, -128, -128, 100, 127, 38, 127, 127, 31, -97, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -44, -128, -128, 127, -128, -128, -128, 123, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 85, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -116, 127, 127, 60, 127, 127, 127, 127, 127, 127, 86, -128, -128, -128, 127, -128, -128, -128, -39, -128, -128, -81, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -85, 127, -128, 127, 127, 127, -128, -1, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 5, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 75, 127, 127, 127, 127, 127, 127, 103, 127, 15, -128, 127, 48, 127, 127, 127, -128, -128, -128, -128, -44, 127, 108, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, 66, -128, 127, -128, 127, -12, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -87, -128, -128, -128, -128, -128, -128, -101, -128, -128, -128, 127, -128, 127, 111, 127, 127, 127, 127, -113, 127, -128, -128, -128, 127, -128, -128, -128, -96, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 122, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 45, -103, -128, -128, 127, -128, 127, 70, 127, 127, 127, 127, 127, 127, 127, -128, 64, -128, -8, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -119, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -124, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 80, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -39, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 0, 86, -128, -128, 106, -102, -128, -128, -65, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -111, -128, -128, -128, 34, -128, -128, 127, 127, -128, 127, -36, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 44, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 3, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -13, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -27, 127, 127, -42, 127, 127, -128, -128, 65, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -124, 127, 127, 127, -128, 21, 127, 127, 127, 127, 127, 127, 127, 44, -128, 127, 127, 121, 127, 127, 0, -128, -128, -128, -128, -128, -128, 44, 127, 127, -128, 127, 33, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 69, -85, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -18, 127, -128, 127, 127, 127, 127, 127, 127, 65, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -18, -128, 127, 127, 127, 55, -91, -128, -128, 127, -128, -128, 127, 127, -128, 6, 127, -128, -128, 127, -128, -128, -128, 127, 127, 49, 127, 127, 127, 127, -128, 12, 127, -128, -123, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 107, -114, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 97, -128, 127, -128, 127, -128, -128, 127, -128, -91, 103, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -59, 127, 127, 127, 127, 127, 127, -34, -128, 127, 127, -128, -128, 127, -17, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -114, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 70, -128, -128, 127, -128, 127, -37, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 68, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -12, -128, 127, -128, -128, -128, -16, -128, -106, 127, -100, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -7, -128, -128, 127, -128, 127, -128, 127, -97, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -121, -128, -128, 127, -128, 127, -128, 127, 127, 107, -32, -128, 103, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -37, 127, 85, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -17, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 81, -128, 127, 127, 127, -128, -128, -128, -2, -128, -128, 127, 127, 127, 127, 127, 127, 36, -128, -47, -128, -128, -128, 127, 70, 0, 127, 127, 127, -128, 26, -128, -128, -128, -31, -128, 24, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 18, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -80, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 79, 127, -128, -128, 127, 111, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 106, 127, 66, 127, 127, -128, 127, -97, 127, -128, -98, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -87, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -85, 127, 127, -128, 79, 127, -128, -128, 127, -128, 127, 18, 127, -64, 127, -66, 127, 1, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -81, 127, 127, -128, 127, 127, -128, 127, -107, 90, -128, 75, -128, 127, -128, 127, -128, -7, 10, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 124, 127, -128, -121, 127, -128, -128, -128, -17, 127, 52, 127, -128, -128, 127, -128, 65, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 76, -128, 127, -128, 127, -49, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -63, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -74, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -53, 127, 81, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 90, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -12, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 58, 127, 127, 127, -128, -128, 127, 127, -128, -128, -7, 96, 127, 127, -128, -128, -128, 127, -128, -109, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 3, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -32, -128, -128, -128, -95, -128, -128, 127, 127, 33, 127, 127, 127, 127, 127, -128, 127, 127, 127, -39, 127, -128, -128, -128, 109, -21, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 98, 127, 119, 127, 127, 127, -128, -128, -128, -128, -119, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -119, 127, -128, 118, -128, 127, 127, 127, 127, 76, -128, -128, 127, -88, 78, 127, -6, 127, 127, -80, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 3, 127, -128, -128, 0, -128, -128, -128, -54, -128, -128, -128, 127, -90, -8, -128, 127, -128, -128, 127, -7, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 27, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -43, -128, -128, -128, -128, -128, -128, -128, -6, 127, 127, 127, 6, 127, 127, 127, -128, 76, 127, -128, 127, -128, -128, 127, 78, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -101, 127, 127, -128, 127, 127, 127, -128, 127, 127, -108, 27, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -86, -18, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 1, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -80, -128, -128, -128, 127, -96, -128, 127, 127, -128, 6, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 106, -128, 127, 127, -128, 127, -32, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -106, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -47, 122, 127, 127, -128, -128, -53, -128, -128, -128, 63, -128, -128, -128, -27, -128, -128, -128, 34, -128, -128, -128, 127, 1, -128, -128, 42, -128, -128, 81, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -107, 127, 127, 127, 127, 127, 127, -122, -128, -68, 86, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 106, 127, 127, 127, 127, 127, 127, 127, 127, 127, -70, 127, 127, 127, 127, 127, 127, -118, 127, -128, 127, -128, -128, -128, 127, 45, -128, -128, -128, -128, 7, -128, -128, -128, 34, 17, -128, -128, -128, -128, -128, -6, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 37, -128, 74, 127, -38, -122, 127, 127, 127, -128, 98, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, 57, -128, -128, -128, -128, 127, -128, -128, -54, 127, 127, 127, 127, 127, 127, 127, -128, 127, -122, 127, -128, -15, -128, 127, -124, 127, -128, -128, 127, 127, 66, 127, 127, 127, -128, 127, -102, -128, 11, 112, -128, 127, -128, -128, 127, 127, -29, 92, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -28, -128, 127, 127, 127, -128, 95, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 118, -128, -128, -128, 127, 86, -128, -128, 127, 11, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -6, -128, -128, 127, 116, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -33, -128, -54, 79, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -111, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 73, 127, 63, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 21, 127, 127, -86, -76, -128, -128, -128, -95, 127, 52, -128, 127, 127, -128, 127, 127, -128, -128, 116, -128, -128, -128, -128, -128, -128, -128, -128, -122, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -93, -128, -128, -128, -95, 123, 127, 127, 127, 127, 127, 127, -12, 127, -128, -128, -128, -55, -128, -128, 127, 127, 127, -119, 127, -128, -128, -128, -128, -52, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -49, 127, 3, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 47, 39, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -103, 127, 127, 127, 43, -128, -128, -23, -128, -128, 127, -128, -128, 127, 127, -128, 86, 127, -128, 127, 127, -3, 127, 8, -128, -128, 36, -128, -128, 21, -11, -128, -34, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -2, -128, -128, -128, -128, -128, -128, 93, -128, -128, 127, 127, 127, 127, -128, -102, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 100, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -86, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -49, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 63, -22, -128, -128, -128, -128, -128, -128, -128, -18, -128, -128, 127, 127, -47, 127, 127, 127, 27, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 73, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 98, -128, 127, -128, -128, -128, -111, -87, 127, -128, 113, -128, -128, -128, -128, 127, 127, -128, -118, 127, -128, -128, -128, 49, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -11, 127, 127, 93, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -98, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 54, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 114, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 26, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, 7, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 109, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -39, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -31, 127, -75, 127, 127, -79, -128, -128, -29, -128, -128, 127, -128, -128, -128, -121, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -1, -128, -128, -128, -128, -128, -128, 36, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -102, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -12, 121, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 66, -59, 127, 127, 127, 90, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 122, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 107, -128, -128, -128, -128, -128, -128, 127, 127, -128, 39, 127, 127, 127, 127, 127, -78, -128, 127, -128, 127, -128, 127, 127, 127, -68, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -11, 127, 127, -128, -128, 127, 127, -128, -128, 97, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 64, -128, 127, -128, -128, -12, 127, -128, -80, 31, 118, -128, 127, 33, -128, -128, 127, 127, 127, 127, 127, 101, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 55, 127, -128, 127, 127, 113, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 58, 127, 127, 49, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 3, 70, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 66, -128, 127, -128, -128, -128, 127, 71, -128, 127, 127, -128, -128, 127, -71, -128, -102, 127, -128, 66, 127, -128, 127, 127, -128, -128, 127, 127, 103, 127, 127, -128, -128, 127, -128, 7, 113, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -65, -128, 127, -128, 127, 127, 127, 29, -37, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 2, 127, -128, -128, -128, -128, 68, 127, 112, 92, 1, 0, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 85, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -106, 127, 127, -128, 127, -128, -128, -128, 127, -87, 127, -3, 127, 127, 121, -128, -128, 127, -128, 127, 1, 127, -128, 127, -15, -128, -128, -128, -128, -128, 127, -128, 3, 127, 127, -128, -128, -128, -128, -128, -128, 63, 43, -109, 127, 127, 127, -44, -118, 127, -95, 127, 127, 127, -69, 127, -114, -128, 127, -128, -128, 113, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 6, -128, 127, 127, 127, 127, 127, -128, -128, 78, -128, -128, 127, 127, -75, 127, 127, 127, -69, 127, 127, 127, -128, 127, -80, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -85, -128, 127, -73, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -16, 127, -128, -128, 127, -128, 63, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 52, 127, 127, -128, 127, 127, 127, 127, -1, 127, 92, -128, 22, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -17, 127, -128, 65, 127, -128, 10, 127, -128, -128, 127, 111, -128, -128, 127, 127, -122, -128, 113, 127, -128, 127, 32, -128, -128, -128, -128, -128, -128, -128, -128, -128, 31, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 27, 127, 127, 127, 127, -128, -128, 127, -17, -128, -128, 127, 127, 127, -128, 127, -128, 97, -128, -128, -128, 127, -128, -128, -128, -109, -128, -128, -128, -128, -128, 127, -128, -128, 2, -38, -128, -128, -128, 93, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -21, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 6, -128, 127, -128, -128, -128, 63, -128, 127, -63, -11, 127, 127, -128, -128, 81, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 15, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 65, 127, 127, 127, 127, 127, -128, -128, -79, 127, -128, -128, 127, -98, -128, 127, 127, -128, -37, 127, 127, 127, -128, 127, -128, -11, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -117, 127, 127, -128, -128, -128, 127, -128, -128, -128, 16, -65, 127, -128, -13, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -44, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 23, -128, -37, 127, 127, -128, 127, 127, 127, -96, -128, 127, -128, 54, -128, 127, -128, 127, 31, 127, -128, -128, -32, -123, -45, -98, 127, 127, 127, 127, 127, 63, -128, 127, -128, 127, -87, -2, -128, 127, 127, -128, -128, 1, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -70, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -64, 24, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, 92, 127, 127, -128, 76, 127, 18, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 64, -107, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -65, 18, 127, 127, -128, -128, 92, -128, -128, -128, 127, -128, -128, 127, -128, 53, -128, 127, -128, 127, 101, 127, 127, -128, -18, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 26, -26, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -22, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -113, 127, 127, 39, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 91, -128, 127, -128, -128, -128, -128, -128, -128, -100, -128, -128, 107, -128, 127, -128, -128, -128, 113, -128, -128, 127, -98, 127, 127, 127, 24, -128, -128, -128, -128, -128, -128, 101, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 91, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 10, 127, 127, 33, 127, 127, -128, 127, -128, -128, -128, 122, -128, -128, 127, -66, 127, -21, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 116, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -57, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -2, -128, 127, -128, 127, -128, 127, -128, -128, -128, -90, -43, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -36, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 34, 127, 127, 127, 127, 127, 127, 127, 127, 17, 127, 127, 127, -128, 127, 2, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 66, -128, 127, -128, -59, -128, 127, -128, -52, -128, -100, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -53, -128, -128, 127, -128, -128, -128, -22, -128, -128, -128, -128, -128, -128, 13, -53, 127, 127, 127, -128, -85, -128, -128, -128, -128, 127, -21, -88, -68, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 111, 11, -128, -128, 124, -128, -128, -128, 127, -31, -16, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -65, 127, -128, -128, -11, -128, 127, 127, 127, -128, 127, 114, -128, -47, -128, -60, -128, 52, 127, -128, 127, 54, 127, 63, 13, -128, 21, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -90, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -32, 127, 127, -128, 127, -128, 127, 17, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -121, 127, 127, 127, 127, 127, 127, 127, -128, 127, 24, 44, 127, 127, 127, 127, 127, 127, 127, 127, 3, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 119, -128, -128, -128, -128, -128, 127, -95, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 59, 42, -55, 127, 127, 127, 127, -128, -12, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 42, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 52, 127, 127, -81, 127, 127, -128, 127, -128, -50, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -113, -128, -128, 127, 55, -128, -128, 127, 117, -128, -128, 127, 127, 127, 127, 93, 112, -11, -128, -128, -128, -128, -128, 127, -128, -128, 10, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 47, -128, 6, -128, -128, -116, 127, -128, -93, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 39, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -8, -128, -128, -128, 127, 127, -76, -128, -128, -128, -128, -128, -128, -128, 37, -128, 127, 127, 127, 43, 127, 127, 127, -128, 124, 127, 127, -95, 47, 127, 127, 127, 127, 127, -102, -128, 127, 127, 127, 33, 127, 127, 127, -128, 45, 127, 116, 127, 127, 127, -128, 127, -42, 127, 18, -128, 127, 127, -2, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -16, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 6, -128, 127, 127, -121, -128, -128, 127, -128, 69, -128, 127, -128, 127, -76, 127, -128, -128, -128, -22, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -121, -128, -128, -128, -101, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 109, -128, -95, -128, -100, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -32, -128, -128, -128, 127, 127, 107, -128, 127, 127, -57, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -42, 127, -128, -128, -128, 127, 69, 127, 113, 127, 127, 127, 127, -128, -128, -128, -128, -128, -81, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -121, 7, -128, -73, 18, 127, 127, 127, -128, -128, 127, 127, -128, -128, -48, 127, -128, -128, -128, -128, -128, 127, -6, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -106, 127, -128, 127, 127, 127, -128, 127, 127, 113, -128, -88, 39, -128, 127, -128, -98, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -11, -128, 127, 127, -128, -128, 123, 127, -128, 127, 108, 127, 127, 127, -128, 127, 127, -128, -128, 59, 127, 127, 103, 127, 107, 127, -128, -128, -128, -128, 39, -128, -128, 53, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 73, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 66, 127, 127, 111, -128, -128, 127, -128, -128, -128, -128, 66, -128, -128, -118, -76, -128, -60, 127, -57, -39, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -79, -128, 127, 127, 127, 127, 114, 10, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 43, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 36, -128, 11, -21, 127, -128, 44, 127, -27, -128, -128, 127, 13, -128, -128, 127, 127, 49, -128, -116, 127, -128, -128, -128, -128, -128, 127, 127, 91, 127, 127, 127, 127, 127, 127, 127, 127, -123, 102, -128, -128, -52, 127, -38, 127, -128, 24, -128, -128, -128, -68, 127, 127, 127, -128, 127, 127, -128, -128, 127, 54, -128, 90, -128, -128, -44, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 71, -118, -68, -128, 127, -128, -128, -128, -128, -128, -128, -128, -27, 127, 127, -128, -128, 127, -128, -128, -128, -128, -80, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -98, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -44, 127, 127, -128, -128, -47, 100, -128, -128, -128, -128, -128, 97, 127, 127, 127, 127, 127, 127, 28, -128, 127, 127, -98, 127, 127, 127, -128, 43, -36, -128, -128, -128, -128, -128, -128, -39, 127, -86, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 32, -128, -128, -128, -128, -128, -128, -128, -1, -80, -12, -128, 12, -29, -128, 127, -128, -128, -128, 38, -128, -128, 127, -128, -128, 29, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 44, -128, 127, -128, 127, -29, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 2, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 10, 6, 127, -128, -128, -128, 127, 127, -128, -128, 34, -128, -128, -128, 33, -128, -128, -81, 65, -128, -128, -128, 127, 127, -128, -128, 127, 127, -71, -128, -93, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 15, -128, 127, 127, 127, 127, 55, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -65, -128, -128, -128, -128, -128, 2, 127, 45, -128, -128, 27, -128, -128, 86, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -116, 127, 127, 127, 127, -32, 127, 127, -128, -128, 127, 127, -128, -71, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -100, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -8, 127, 127, 127, -128, 127, 31, -128, -128, -128, 127, -128, 64, -128, 127, -128, -128, -128, -128, -128, -128, -38, 86, -96, -128, -79, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 59, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -31, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 2, 10, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 88, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -24, -128, -27, 127, 127, -68, 127, 127, 127, 127, 127, -128, -8, 127, -128, 127, -128, 127, -128, 127, 73, 127, -128, -128, 127, -128, 11, 127, 127, -128, 27, 127, 11, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -49, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -52, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 45, -128, 127, 127, -103, 127, -128, 127, 127, 127, -44, 127, 27, 127, -128, 127, -128, -128, 102, 29, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 64, -128, 127, 127, 127, 127, 127, -128, 127, -128, 28, -87, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -111, -128, 127, -128, -128, -128, 127, 0, -128, 127, 127, -128, -47, 127, -128, 45, -68, -128, -128, -128, -128, -128, 53, 127, -128, -128, 127, -128, -128, -75, 127, -128, 127, 127, 127, 127, 127, 127, 23, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 2, -128, 127, -128, -24, -128, 127, -128, 127, -128, -128, 24, 127, 127, 127, 127, 127, 127, 127, -64, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 5, 127, -128, -128, -128, -128, 127, -128, -18, -128, 127, -128, 127, 103, 127, 127, -128, 127, 127, -128, -128, 127, -63, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -39, -128, -128, -128, -128, -128, 54, -39, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -98, 127, -128, -128, -24, -128, -128, -128, 127, -128, -32, -128, 127, -128, -128, -128, 127, -128, -128, -22, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -2, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -6, 127, -128, -128, -128, 36, -128, -128, 127, 127, 21, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -48, -128, 127, 127, -128, -128, 127, -71, -128, 127, -128, -128, -128, 98, 127, 127, 49, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 29, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -73, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -3, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -65, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 12, -128, -128, -128, 68, 127, 127, -107, 127, 127, 127, -128, -106, -128, 127, 127, 127, 127, 127, 127, 127, 7, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 88, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 24, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 78, 127, -128, 127, -128, -53, -95, -128, 66, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -54, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 54, -128, -43, -128, 127, 127, 127, -128, 127, 127, -128, 42, 127, -128, -128, 127, -79, -128, -59, 127, 127, 124, -128, 127, -128, -128, -128, 127, -54, 36, 127, 127, -128, -128, -128, -128, -128, 103, 127, 127, 127, 127, 127, 127, -128, -119, -128, 114, -128, -128, 127, 97, -128, -124, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 7, -128, 127, 127, 127, -128, -128, -128, -128, -128, -79, 127, 127, 127, 127, 127, 98, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 33, 127, -57, -128, -53, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -52, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -116, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 123, -128, 127, 23, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -32, -128, -128, 3, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 93, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 29, 127, 45, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -97, -27, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -87, 127, -128, 127, 36, 127, 76, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 50, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 32, -128, -128, -128, -128, -128, -128, 127, -33, 127, -128, -12, 60, 24, -128, -91, 29, 127, 33, 127, -34, 127, 109, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -33, 127, -107, -128, -65, -128, -128, -128, -128, 1, 119, -43, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -37, -128, 0, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -10, 127, 76, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 3, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 2, -128, -128, 16, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -15, -128, -128, -128, -128, -128, -128, -44, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 11, -128, -88, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 27, -10, 127, 127, 127, 127, -73, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -18, 127, -128, -128, -128, 127, -128, 109, -128, 127, 127, 127, -128, 127, 55, -128, 127, 127, 127, -128, 127, 127, -70, -128, 127, 127, 127, 127, 127, -128, 91, 127, 127, -128, 127, 127, 127, -106, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 93, -128, -49, -128, 43, -128, -5, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 91, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 123, -128, 127, 127, 127, -128, 127, -128, 127, -128, 111, 10, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 2, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -29, -128, -128, -128, -128, 127, 107, -128, -128, 127, -128, -128, 13, 69, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -33, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 102, 116, 127, 127, 127, -117, 127, 127, -128, -13, -128, -128, -128, -15, -128, -128, -128, -128, -128, -128, -128, -128, 127, 1, -128, -128, -43, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -6, 127, 127, 127, 127, 0, 127, -128, 127, 13, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 23, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -29, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 43, 127, 127, 127, -128, 127, 36, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 10, -128, -128, -128, 127, -128, -64, -128, -128, -128, -128, -128, 54, -91, 127, 127, 127, -128, 111, -128, -128, -128, -128, -128, -128, 88, 127, -128, 127, 127, -128, -128, 34, 45, 127, -128, 127, 127, 127, -128, -106, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 54, 127, 127, 127, 127, 127, 127, 127, 70, 2, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 117, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 45, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -78, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 93, -128, -128, -101, -128, 90, -128, -53, -98, -26, -128, 127, -44, 127, -128, -128, -128, -36, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 42, -128, -128, -128, 97, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -44, -128, 127, -128, 3, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 73, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -69, -128, 127, 127, -29, -128, -128, -50, -90, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -15, -128, -128, -128, 31, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -43, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 96, -128, -93, -128, 127, -128, 127, -128, 127, -128, 118, -128, 127, -128, -128, -23, -128, -128, -128, -91, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 87, 127, 127, -117, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 98, -128, -128, -11, -128, 127, 127, 7, -128, 31, -128, -128, -128, 44, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 0, 127, -26, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 47, 119, -128, -128, -114, 127, 7, -128, 8, 127, 127, -128, -128, 86, -128, -128, -128, -128, -128, -128, 74, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 11, 127, 121, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -1, -128, -128, 127, 127, -92, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 49, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 11, -128, -128, -128, -128, -128, -128, 106, 127, -128, -128, 127, -103, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 76, 127, -128, -42, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 45, -128, -128, -128, 127, 127, 127, -128, 98, -128, 60, -128, -128, -128, 78, -128, 127, 127, 127, 101, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 58, 127, -128, 127, 127, 111, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -113, -128, 6, -64, -128, -128, -128, 1, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -80, -128, 127, 127, 127, -53, -15, 127, 90, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -43, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 123, -128, 127, 127, 97, 127, 127, 127, 127, 127, 127, -123, -128, -128, -128, -128, -128, 63, -128, -128, -128, -2, -128, 27, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -127, -128, 65, -128, -128, -128, 127, 127, -128, -74, -128, 127, -128, -128, 127, -107, 127, -18, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -114, 127, -71, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 91, -22, -128, -128, -128, -128, -122, -128, 127, -128, 97, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -106, 127, -128, -123, -128, -128, -128, -128, 127, 95, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 0, 127, 127, 127, 111, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 23, 127, -128, 127, 117, 127, -128, 127, 48, 127, -128, 127, 36, 127, -128, 127, 127, 127, -128, 127, 127, -53, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -113, -128, -128, -57, 127, -47, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 23, -128, -128, -128, -79, -128, -128, -128, -128, -128, -128, -128, 57, 127, -128, 127, 103, 127, -128, 127, 127, 127, -128, 127, 127, 127, -97, 127, 127, -128, 127, -12, 127, -128, 127, -64, 127, 2, 127, 127, -128, -128, -128, 127, -128, 7, -128, 127, -128, 127, 127, 127, 127, -117, 127, 127, 127, -128, 127, 127, 0, 127, 127, -128, 127, -128, 1, -128, -128, -128, -128, 127, -128, -102, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 43, -44, 127, 127, 127, -128, 127, -128, 127, -128, 127, 17, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 101, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 3, 127, -128, 119, -128, -128, 127, -128, -85, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -31, -128, -128, -128, -128, -128, -128, 127, 127, -90, -128, 127, -128, -128, -128, -128, -128, -128, 11, 108, 127, -21, -128, 119, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 18, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 109, -128, -128, -128, 127, -128, -128, -128, -107, -128, -128, -54, -128, -128, -128, 127, 6, -128, 127, -128, 127, 127, 127, 127, 86, 127, -34, 127, -123, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 39, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 11, -128, -128, -128, 73, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -119, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -33, 127, -128, 127, 47, -75, -128, 86, -128, -128, 127, -128, -128, -128, 1, -128, -128, -128, -128, -128, -128, -128, -128, 127, -59, -68, 127, 127, 127, 127, 127, -128, 127, 122, 127, -39, 127, 127, 127, 127, 127, -85, 90, -128, 127, -128, -113, -128, -128, -128, -128, -128, 63, -128, -27, 109, 127, 42, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -42, -128, 127, -76, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 90, -128, -128, 127, -128, -128, -128, -128, -128, 39, 127, 127, 127, -50, -128, 127, -128, -128, -128, 127, -128, -128, -52, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -96, -128, 127, 102, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 95, -128, -128, 127, -128, -128, -128, -128, 96, -28, 127, 127, 127, -95, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -8, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 8, -128, -128, -128, 127, -128, -128, 127, 45, -128, -128, 127, -128, -128, -118, -128, 45, -128, -128, -128, 127, -100, -128, 127, 127, 32, 127, 127, 127, -128, 127, -128, -128, -128, 127, -58, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -38, -128, -16, 127, 127, 127, 127, 127, 127, -128, 127, 53, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 79, -128, 127, -2, 127, -128, 127, 127, 127, 48, -117, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 119, -128, 127, -97, 127, -128, 127, -128, 127, 127, 103, 127, 127, -13, 123, 127, -128, -128, 127, -128, 127, 127, 127, -16, 127, 127, 127, -128, 127, 57, 13, -128, 127, 127, -128, -128, -128, -128, -128, -79, -128, -50, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -66, 127, -128, 127, 0, 127, -128, 127, -128, 127, -128, 108, -128, 127, 127, 127, -128, 127, 127, 118, -128, 31, -128, -128, -128, -128, -128, 127, -128, -68, -128, 127, -116, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 65, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -85, 127, -109, 10, -128, -121, -128, -128, -128, 127, -128, 127, 96, 98, -128, -128, -128, -128, -128, -124, 60, 127, -85, 127, -128, -128, 127, 73, -128, 68, 127, 127, -128, -128, 127, 102, 127, 127, 127, 127, 127, 127, 127, -63, -128, -71, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -24, -128, -128, -128, -108, -128, -128, 127, 127, -128, 123, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -45, -128, 127, -128, -90, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -100, -128, 127, -128, -55, 127, 127, 50, -5, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -3, -128, 127, 127, -128, -128, 127, 127, -24, -98, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 33, -128, -128, -128, -128, -96, -128, -128, 127, 127, -128, -88, 127, 50, -128, 127, 127, -128, 71, 127, 127, 127, -43, 37, 127, 127, 127, -23, 127, 127, -128, 2, -128, -128, -128, -128, -128, -128, 37, -128, -128, 127, -128, 114, 127, 127, 91, 127, 127, 127, -128, 127, 127, 127, -68, 127, -128, 127, 127, -74, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -12, 122, 127, 127, -128, -128, -91, 127, -128, 127, -128, 91, -128, -128, -128, -128, -128, 47, 127, 127, 127, 127, 127, 127, -128, -128, -55, 127, -128, -128, -69, 127, 38, -128, -128, 34, -128, -128, -128, -128, -76, 127, -128, -128, 127, 127, 127, -128, 127, -128, 16, -128, -128, -128, -6, -128, -128, -128, 127, 127, 0, 127, 127, 127, 127, 127, 71, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -47, 127, -128, 127, 127, -33, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -123, 127, 127, -128, 127, 127, 127, -128, 127, -128, 3, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -58, 106, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -1, -128, 127, -128, -128, 58, 127, 127, 127, 127, 127, 127, -128, -128, -128, 0, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -39, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 47, 127, -128, -128, -128, -128, -128, -128, 60, -15, 127, 127, 127, -128, -128, -109, -128, 45, -128, -128, 127, -128, 23, -75, 127, 127, 127, -128, -128, 127, -128, -128, -128, -36, -124, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 117, 127, 127, 127, -128, 98, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -24, -128, -128, 0, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -58, 95, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -74, -128, 127, -128, 127, -128, -128, -128, -96, 127, -128, -128, 127, -11, -128, -128, 127, 0, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 53, 127, -2, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 109, 127, 127, 13, 127, 127, 127, 127, 127, -123, -128, 127, 97, -128, -128, 127, 127, -128, -128, 75, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 10, -128, -128, -128, 127, 127, 127, -122, 127, 127, -128, -128, 127, 127, 127, -128, 0, -128, -128, -128, -128, -128, -128, -128, 0, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 59, 127, -128, 127, 127, -128, 127, 111, 127, -128, 127, -10, 127, -128, -128, -128, -128, -128, 127, 127, -95, 127, 127, 127, -128, 127, 127, 127, 90, 127, 127, 127, 127, -71, 127, 127, 127, 127, 116, 127, -128, -128, -128, -128, -128, -128, 127, 127, 13, 127, 127, -128, -128, -128, -128, -128, 12, -128, 127, 127, -128, -128, -3, -128, 48, -128, 31, -29, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 95, -128, 127, 127, -128, 112, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -11, 7, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 70, 127, 127, 127, 127, -128, -128, 59, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 106, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 23, -128, 127, 127, 39, -85, 127, -128, -128, -128, -128, -128, -128, 127, -32, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -29, 127, -10, 127, 127, 117, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -76, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 31, -128, 127, -50, -128, -128, -128, -128, -85, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 73, -34, -128, 6, 127, 127, -128, 127, -10, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 7, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -34, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -8, 127, 127, 127, 127, -37, 127, -128, 98, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 34, -128, -128, -128, 127, 127, -128, -128, -128, 127, 24, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -102, -29, -128, 111, 28, 127, 127, 127, 127, 127, 127, -128, 127, -128, -101, -128, -128, -128, 127, -128, 127, -97, 58, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -116, -128, 127, -128, -128, -128, -52, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -124, 127, 113, -128, -128, 127, 124, -128, -128, -128, -128, -128, -128, 127, -128, -86, 3, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -43, 74, -22, 127, -128, -128, -128, -128, -128, 100, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 122, -128, 127, -128, -128, -128, 127, 79, -128, 127, -96, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 118, 127, -128, 8, 127, 127, 127, -128, 74, -128, 127, -128, -128, -128, 127, -128, -128, 11, -128, -128, -128, -128, -128, -128, 127, -90, 53, -50, -128, -128, -128, -128, -128, -128, -57, -128, 127, -128, -128, -128, 127, -128, -13, 53, 127, 127, 127, 127, 127, 127, 127, 24, -128, -128, 114, 127, -17, 127, 127, 127, 50, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -47, -128, -128, -128, -128, 127, -128, -39, -128, 127, -128, 127, -2, 97, 124, 127, 127, 127, 127, 106, 127, 42, 127, 127, 127, 127, 127, 92, -128, -29, -128, -128, -128, -128, -128, -128, 6, -128, 127, 127, 127, 127, 127, 127, 127, -128, 2, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 58, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 23, -128, 127, 28, 127, 79, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 80, -50, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -81, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 31, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -29, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -32, -128, 127, -128, -128, 127, 127, -59, 127, 127, 127, 127, 127, -79, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -15, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -33, 127, 127, 127, -100, 100, -128, -128, -128, -100, -128, 127, -128, 127, 0, 113, 45, 127, -88, -128, 71, 127, -128, -128, 127, 57, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -38, -128, 127, 127, 127, -128, 80, 127, -128, -128, 127, 127, 127, 64, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 3, -128, -128, 127, -128, -128, -128, 127, -128, -55, 127, 0, 112, 127, -128, -128, -128, -128, -128, -128, 88, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -63, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -33, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -31, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -26, 127, 127, 127, 127, 127, 127, 127, 127, -59, 127, 127, -128, -128, -128, -58, -127, 127, -128, 127, 127, -128, -128, -128, -128, -28, -128, -128, 127, 127, 127, -34, 0, 127, 127, 127, -128, 127, -128, 34, -128, -128, -128, -128, -128, -128, 23, -128, 102, 113, -128, -128, 127, -128, -128, -123, 127, -128, -128, -128, -128, -128, -88, -128, -128, -128, 63, -128, -128, -128, -128, -128, -128, -128, -128, -128, -5, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -75, 127, 127, -128, 127, 127, -100, -128, 127, -128, 127, -128, -1, -97, 127, 127, 81, 127, 127, 127, -128, -85, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 50, 127, -5, 127, 127, 127, -128, 127, 2, -128, -128, -128, -128, -128, 0, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 58, 127, 127, 127, 127, 127, 127, 127, -128, 86, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -73, 127, 127, 48, 127, 22, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 27, -128, -128, 127, 127, 127, -128, 33, -128, -128, -128, -128, -128, 108, -128, 127, 127, 127, -128, 127, 127, 127, 108, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 29, -107, -128, -128, -128, -128, -128, -128, 127, -128, 127, -47, 127, -71, 127, 127, 127, 127, 127, -128, -100, 127, -128, 127, 90, 127, -128, 127, 127, -128, -128, 127, 127, 93, -128, -128, -95, 70, -65, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 85, 127, 127, 127, -71, 127, -106, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -44, 127, -128, 127, 127, 127, 127, 127, 127, -128, -114, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -73, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -57, -128, 127, -128, -128, -128, -128, 127, -128, 53, -128, -128, 127, -78, -128, 127, 127, 127, 127, 127, 127, 127, 127, 59, 127, -128, 127, -128, 33, -128, 127, -128, -128, -128, 127, -128, 127, 102, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -28, -128, 127, -128, -128, -128, -36, -17, -128, 1, 127, 127, 127, -128, 13, -128, -37, -128, 3, 127, 127, 127, 127, 127, 127, 127, 121, -128, 127, 39, 127, 118, 127, -128, 127, -128, 127, 127, 127, 127, 12, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 52, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -111, 127, 127, 127, -128, -128, 127, -128, -128, -66, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 53, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -111, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -44, -128, 127, -128, 127, 127, -128, -128, 23, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -95, -128, -109, -128, -128, 98, 127, -128, -22, -92, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 17, -15, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -109, 127, 127, -128, -128, -128, -128, -128, -103, -128, -128, -128, -128, -128, -128, 127, -128, 127, -74, -15, -128, -128, 127, -128, -128, 127, 127, 127, 64, -128, -128, -128, -128, -128, -42, -128, 127, -128, 127, 127, -128, -128, -63, -128, -128, -128, 127, 127, -128, -39, -128, 127, -128, -128, 37, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -3, 33, -128, -128, -70, 127, -128, -128, 127, 127, -128, -128, 127, 79, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -39, 127, 127, -128, -18, -128, -128, -128, 127, -128, 127, -128, 86, -128, 127, -128, 127, -128, 81, -128, 127, -128, -128, -128, 127, 21, 127, 127, 127, 127, -128, 127, -57, 127, -128, -68, 127, 127, 22, 0, 127, 127, 17, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 45, 127, -98, 127, -128, 127, 102, -128, -128, -128, -128, -91, -29, 127, 5, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 38, 127, -128, -128, -128, -128, -128, -75, -128, -128, 127, 127, -128, 127, 127, 7, -128, -128, -128, -128, -128, -128, -128, -128, 87, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -1, -128, 18, 127, 127, -106, 127, 127, -128, -128, 17, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -36, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 0, 127, 127, -128, -128, -128, -128, -128, -128, 127, -6, 127, -128, 127, 127, 127, 73, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 121, 127, 127, -85, 127, 127, -128, -128, -128, 21, -128, -128, 127, 127, 127, -128, -128, 127, 59, -128, -128, 127, -128, 127, -128, 127, 55, 127, 127, 127, 96, -128, -74, 90, 87, 127, 127, 127, 127, -128, -80, -128, -128, -128, -128, -128, -128, 127, -128, -66, 127, 127, -128, 127, 127, 127, -57, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 59, -38, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -1, -27, -128, 127, -128, -101, -26, 127, 127, 127, 127, 127, 109, 127, 121, 127, 127, 111, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 18, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -76, 127, 127, -108, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 124, 127, -64, -128, -92, 127, -128, -118, -128, -128, -128, -8, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -43, 97, -128, 127, 127, -103, 127, 127, 127, 127, -128, -98, -47, -31, -128, -128, -128, -128, -128, -128, -128, -128, -128, 122, -128, -128, -128, -128, -128, -128, -128, -128, 59, -128, -128, 127, -38, 127, -128, 127, 127, 127, 31, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -75, 127, 127, -128, 44, 127, 127, 127, -128, 127, 102, -128, -128, -128, -128, -128, -128, -128, -128, 127, -48, 127, 127, 127, 127, 127, 127, -128, 127, -128, 118, 0, 127, 97, -128, 127, 127, 127, 127, 127, 127, 127, 127, 37, 127, 127, 127, -128, 127, 127, 127, 69, 124, 127, 127, -128, -128, 127, 127, -128, 127, -128, -24, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -78, -128, -128, 0, -128, -8, -128, 127, -128, 24, -128, 127, 127, 127, 127, 127, 127, 127, 127, 27, -128, 127, -128, -128, -128, -128, -91, 127, -128, 22, 127, -128, -128, -128, -128, -128, -128, -128, -31, -128, 127, 127, 127, 127, 127, 38, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -12, 27, 127, -128, 34, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -87, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 57, 127, 127, 127, 127, 127, 127, -22, 127, 127, 64, -128, -128, 127, -128, -128, -128, -128, -128, -128, 12, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -31, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -118, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 26, -128, -128, 127, -128, 127, -128, 127, 127, 127, -119, 127, -128, 127, 127, -128, 127, -3, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 49, -128, 127, -128, 127, 113, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 39, -128, 127, 73, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -59, -128, -111, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -106, -128, -128, -128, -58, -128, -128, 127, 90, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -68, -128, 127, -128, 127, 93, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -63, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 117, -112, -128, 127, -124, 127, -128, 127, -128, 127, -33, 28, -5, 127, 127, -26, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 22, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -47, -128, -128, 127, 69, -128, -128, 127, -128, -128, 127, -92, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 69, 68, 127, 127, -128, 127, 127, -37, 127, 127, 42, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 68, 127, 127, 127, 11, -128, 127, -108, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -64, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 38, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -80, -128, -128, -128, 127, 127, -47, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -18, 127, 127, -128, -128, 127, 78, -128, -128, 88, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 101, 33, -116, -31, -123, 33, 127, 127, 2, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -127, -128, -16, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 121, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 22, -128, -128, -127, -128, 127, 127, -128, 3, 127, -128, -128, -128, -11, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 23, -128, 13, -128, 127, 116, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -114, -128, -128, 88, -128, 127, 59, -128, 127, 70, -128, -128, 5, -128, -79, 127, -119, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -68, 127, 127, -92, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -107, 127, 127, 127, -128, 127, 127, 127, 127, 127, -58, -128, -128, -128, -128, -128, -128, -49, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, -118, 127, 127, -128, 127, 127, -128, -95, 127, -128, 88, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -68, -60, -128, -15, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 90, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 123, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -8, 127, 127, 127, 127, 127, 127, 127, 91, 106, 127, -128, 127, -128, 127, -128, 92, -128, -8, -128, 127, 127, -128, -128, 127, 116, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -11, 127, 127, 127, -128, 127, 90, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 15, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -44, 127, 127, 127, 127, 127, 127, 127, 87, -26, 127, -128, 127, -128, 127, -128, 127, -81, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 85, 127, 127, 127, 127, 13, -128, -128, 127, 127, -128, 127, 127, 7, -128, 127, -128, -128, 127, 101, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -42, -128, -128, -128, -128, -128, -128, -128, 127, 106, 24, -128, 127, -128, -128, 127, -128, 127, -128, -13, -128, -28, -128, 96, 127, -128, 127, 127, 127, 127, 127, 127, -128, -119, 87, -128, -128, -128, 127, -128, 127, -117, 127, -128, 127, -128, 127, -128, 47, -128, 127, -128, -55, 7, 66, -128, -128, -128, -128, 127, -128, 127, 127, 127, -34, -53, -128, -128, -128, -128, -128, -128, -128, -128, 95, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 76, 127, -128, -96, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -15, -128, 26, 127, -128, -26, 127, 127, 92, 127, 127, 127, -97, -128, 127, -128, 127, -128, -128, -128, 45, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -45, -128, 127, 127, 127, -47, 127, 127, 127, 127, 127, 127, 127, 127, -79, 127, 26, -128, -128, 54, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 39, 127, -128, 127, 127, 127, -128, 127, 127, 36, 127, 127, 127, -128, 127, 127, 127, 127, 127, -80, -128, -128, -128, -128, -27, 127, -124, 127, 127, 127, -128, 127, 127, 127, -121, -128, 127, 127, -128, -128, 73, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -13, 127, -128, 127, 127, -112, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 24, -128, 127, -128, -128, -128, 16, -128, -128, 127, -128, -128, 127, 7, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -80, 127, 127, 106, -128, 127, -78, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 102, 127, -128, 33, -128, 127, -128, 127, -128, 37, -128, -128, -128, -128, -128, -15, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 0, -103, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -49, -128, -97, -128, 93, 127, 1, 127, 127, 127, -128, 127, -85, -128, -128, 127, -128, -128, 127, 127, -128, -8, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 54, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 22, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 73, 127, -128, -90, -128, -128, -128, -128, 127, -128, -92, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 92, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 100, 127 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
