-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
            -77, -17, 68, 57, -115, -94, 36, -117, 94, -18, 120, 110, 92, 89     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -32, 11, -47, -121, -4, -95, -70, 30, -12, 96, 95, -12, -54, 105, 114, -91, -58, -97, -10, 39, -115, 39, 103, -90, -7, 51, -83, 102, -81, -109, -66, -55, -54, -115, -125, -126, -127, 109, -80, 100, 119, 60, 44, -102, -50, 87, -80, -26, 107, 84, 63, -20, -81, 92, -34, 59, 28, 61, -32, 96, -46, -70, -79, -17, -24, 103, 20, 37, 105, -32, -97, 70, 62, 64, -30, 61, 18, -65, 118, -73, 21, 6, 87, 119, 31, 12, 61, 64, -106, -29, 97, 11, 91, -105, -121, 23, -79, 85, -99, 47, -40, -1, 14, -8, 80, -47, 62, -36, -42, 7, 110, -31, 45, -37, 36, -21, -92, 74, 1, 37, -67, 65, 21, -28, 40, 107, 49, 124, 54, 52, -109, -122, 113, 10, 106, -72, 97, -54, 37, 75, -2, -125, -21, 105, -33, 28, 44, 84, -47, -11, -16, -33, 116, -44, -116, -18, 93, 19, -46, -106, 17, 65, -80, 113, -89, -91, -32, -73, -69, 90, 42, -101, -99, 44, -73, 72, -60, 59, -97, 94, 63, 92, 40, 14, 39, 82, 11, -117, 10, -93, 83, -6, 13, -79, 121, -75, -117, -45, -115, 73, 37, 101, -118, -122, -122, 44, -89, 85, 124, -55, 120, -74, -124, 11, 119, 124, 43, -123, -85, -88, 5, 94, -68, 104, -70, -30, -92, -88, -34, 100, 26, -25, 121, -73, -42, -10, 12, -22, -38, -35, -56, 105, -39, 64, -29, -21, 59, 12, -112, 7, 37, 111, -95, 29, 54, 37, -75, -77, 50, -108, -30, -11, 103, -44, -91, -53, -100, -104, -25, 108, 31, -80, 87, -78, 80, -46, 112, -7, -61, 26, 8, -46, 32, -88, 69, -37, 126, -24, -113, 28, 52, -35, 119, 123, -7, 32, -27, 56, -70, 68, -70, -81, 123, 7, -63, 16, -6, 52, 56, -116, -51, -87, 76, -115, 84, 102, 111, 30, 19, -126, -112, 28, 3, -126, 63, 114, 7, 42, 38, 36, 27, -10, -90, -19, -70, 61, -11, -103, 37, 49, 103, -79, -16, -45, 68, -106, -49, -17, 48, -53, -92, 22, -119, -118, -117, -92, -50, -41, 110, -67, 115, 122, -59, -5, -13, -24, 63, 103, 53, 117, 107, -110, 51, 117, 33, -60, -123, 101, 16, -40, 2, 51, -39, 110, 31, 75, -23, 116, 91, 104, -43, -124, 29, -90, 11, -101, 59, -58, 18, 7, -107, -62, -10, -128, 115, -23, 17, -117, -38, 48, 26, 45, -64, -41, 36, -22, 51, 57, 102, -28, -4, -102, 11, -60, 10, 109, 97, -100, -77, -79, 105, -110, 12, -4, 38, -114, -61, -29, -10, -71, 89, 2, -13, 39, 45, -46, 89, -37, -54, -27, 41, 106, 45, 49, 111, -66, 87, -41, 106, 91, -39, 97, 68, 63, 106, 84, -58, -82, -125, -93, 50, 55, -88, 102, 96, -1, 30, -76, 85, 90, 18, -3, 55, 115, 99, 89, -77, 64, 46, 77, -27, -19, -65, 50, 65, 52, 28, 101, 38, -2, -4, 2, 74, 4, -106, 31, -27, 21, 76, 32, 93, -12, -118, 100, -2, -7, -117, -90, 0, 116, 105, 18, 27, 85, -53, -91, -17, -96, 47, -11, 75, -30, -35, -87, -23, -6, -3, 126, 6, 31, 99, 122, 103, -68, -72, -108, -120, 4, 93, -86, -52, -63, 6, -23, -120, -69, 50, 25, -79, -9, 57, 74, 77, 84, 121, -85, -24, 107, 46, 44, 120, 49, -51, -122, -12, 49, -45, 78, -68, 12, 63, 86, 73, -2, 72, -96, -70, 98, -116, -34, -77, 101, -112, 62, 83, -58, -71, 78, 25, -31, -103, 104, -27, -13, -10, 84, 39, -68, -20, 48, 0, -16, -127, 97, 79, -44, -117, -67, -44, -58, 4, 23, 46, -55, 90, 94, -83, -123, -36, 109, -73, 94, 11, 39, -8, 99, -56, 97, 113, 40, 52, 119, 24, -51, -125, 61, -47, 16, 37, 11, 42, 67, -56, 61, 36, -35, 72, 25, -10, -47, 82, -106, 107, 104, -24, 82, 7, -61, -119, -122, 109, 103, -70, 12, 65, 46, 121, 27, 73, -94, 94, 98, -4, 126, 125, 67, -74, -121, 83, 84, -55, -4, -20, -124, 58, 118, -30, 12, 10, 70, 34, -63, -55, 74, -62, 109, -50, -62, 75, -70, -70, -107, 9, 120, -47, -25, 41, -80, -69, 41, -58, -14, 111, 46, -78, 47, 94, -86, -61, -4, -114, 10, -41, 110, -69, -12, -111, -50, -52, -4, 70, -57, -82, -66, -116, -23, -110, -90, -76, 94, 81, 81, 53, 93, 106, 56, 7, 39, 71, -14, -42, -30, 57, -86, 68, 42, 94, -53, -72, 48, 47, 122, 4, -96, -1, 75, 121, -11, 66, 122, -2, -18, -50, 63, 60, 92, -88, -89, 90, -123, -51, -50, 60, -9, 9, -22, 113, -3, 84, 70, -113, -68, -28, -112, -76, 33, -59, 2, -19, 98, -35, 1, 127, -126, -39, -12, 108, 117, 87, -68, 29, 107, 78, -91, -26, 17, 32, -110, -96, -63, 110, -118, -11, 83, 83, -67, -122, 68, -34, 82, 113, 43, -102, -62, -10, -113, -56, -44, -87, 107, 126, -30, 116, 83, 123, -80, -13, -17, 101, -9, 79, 114, 55, 118, 114, 21, -30, 97, -21, 103, -77, -95, 48, 37, 8, -81, -73, 81, -59, 116, 69, -86, 5, 118, -14, -97, -55, -5, -83, 7, 55, 56, 26, -10, 3, 62, -47, 107, -25, -112, 35, 48, -81, 1, 95, 118, -77, -8, -125, 109, -91, 112, -52, -76, 35, -30, -107, 102, -57, -61, -111, -64, -23, -40, -29, 50, 27, 80, 55, 110, -47, -5, 114, -50, -111, 25, -41, 11, -41, 108, -90, -22, 54, -15, 27, 82, -66, -118, -110, -51, 60, 35, -27, 44, -1, 49, 90, -2, 30, 77, 101, -5, -72, -125, 64, 39, -31, -112, 37, -126, -36, -26, 13, -118, 26, 76, 21, 9, -9, -44, 24, -36, -92, -88, -112, 5, -50, -117, -25, -6, 83, 126, -105, 93, -41, 84, 123, -91, 30, 47, 26, 29, -126, 16, -43, 40, -21, 66, -122, 81, -128, 78, -102, -113, -90, 59, 33, 82, -120, -83, 58, 23, 26, -39, -43, 22, -123, -46, 6, -125, -13, 85, -63, 70, 26, 75, 25, 118, 89, -84, 79, -79, -22, 77, 24, -6, -124, 86, -23, 87, 57, -54, -54, 22, -1, 71, 85, 61, -77, 59, -10, -122, 38, 2, 34, -67, -125, -82, -73, -66, -2, -18, 87, 120, 96, -66, 23, 24, 31, 119, -31, -36, -76, -51, 19, -43, -104, 57, 106, 105, 96, 88, 57, -88, 100, -40, -66, -91, 18, -76, -77, 118, 58, 97, 78, -30, -22, -50, 102, 49, 26, 27, 79, 112, -119, -48, 41, 93, -88, 19, -123, 87, -15, -39, -12, 9, -94, 4, 5, -25, -4, -101, -73, 43, -47, 17, 43, -21, 99, -80, 65, 116, 26, 74, 32, -46, -39, -21, 0, -58, -20, 69, 78, -35, 113, -69, -85, -80, -110, -124, -49, -126, 70, -43, 75, 98, -10, 74, 121, -117, 60, -101, -110, 89, 6, 30, -67, 78, -23, -70, -23, 106, -122, 113, -107, -112, 62, 82, -37, -96, -43, 101, 33, 93, 17, -85, 101, -122, 52, -109, -31, 114, 19, 17, -10, 92, 49, -37, -2, -29, 61, 73, 57, -3, -7, -11, 68, 40, -87, -29, -89, -59, -33, -16, -13, 112, -120, -111, 22, 121, -55, -115, -106, -93, 97, -71, 25, 122, -82, 80, -42, -128, 26, -44, 89, 25, 27, 99, -128, 113, 63, -44, -123, -11, -54, -49, 10, 85, 3, -93, 95, 32, 60, 31, 63, -9, 121, 0, -115, -19, 4, 1, -15, -84, -83, 112, -108, -79, -35, -83, -78, -41, -54, -28, -38, -60, -91, -97, 46, -104, -104, -4, -57, 40, 78, 73, 81, -96, 16, 99, 70, -113, 78, 33, -90, 0, 12, -74, -53, 51, -3, 116, 52, -19, -114, -86, 14, 81, -68, 6, -123, 17, -82, 16, 91, -71, -14, 37, 97, -122, 45, 19, -67, 11, -33, -34, -14, 66, 94, 69, -106, -118, 112, 39, 18, -69, -116, 88, 58, -36, -117, -40, -119, -40, 66, -110, -9, 21, 42, 49, 65, -110, -77, -126, -54, 9, -99, 7, 20, 23, -111, 18, 82, -27, 26, -122, -54, 107, -97, -95, -78, -14, -27, -107, -37, 45, -92, 110, 86, -48, 120, -109, 47, 35, -22, 19, -50, 99, 76, 29, -83, -120, -62, 96, 109, -116, -71, -79, 78, -67, -114, -47, -26, 36, -105, 98, -51, 2, 30, 78, 122, -102, -104, 71, -125, -22, -22, 32, 1, -50, -35, -10, 37, -110, 107, -64, -92, 44, -3, 124, -67, 21, 120, -61, 70, -13, 108, 100, 64, 32, -30, 74, 33, 95, -32, 2, -107, -44, 126, 54, -27, 21, 26, -9, -126, -26, -66, 74, 90, 15, -121, -127, 110, -119, -69, 46, 51, -40, -82, 112, -7, 23, 39, 34, -59, -123, 10, 26, 41, -98, 121, -82, 66, -90, -87, -69, -88, -29, 127, -67, 34, -126, -69, 18, -108, -7, -53, 93, 55, 8, 21, 11, 47, 84, 99, 88, -48, 74, -118, -8, -88, 91, 98, -63, -87, -80, 31, -39, 57, -21, -87, -54, -94, 62, 86, -94, -50, 97, 97, -97, -24, -43, -17, -9, 32, 127, 36, 21, 115, -127, -23, 118, -60, -64, -114, 112, -81, -63, -10, 2, -115, 4, -26, 0, 109, 89, 32, -38, -63, -116, 73, 39, 59, 63, 29, 60, -28, 95, -86, -72, 87, -83, -85, 104, 92, 27, -106, 60, 50, -82, 84, -39, 43, 115, 54, 126, -46, 81, 36, -113, 68, 98, 28, 36, -68, -72, 96, 80, -75, -6, 7, -60, 68, -62, 48, -63, -85, 8, -12, 81, 3, -92, -77, -69, 57, -55, -101, 125, -75, -109, 54, 53, -26, -13, 26, -18, 7, -14, -124, -21, -107, -31, -30, -118, 29, 16, -59, -109, -101, -110, 21, -108, -114, 19, 88, -41, -112, 87, 4, 41, -121, -13, -80, -57, -13, -47, 35, -119, -128, 26, -36, 123, -109, -58, 112, -27, -48, 121, 114, 14, -126, 51, 50, -116, 11, 84, -107, 5, -42, -59, -50, 52, -89, 17, -115, 73, 44, 20, -120, -116, -112, 48, 7, 61, -122, -17, 97, -62, -15, -21, 125, 18, 56, 30, 15, -61, 77, 127, 68, 35, -73, 94, -25, -117, 100, -4, 105, 95, -4, 49, 123, 118, -49, -27, -86, 1, 55, -30, 104, -58, -117, -55, -14, 94, -36, 78, -5, -9, -125, 61, 4, 84, 51, 60, -22, -88, -7, -100, -64, -30, 65, -11, 61, 116, 15, 10, 64, -55, 45, 116, -12, -100, 96, 72, -75, -70, -20, -26, -70, 56, -84, 73, 97, -119, 107, -21, 69, -38, -96, -54, -37, -109, -66, -112, 51, -66, 60, 28, -64, 0, -43, 40, 9, 16, 61, 102, -33, 110, 75, 58, -2, 40, 42, 122, 19, -53, 103, 100, 46, 76, 79, 91, -11, -26, -46, 88, 121, 38, -122, -5, 39, -116, -7, -65, -91, 90, -21, 20, 23, -69, -79, -16, -28, 51, 2, 105, 115, 28, 104, 79, -44, -44, -117, 58, -76, -53, -101, -107, 34, -112, 71, -104, -65, 79, -122, 70, 59, -2, -92, -39, -66, 32, 112, -112, -110, 19, -47, -103, 113, 102, -82, 46, -10, -60, 30, 110, -95, -119, 8, -69, -37, -88, -42, -60, -1, -33, 15, -34, -12, -41, -118, -52, -115, 13, 109, -23, 83, -50, 115, -95, -92, 63, 70, -49, 57, 27, -6, 42, -37, 7, -107, 39, -36, 19, 102, 63, 41, -14, 5, 111, 3, -27, -20, 115, 74, -35, -15, -2, 1, 101, 43, -126, -38, -110, 4, 111, -76, -99, 23, -1, 11, 3, -1, -20, -25, 43, -37, 70, -68, 92, -90, -56, -29, -63, 80, 126, 3, -50, 54, 90, 104, 0, 66, -107, -124, 2, -94, -25, 80, -69, 83, -91, -10, 59, 47, -101, -118, -113, -75, 108, -117, -112, -97, -85, -2, 107, -68, 19, 53, -62, 121, 100, 25, 98, -95, -33, -109, 9, 71, 72, -85, -24, 3, 118, -88, -58, -94, -66, 63, -22, 108, 101, -80, -35, -76, 30, -96, -102, -31, 106, -65, -93, -123, -96, -19, -50, 12, -41, -3, -38, -93, -124, 35, 19, -56, 61, 8, -107, 122, -117, 17, 98, 13, 17, 87, 94, -62, -82, -36, 50, -58, 61, -127, 92, 43, 24, -94, -76, 15, -103, -101, 75, 14, 94, -47, -81, 28, -95, -70, -110, -85, -112, 90, -17, -98, -38, -57, 111, 28, -62, 122, 81, -7, 110, -72, -47, -73, -109, -124, -11, -50, -48, -17, -95, -125, -128, -77, 28, -70, -34, 65, -66, -20, -42, 58, -54, 29, 37, -53, 79, 92, -124, -9, 107, -22, 80, 24, -104, -28, -53, 80, 30, 63, 31, -109, 120, 121, -36, -67, 38, -50, -35, 75, -54, 6, -85, 30, -6, -24, -33, 2, -30, -124, -123, -33, 31, 44, 85, -99, 15, -100, 96, 108, -23, -115, 47, 95, -71, 2, 25, -33, -85, 24, 36, -41, -26, 120, -8, 81, -72, -100, 22, 115, 3, 55, -44, -52, -84, -7, 75, 92, 39, -42, -34, -91, 25, 70, 13, 58, -3, 105, 121, -26, -7, 48, 87, -13, -96, -107, 92, -67, 42, -120, 82, -21, -22, -54, -74, 106, -119, 88, -114, 86, -86, -76, -35, 21, 97, 97, -112, -106, 10, -102, 82, -78, 114, 42, -107, -121, 31, -19, -2, 99, 85, -125, 71, -63, 55, 2, -109, 28, -118, -6, -18, 33, 49, -116, 35, 84, 126, -83, -17, -45, -73, -85, 76, 17, -121, -67, 59, -2, -54, 22, 87, 53, -20, -40, -59, -76, -124, 65, -89, 92, 81, 3, -58, 13, -21, 13, 97, -33, -61, -20, 126, 0, 67, 113, 56, 115, -80, -57, 51, 78, -59, 60, 63, 17, 44, 89, 41, -124, -87, -97, 21, -75, 88, 119, 118, 67, 69, 17, -41, -112, -96, 119, -39, -127, 109, -33, -60, 114, -48, -24, 67, 102, -120, 64, -117, -59, -4, -61, 82, -11, 86, 5, -104, -11, -36, -79, -42, 38, 64, 44, 118, -116, 71, -20, 116, -74, 87, -16, -124, -81, 84, 21, -53, 28, 124, 58, 67, 22, -58, 74, 73, 89, -88, -51, -45, -42, 47, -44, 24, -107, 64, 111, 116, 120, 8, -58, -31, -75, -122, -105, 114, -51, -74, -85, 62, 85, -4, -103, 29, -87, 5, -41, -11, -84, -104, 110, -24, -2, -89, -124, 16, 96, -52, -53, -12, 62, 95, -96, -98, 29, -21, 54, 123, -110, -93, 100, -3, 60, 54, -60, 112, 12, -25, 87, -100, -46, 109, 19, 80, -44, 29, -79, 46, -115, 29, 75, 120, -127, -65, -67, 68, 23, -10, -22, 88, -27, -91, 89, -88, 10, 25, 127, -93, 49, 29, 0, -113, 60, 25, -72, 91, 38, -31, 12, -78, -119, -104, 120, -45, -46, -86, -100, -75, -90, -72, 109, -83, 119, -103, 11, 97, -37, -124, 123, -24, 36, -40, -62, -85, -32, -46, 96, 97, -95, 121, 24, -54, 49, 105, 39, -106, 21, -72, -20, -30, 21, 25, 77, 19, 110, -106, 40, -47, 107, 37, -36, 77, -111, -38, -128, -12, -57, -46, -89, -85, -57, 112, -29, 43, 62, 59, 33, -68, 2, -25, 67, 94, -24, -36, -57, -121, -70, 113, 102, -26, 23, -119, -26, -115, -83, 67, 125, 75, 14, 29, -16, -71, 19, 64, -93, 105, -27, 60, -42, 127, 81, 29, -42, -127, -8, 20, 29, -68, 82, -28, 125, -107, 65, 6, 104, 80, -46, -99, 110, 123, 43, 72, 38, 19, -81, -114, -100, -2, 57, 103, -88, -96, -103, 97, -17, -113, -58, -19, -50, 111, -112, 5, 46, 127, 46, -116, 99, 96, 31, 15, 34, 64, 13, -74, 68, 13, 125, -18, -59, 87, -76, 86, 125, -8, -38, -112, -49, -24, 118, -85, -117, 65, -74, -78, -27, -79, 123, 87, 85, -69, -34, 33, -41, 63, -80, -123, 39, 61, 15, 64, 115, 122, 7, -62, -98, -109, -123, 102, 59, 109, 70, 104, -30, 9, 49, 69, -14, 4, -116, 126, 88, 25, -36, -65, 21, 18, 7, 82, 121, -88, 122, -114, 22, 48, -98, 49, -53, 112, -70, -109, 53, 44, 95, 64, -36, 91, 126, 62, 54, 117, 107, 87, 76, -83, 109, 123, 124, 99, -13, -24, 35, -116, 98, -16, -33, 71, 17, 99, -42, -64, -36, -21, -95, -36, -76, -95, -96, -54, 49, 56, -19, -121, -4, 105, 11, 71, 33, 43, 40, -1, -109, 6, 36, 24, 86, 11, -7, -19, 109, 3, -47, -114, -7, -55, -47, 62, -17, 100, -22, 40, 63, 110, -89, -105, 65, -118, -109, 50, -119, 5, -29, 67, -95, 77, 85, -98, -109, 77, -82, -3, 34, -32, 106, 83, -33, -83, 31, 72, 76, 48, 91, 122, -76, 5, -36, -123, -51, -12, 47, -13, 35, -110, 20, -46, -115, -78, 44, -59, -38, -109, 14, -75, -17, -25, -73, 17, 82, -106, 36, 56, 51, 75, 100, -77, -75, -81, -21, -60, 25, -10, -19, -29, 43, 52, -4, 4, 6, 95, 7, 93, 104, 68, 34, -89, -81, 22, 20, -93, 72, -98, 34, -119, -24, 112, 30, -51, -1, 32, -95, -123, -100, -44, 125, -67, -78, -14, -107, 99, -114, -62, -58, 59, -16, -85, 34, 2, 25, 30, 17, -72, -48, 61, 18, -106, 74, -4, -122, -51, -64, 23, -41, 0, 98, 126, -122, -1, -10, 107, -86, -127, -124, 58, -85, -103, -111, 14, 43, 109, -90, 104, -53, -17, -66, 32, -21, 90, -72, -115, 115, 102, 42, 64, -48, -64, -94, -67, -12, 48, -79, -74, 16, -51, -58, 55, 23, 81, -104, -116, -23, -67, 44, 29, -107, 72, 26, 46, 93, 81, -40, 18, -11, -11, -14, -53, -106, -10, -96, -97, 52, 105, -7, 88, -106, -60, 65, 91, 3, -124, -50, -93, -84, 112, -123, 123, 23, -32, 15, 18, 1, 87, 52, -84, -125, -36, 117, 70, 40, -97, -118, -118, -11, -97, -74, -37, -3, -113, 10, -123, 50, -41, -35, 81, -45, -62, -41, 76, 15, -116, 48, -105, -127, 24, -122, 78, 127, 20, 19, 108, -44, -28, 76, -46, -33, 121, 125, 108, 11, 58, -109, 61, -12, 72, 43, 33, -14, -90, -26, -115, -123, -1, -44, -92, -39, -39, 20, 94, 0, 50, 90, 62, 28, 114, 15, 5, 57, 127, 42, -45, -87, -52, -27, -90, 99, -36, -125, 11, -109, 86, -63, 64, -30, 44, 0, -103, -40, -84, -20, -97, -70, -121, 15, 89, 1, -5, 97, -121, 8, -36, 85, -77, -57, 62, -64, -20, 70, -120, -45, 76, 24, 93, -116, -28, -31, -118, 43, 32, -29, 40, 97, -66, -24, 79, 65, -16, 39, 75, -79, -124, 55, -76, 72, -112, -72, 82, -43, -80, -36, 101, -66, 27, -126, 51, 5, -33, -57, -89, 76, 38, -87, -43, -101, -100, -46, -36, 99, 80, -51, -40, 13, 70, 97, -30, 127, -76, 105, 68, 68, -40, 35, -77, 9, 15, 59, 34, -85, -116, 35, 8, 100, -68, 19, 44, -25, -40, 57, 66, -60, 23, -48, 38, -62, 30, -30, -18, -4, -95, -67, 111, -90, 106, 26, 112, 119, -16, -6, -86, 22, -4, 68, 46, 117, -31, -10, -125, 39, 122, 123, 14, 122, 38, 19, 125, 81, -107, 100, 75, -97, 75, 108, 31, -100, 28, 45, -5, -106, -3, -3, -98, -104, 17, 18, -108, -24, -61, 102, -12, -23, -7, 37, 96, 19, 38, 91, 70, 20, 67, 37, 127, -37, 117, -30, -8, 123, 5, -115, -98, 37, 29, 20, 46, 7, 106, 30, 94, 17, -70, 2, 106, 57, 119, 78, 121, -84, -32, -127, 69, -124, 39, 24, 53, -96, 24, -126, -93, -34, -55, -95, -63, 121, 16, 96, 56, -59, -64, 124, 44, 63, -89, 87, -120, 116, -40, -6, 86, 99, 38, 22, 89, -33, -62, -113, -89, -120, 109, 6, -113, -13, -36, 60, -42, -86, -100, -85, -122, -21, -112, 36, -120, -125, -67, -8, 110, -26, 56, -71, -85, -88, 53, 7, -74, 12, 101, -4, -100, 4, 113, 23, -70, -107, -8, 98, -118, 97, 115, 76, 61, 40, -60, -112, -15, 73, -67, 96, 59, 110, 35, 56, 87, 14, 73, -49, -53, -50, -49, 93, -52, 40, 120, 56, -112, 94, -77, 82, 95, -127, -96, 0, 118, -121, 100, -79, 27, -1, -70, -89, 14, -87, 45, 108, -125, 50, 76, 54, 27, -6, 54, -97, 75, -30, -76, -66, 100, 17, -35, -50, -4, -25, 13, 113, -123, 113, 98, -28, 33, 91, 93, -54, 100, 109, -76, -50, 66, -113, 81, 48, -29, -90, -41, 75, -120, 95, 106, -79, 100, -80, 43, -22, -3, 51, -69, -114, -110, -18, -58, -87, 109, -49, 59, -109, 98, -54, 40, -106, 26, -26, 22, 50, -124, 62, 116, -111, 102, -26, -48, 103, 10, 108, 46, 22, 17, 11, 119, -8, 15, -123, 53, 80, 38, 66, -12, 64, 91, 23, -101, 111, -83, 110, 88, -41, 113, 124, 52, -83, -54, 82, 57, -60, 6, 79, -37, 76, -127, 127, 98, -47, 33, 127, 110, -46, -15, 119, 86, -81, -54, -13, 35, 81, 80, 9, -12, 80, 38, 3, 113, 103, 56, -15, 24, -30, 6, -74, 63, 98, 35, 72, -36, 78, 78, -47, -85, 87, -78, 83, -19, 27, -118, -105, 51, -5, 18, 53, -24, -126, -111, -59, -15, 36, -93, 22, 4, 108, -125, -118, -7, -34, 123, 79, -89, -125, -25, -50, 124, 98, -104, 43, -59, -53, -93, 11, 92, 91, -6, -121, 77, 116, -33, -65, 107, 33, -60, -65, 34, -128, 33, -71, 115, 66, 109, -121, 36, -39, 72, 104, -111, 21, 109, 20, -55, -98, -23, 87, -115, -5, 58, 69, -70, 64, 103, 65, -50, 111, 103, 88, 125, 54, -67, -56, -88, -124, -55, 117, 83, -61, 28, 45, 114, -6, -73, 109, -61, 70, 45, 5, -100, -7, 112, -48, 97, 111, 32, -51, -89, 33, 124, -106, -24, -25, 71, -80, 110, 55, -65, 21, 104, 44, -44, 52, -56, 80, -13, -116, -94, 45, -113, 25, 93, 116, -85, 16, -107, -82, 18, -46, -117, -107, -41, 115, 110, 24, -58, -61, 50, -5, 75, -46, -89, 8, -93, 47, -123, 121, 69, -54, -122, -88, 3, 26, -23, -14, 61, 121, 24, -74, -10, 84, -60, -126, 59, 0, -47, -20, 90, 115, 123, 11, 88, -45, 86, 14, -70, 108, 90, -32, 24, -32, 121, 105, 112, -3, -93, 78, -23, 110, 20, -93, -96, 14, -68, -62, 66, -4, -57, 23, 105, -64, -98, -56, 67, -29, 21, 60, 120, 37, -72, 24, 80, -80, -80, 28, 78, -31, -34, -59, -69, 4, -112, -110, -93, -46, 66, -1, 30, 6, 51, 38, -13, 49, 93, -39, 79, 45, 77, -38, -4, 30, -83, 21, 104, -50, -51, 13, 67, 47, 65, 87, 91, 0, -123, -121, 101, -70, 108, -65, -58, -67, -36, 47, 113, -77, -49, 83, 18, 53, 39, 61, -16, -123, 27, 4, 11, -10, -66, 11, 106, 73, -55, -120, 69, -87, -16, -112, 13, -36, -95, 12, -73, -66, -59, -126, -17, 118, 49, -48, 48, 87, -18, -121, 124, -44, 19, -44, -33, 41, 10, -60, 112, -32, -121, 95, 99, 60, 83, 15, -21, -21, 88, 83, 28, -38, 74, -69, -110, 113, -74, 70, -22, -99, 87, -34, -67, 126, 123, -120, 116, 123, -78, -92, 15, -126, -37, -64, 99, 43, 106, 15, 42, 10, 6, 36, 61, 52, 81, -23, 80, 27, -13, -102, -29, 5, -128, -32, -42, -73, -33, -123, 74, 20, 125, 30, 93, -22, -113, 78, 119, -91, -38, 35, 4, -92, -46, -55, 60, -23, -7, 10, -29, 57, -60, -29, 107, -85, 47, -23, 7, 23, -18, 122, 37, 94, -80, -82, 109, 108, 4, 29, -34, 48, -24, -74, 32, 61, -111, -5, 57, -113, 46, 22, 42, -92, 121, -58, -39, -122, -75, -13, -119, -9, 49, -115, 3, -19, -94, 93, 73, 16, -110, -26, 14, 104, 54, -28, -24, -112, -72, 71, 117, 11, -43, -110, 7, 82, 123, 0, 100, 28, -22, -120, -109, 73, 127, 100, 79, -126, -84, 60, -100, -63, -64, -16, -118, 58, 101, -35, 22, -99, 29, -88, 58, -111, 47, -20, -36, 68, 56, 99, 81, 69, -124, 27, -107, -125, -23, 41, -110, -98, 106, -31, 111, -2, -55, -46, -54, 10, 64, 34, -24, 7, -90, 125, -106, -28, -9, -107, -41, -16, -30, 92, 36, -44, 77, -3, 96, -35, 69, 2, -37, 50, 63, -53, -56, -103, 28, 71, -32, 126, -93, 79, -46, -81, -30, -54, 48, 5, 17, 127, -14, 94, 98, -49, 51, 51, 29, -114, 67, 104, 34, 20, -82, 39, -111, 96, -21, 110, -4, 127, 109, -82, -66, 98, -18, -27, -36, -101, 120, -58, 68, 112, -72, -94, -15, 56, 104, -7, 116, 93, 101, -25, 123, 57, -103, 80, -124, 81, 117, -34, 6, -114, -10, 45, 13, -100, -87, 41, -32, -106, 82, -33, -76, -72, 109, 125, 52, 55, -3, 89, -28, -45, -45, 95, 62, -58, -62, 52, 67, -100, -99, -56, 108, -42, 116, 81, 29, 30, -17, 126, 126, -94, 28, 57, 91, -73, 82, -92, 55, 119, 45, -47, 77, 73, 22, -37, -24, -104, -22, 66, 117, 43, -61, 26, 17, 60, -103, -78, -75, 19, 54, -40, 62, -73, 35, -120, 26, 86, 32, 35, -94, -108, 126, -81, -118, -55, -83, 60, 81, -10, 52, -87, 69, 66, 95, -125, 9, 94, -31, 121, -106, 37, -48, -115, 108, -111, -1, -42, -85, 13, -55, 81, 97, -47, -38, 78, -14, 14, -43, 38, -69, 27, -108, 106, -60, 77, 96, -70, 51, -5, -94, -58, -45, 71, 24, -60, -20, -33, -37, -100, -88, 22, 84, 33, 88, -2, 92, -36, -8, 17, 69, 40, 117, 104, -47, 112, -6, 32, 52, -107, -70, -18, -111, -10, -19, -116, 8, 43, -52, 40, -86, -86, -88, -101, 11, 74, -81, 14, -42, 100, -82, -58, 34, -127, -43, 80, 122, -85, -97, 94, 109, 40, 103, 35, -46, 61, 91, -59, 24, -81, 47, -96, 121, 115, 56, 29, -127, 43, -113, 5, 97, 76, -58, -63, 6, 17, -76, 108, -92, -83, -83, 2, 54, -122, 101, -125, 3, 85, 72, 105, 74, -13, -45, -109, -74, 49, -11, 114, 103, 122, -45, -104, 95, -112, -96, 93, -11, -118, 127, -98, -7, -29, 67, -50, -25, 73, -16, 0, -67, 84, -50, -73, -50, -114, -36, -53, -127, -5, -44, -27, -117, 34, -96, -50, 90, -40, 107, 14, 86, -76, 94, 50, -20, -88, -53, -124, 34, 32, 27, 84, 9, -53, 24, 71, 53, 98, -99, -17, -116, -39, 15, -36, -64, -90, -36, 53, -78, 31, -122, -105, -29, -107, 8, -8, 29, 19, 12, 3, -79, 23, -82, 45, -127, 67, 104, -108, -78, 88, -50, 30, -94, 91, -108, 92, 66, -4, 17, -46, -7, -30, 84, -49, 104, 75, 52, 99, -91, 13, -61, -80, -35, -21, 15, 76, -86, 102, 53, 40, 48, 74, -39, 109, 1, -45, -13, 102, 72, -122, -88, 9, 30, -79, -102, 96, 54, 52, -52, 6, 80, -25, -25, -99, 0, -78, -62, -93, -36, -48, 54, 26, -79, 39, -98, -75, 106, 92, -66, 64, 9, -119, -107, 89, -80, -52, 55, -44, -55, -44, 93, 31, 71, 55, 44, 22, -7, 9, 108, -75, -61, 57, -95, -24, 95, -11, -45, -110, 36, 108, 17, 79, -63, -108, 87, 107, 69, 94, -124, 49, 39, 83, 70, 51, 12, -6, 24, 123, -38, 61, 78, -83, -96, -52, -29, 23, -44, 90, 65, -88, -3, -90, -37, -19, 47, 29, -59, -117, -14, -6, -37, 76, 0, 76, -104, 91, -51, 63, 26, -19, 127, -32, 30, -101, 87, -25, -85, -95, 68, 26, 89, -14, 40, 30, -16, -21, 40, -127, 11, -25, 37, -111, -43, -95, -113, 60, 95, 99, -79, -127, -80, -68, -57, 7, -104, 88, -45, 58, -4, 9, 35, 1, 6, 82, 35, 73, -110, -104, 108, 33, 118, -20, -8, 113, -62, -107, -15, -75, 93, -99, -27, -63, 125, -18, 72, -1, -117, -66, 61, -4, -37, -77, -123, -71, 20, 37, 53, 74, -80, 106, 103, -7, -38, -105, -82, 78, -92, 116, -110, 19, 63, 123, -2, 67, 41, -55, -115, 43, 24, -77, -26, -9, 105, 101, -50, -15, -42, 70, 12, 57, -95, 50, -54, -102, 51, 127, 29, -80, 81, -31, -126, -58, 12, 123, 80, -74, 14, -111, 15, 40, -126, 103, -96, -43, -5, 58, 31, 50, -2, -116, 62, 21, 14, -8, -73, 94, 59, 19, -10, -113, 118, 75, -99, 53, 91, -128, 119, 122, -43, -5, 33, 20, 79, -6, 70, 121, 105, 78, 66, 40, -45, -67, -24, -90, 76, -30, -119, 102, -98, 51, -51, -92, -84, 84, -7, 47, 73, 65, -107, 76, 30, 87, -52, -82, -30, -111, -104, -29, -4, -75, 40, 66, 21, 9, -113, -96, 112, -80, 7, -92, 27, 30, -80, 108, 71, -118, -123, 2, 15, 49, -58, 42, 91, 35, 73, -92, 110, 94, -121, -28, -110, 79, 56, 31, 63, 39, -90, -2, -121, 11, 59, -8, -70, -28, 57, 30, 24, -98, 64, -51, 55, 96, -9, 83, -96, -54, 4, 126, -51, -23, -63, -78, -93, -98, -118, -94, -42, -45, -47, -37, -116, -63, 84, 123, 85, -72, -13, 118, 119, 100, 43, 92, 93, 63, 7, -16, 98, -54, 105, -50, 57, 117, -86, 14, 47, -128, 47, -27, -11, 19, 114, 74, -6, -21, 101, 2, 25, -11, 17, -118, -75, -107, 127, -115, -69, -1, 89, -24, -22, -97, -99, 25, -110, -84, -123, 47, 119, -39, 86, 43, 29, -14, -41, -72, -117, -81, 83, 85, -63, 46, 85, 126, 87, -70, -116, -62, -83, 108, 42, 124, -20, -39, -84, 7, -100, 32, 109, 35, 16, -13, 84, 52, -35, -46, 35, -39, -54, -106, 55, 38, -122, -56, -103, 49, 76, -96, -16, -82, 85, 92, -34, 32, -36, 5, 57, 92, 51, -99, 126, 58, -61, 123, -98, -30, -115, 112, 123, -82, -123, -65, 33, 76, 85, 5, -1, -98, 23, 104, 6, 25, -61, 18, 37, -22, 11, 126, -27, 76, 91, -47, 57, -8, 68, -40, 34, -51, 123, -123, -16, 94, 27, -94, -118, 114, 41, 64, -4, -48, 120, 43, -72, 26, -91, -6, -15, 43, -29, 55, -87, 21, -83, -58, 117, 50, 37, 99, 121, 30, -91, -69, 112, -77, -65, -45, -85, 85, -16, 73, 98, -8, -49, -128, 98, 93, 62, -40, -108, -94, -16, -36, -69, -67, 59, 103, 32, -100, -30, 102, -106, -45, -73, 104, 100, 67, 54, -92, 21, -122, -126, -109, -32, 96, -67, -24, -44, 60, 63, -51, -126, 74, 33, -99, 80, -105, 26, 18, -19, -105, -100, 80, -33, -104, 123, -60, 7, -46, 126, -42, -84, -27, -46, -60, 99, 78, -24, -103, -52, 12, -69, 69, 49, -109, -78, -9, 44, 34, 110, -10, 81, -59, -39, -111, 74, 15, 83, -48, 44, 27, -120, 31, 25, 28, 76, 51, -74, 22, 106, -40, -103, 0, -101, 18, 76, 47, -27, -110, 51, -95, 64, 117, -31, -75, 59, 65, -116, 67, 95, -80, -76, 78, -83, 16, -107, -38, -51, 45, 22, 73, -68, 27, 20, -70, -113, 40, -93, 83, -20, 17, 117, 7, -93, 87, 60, 4, -107, 3, 50, -27, 16, 83, -64, 28, 125, -76, 114, 70, 108, -115, 120, 93, 26, -92, -109, -57, 102, 95, 52, 72, 126, -38, -74, -7, -121, 35, 100, -44, -71, 118, -72, 108, -49, -68, -74, 64, 49, 29, 60, 88, 27, 123, -115, -105, 77, 124, -106, -57, -100, -99, -15, 92, -72, -55, -54, 51, -82, 18, 119, 52, -3, -24, -35, 114, 36, -59, 56, 50, -118, -5, -101, 108, 69, 53, -40, -103, 22, -127, -65, -100, 34, -100, 92, -49, 4, -124, 119, 79, 46, 95, -77, -49, -55, -95, -7, 112, -56, -6, 125, 4, 48, 91, -28, 12, 117, 40, -42, -105, -38, -82, -62, -78, -38, -70, 104, 124, 29, 54, -86, 83, -104, 53, 127, 17, -70, -63, -89, -125, 55, -45, 46, 84, -98, 103, 50, 45, 115, 117, 118, -81, 79, 14, -54, -63, -124, -92, -78, -40, 102, -23, -114, 122, -10, 118, -36, 56, -121, -43, 100, 70, 68, -14, 105, -110, -67, 38, -20, -70, -124, 60, -61, 10, 18, 125, -66, -114, -67, 84, 81, 53, 88, 9, 63, 59, -56, -84, -4, 111, 8, 91, 62, -48, 26, -53, 24, 16, -18, 79, -22, 33, 79, 0, -115, 37, -58, -35, 71, 38, 69, -4, 58, -9, -20, 46, -114, 109, 79, 116, 103, 3, -107, 69, -100, 19, 96, 42, 96, 70, 5, 1, -110, 85, -105, -94, 8, 77, -100, -91, -113, -73, -63, 79, 113, -108, -54, -45, 53, 76, -108, -21, -57, 21, -102, 62, 63, 42, -42, 34, -88, 125, 45, 20, -86, -77, 90, -24, -62, 13, -80, 22, 76, 91, 91, -124, -94, 56, 115, -42, -16, -102, -11, -116, 111, 17, -2, -126, -43, -79, -41, -106, 58, -28, -14, -50, 124, 26, -75, 97, 56, -53, 29, -68, -96, -11, -15, -83, 9, 13, -68, -14, -53, -49, 46, -112, -94, -25, -62, 23, 73, 82, 85, -4, -101, -98, 57, 7, -49, 63, 70, -74, 69, -108, -37, 33, 1, 18, -116, -12, 24, -98, 64, 62, -13, 34, 49, 26, -32, 20, 92, -53, -63, 7, 47, 99, 1, 97, -25, -68, 31, -101, -27, -107, 22, -89, 46, 7, 84, 55, -37, 80, -53, 7, -97, -97, -26, 53, 104, 100, 67, 2, 7, -99, 69, 53, -3, -87, -40, -26, 106, -31, -73, 62, 95, 7, -35, 117, 56, -52, 51, -74, -93, 2, -62, 127, -56, 98, -53, 105, 41, 46, -7, 29, 52, 113, -127, -2, 101, 111, 48, 7, -106, -96, -7, -22, 14, -101, -128, -61, 121, 32, -66, 42, 13, -33, -91, 114, -95, -71, 58, -70, 117, 4, -99, 57, -35, 94, 43, -29, 109, 41, -21, -48, -126, -109, 96, 44, 55, 68, 19, -68, -24, -126, 57, -28, 79, -46, -105, -102, -36, 45, 84, 12, 33, 122, -46, 80, 20, -72, -102, 56, -7, 44, -39, 40, -85, -54, 68, -127, -98, -29, -90, -121, 13, -25, 86, 3, 61, -80, 79, 19, -31, -59, -125, 5, 24, 10, -123, 9, 71, 17, -107, -78, -10, -82, 5, 3, 87, 91, 44, 112, -46, -69, 28, 20, -44, -121, -30, 123, 121, -88, 83, 79, -90, 77, -95, 110, -49, -50, 110, 7, -15, -1, -11, 120, 38, 5, -88, -56, 101, 3, -121, 6, -9, 48, -53, -11, -86, -19, 5, 63, 39, 86, 122, -99, 105, -120, -81, 117, -44, 13, 126, -19, 96, -38, 20, 42, 124, -41, -4, 15, 13, 45, 34, -62, 95, 115, -60, 125, 31, 102, -58, -24, 114, 24, 35, 56, -31, -21, -42, 85, -78, -37, 57, -118, -7, 103, 59, -83, -7, 61, -58, -116, 122, -128, -54, -96, 49, 72, 89, -30, 55, 89, -110, -111, -6, -11, -94, -106, 45, -29, 13, 99, -99, -2, -106, 74, 58, 99, 54, 4, -13, -65, -104, -116, -36, 111, -12, -121, -122, 70, 124, 28, 46, -39, -58, 115, -93, -55, -13, -24, 50, 62, -61, -14, 48, 102, 30, 76, 76, 106, 42, -68, 123, -57, 8, -119, 16, -78, 19, -53, 23, 64, -54, -30, 124, -30, 99, -44, 20, 19, 6, -55, 6, 61, -46, -52, 74, 93, -7, 104, 127, -31, 98, 110, 45, 16, -111, -21, -59, -124, 83, 32, -104, -32, 77, -44, 62, -64, 93, -81, 108, 89, 29, 24, 70, 89, 78, 51, -60, 58, 85, 83, -128, 109, 96, -124, 83, 33, 51, 63, -28, 40, -31, -27, -37, 59, -43, -43, -20, -112, -91, 120, -106, 44, 37, 41, 45, -53, -36, -84, -125, -46, 124, 124, -50, 99, 113, -47, 74, 125, -27, 106, 90, -15, 119, -96, -107, -58, 92, 64, -125, 0, -44, -52, -121, -87, 12, 81, 110, -46, -118, -94, -34, -47, -12, -103, 50, 26, 2, 106, -21, -7, -4, 111, -111, 78, 10, 118, 97, -100, -71, 14, 35, 62, 80, -117, 100, 47, 66, -30, -63, 32, 27, -117, -60, 70, -7, 66, 127, 27, 22, 10, 4, 75, 31, -108, 56, 117, 50, -13, -66, 127, 21, -27, 21, 16, -125, 104, -115, -127, -57, -6, 46, -45, -110, -38, -39, 71, 111, -57, 68, -118, -86, 72, 123, 122, -96, 47, -14, -27, 44, 84, -47, 20, -54, -80, -48, 27, -6, 125, 127, 61, 82, 87, -38, 76, -73, -98, 28, 95, -71, 101, -39, -55, 121, 68, 24, 84, -77, -93, -93, -119, 98, 22, 61, -6, 121, 101, -55, -49, -75, 62, -80, -106, -58, 68, 8, 15, -2, 31, -8, 100, -82, -22, 70, -109, -11, 40, 2, -121, 24, -23, -55, 73, 74, -36, 53, 27, -101, 75, -7, 31, -2, 76, 26, -12, -17, -88, 57, -112, -34, 32, -42, 67, 86, 54, -65, -3, 55, -94, -110, -110, 116, -112, 11, -50, 50, 54, -99, 103, -11, -20, -126, 103, 10, 86, 109, -64, -127, 61, 67, 99, 104, -18, -66, 80, 114, 51, -68, -92, -128, -55, 86, 45, 78, -70, -10, -90, 37, 126, -50, -104, 35, -87, -32, 110, -116, 73, -7, -89, 25, 59, 91, 92, -81, 116, 39, -119, -110, -112, 125, 88, -100, -122, -66, -60, -34, 63, 99, -68, -8, -61, 38, -21, 34, 30, -89, -50, -118, 33, -32, 95, 25, -32, 5, 46, 80, 6, 2, 89, -25, -14, 55, 104, 82, -34, 21, -71, 108, 111, -35, -81, -39, 9, 11, 35, -122, 51, 58, 103, 97, -79, 59, -128, 41, 70, -85, -19, -127, 45, 56, 63, -6, 77, 54, -66, 32, -9, -77, -117, -12, 103, 86, -4, 80, -70, -6, -83, 35, 114, -14, -4, 112, -118, -55, 63, -32, -105, 80, 107, 120, 115, 106, -64, 84, -94, -4, -26, 47, -39, 64, -77, 114, -65, 105, 37, -95, -44, -11, -33, 26, -126, -14, 63, -13, 120, -96, -56, 73, -79, 101, 47, 33, 115, 68, -21, 89, -99, 48, 60, 57, -46, 45, 60, 1, -112, 59, -4, 50, -121, 34, -33, -17, -74, 106, 102, -107, 11, 119, 49, -78, -1, 112, -18, 117, 40, -72, -18, -110, 66, -91, 35, 79, -112, -78, 31, 40, -73, -61, -61, 58, 89, -51, -105, -32, 114, -110, 78, -55, -24, -106, -40, 52, 94, 83, -60, -7, -22, -4, 13, -37, 42, -98, -30, 25, -81, 6, 83, -124, 38, 78, 68, 35, 118, -47, 104, -72, -82, -44, -1, 42, 121, -92, -113, -101, 114, 99, -105, -37, 1, -54, 91, 91, 1, -86, 68, 126, -50, -67, 127, 76, 106, -127, 58, 77, -110, -85, 105, -20, 80, -93, 113, -45, 98, -57, -100, 82, 115, -45, -34, -106, -69, -82, -15, -30, -15, -68, -103, -66, 51, -109, 21, 124, -115, -64, -56, -74, 68, -109, -111, 83, 2, -23, 11, 84, -66, 31, 52, -43, 70, 13, 104, -59, 80, 31, -111, -93, -104, -70, -58, -105, -106, -46, -54, -88, -99, -70, 49, 66, 80, 35, -94, -78, 42, -20, 42, 39, -44, -18, 18, 23, -41, -53, -46, 76, 59, -37, 26, -42, 81, -87, 96, -9, 88, -95, 64, 92, 8, -60, 79, -125, -5, -26, -36, -45, -62, -112, 30, 96, -27, 107, -82, 9, -51, -114, 37, 75, -8, -125, 111, 94, 39, 94, -113, -47, -33, -115, 16, -110, -13, 117, 40, 21, 72, 34, -116, 110, -85, -115, 99, -21, -120, -76, 90, -117, -6, 43, 116, 74, 82, 30, -15, 120, 55, -79, 98, -123, 124, 86, 108, 61, 122, 48, -46, 100, 96, 26, -95, -67, 104, 58, 34, 10, 25, 125, 104, -104, 118, -15, 22, -97, -68, -87, 89, 42, 64, -1, -102, 69, -53, -59, 48, 59, 54, 108, 39, 30, -18, -124, -43, -82, 31, -82, -73, 97, 97, -40, 61, -124, -6, -124, -32, 109, -73, -104, 18, -83, -102, 108, -106, -93, 43, 115, -1, 75, -31, -117, 20, 9, -53, 71, 73, -54, -107, -19, -12, 124, 118, 81, 98, 5, 36, -39, 77, 57, 81, -127, -53, -49, 58, 30, -62, -5, 22, 109, -111, -12, 123, -66, 82, -102, 51, -43, -73, 97, 120, -83, -19, -107, -83, 18, -11, 1, -77, 61, -79, -36, 54, -26, 111, -5, 93, -76, -114, 31, -53, -91, 34, 22, 111, -54, 43, -97, -123, 122, 121, -15, -63, -59, 69, -16, -85, 119, -80, -128, 48, 120, -121, 37, -62, -74, -105, 31, 94, 125, 31, -78, 92, 51, 35, 36, 101, -99, 55, 62, 91, 92, -39, 107, 7, 5, -118, -33, -91, 43, -18, -105, 115, -30, 65, -47, 115, -54, 101, 98, 30, -126, 32, 0, 117, 1, 24, 126, -4, 126, -68, -52, -7, 2, -2, 118, 92, -12, -100, -94, -114, -42, 19, 5, 90, 80, 110, -37, 58, 64, 86, 9, -26, -25, -7, -73, -114, -54, 6, -49, -37, 74, -44, 5, 98, 48, 29, -83, -108, -38, 75, 71, -33, -103, 106, 94, -128, -87, -75, -64, -77, 54, -68, 5, 8, 22, 11, -44, 117, -108, -99, -93, 22, 91, -29, 78, 39, -90, -1, 54, -22, 34, 67, -77, 89, 70, 3, -122, 65, -50, -123, -97, -47, 93, -51, -110, 84, 110, -86, 127, 6, -46, 63, -64, -88, -61, -122, 112, 108, 95, 11, -99, 99, 56, 104, -92, 55, 35, 8, -33, -14, -10, -21, 88, 69, 51, 82, 98, -82, -105, -74, -112, -102, -89, -31, -101, 83, 115, 91, 35, -60, 71, -17, -106, 29, 93, 80, -94, -98, -99, 58, 89, -109, -21, -22, -85, 27, 74, -47, -63, 9, 22, 124, -44, -1, 15, 42, 49, 87, 118, -62, 18, 36, 69, 77, -96, 63, -101, 68, 10, -73, 44, 24, -118, 29, -124, 117, 3, 87, 26, -79, -119, 12, -104, -114, 29, 31, 49, -111, 36, 64, -85, -111, 18, 119, -77, 28, 90, -83, 38, -106, 6, -41, -45, 120, -126, 54, -74, 80, 3, 73, 104, -32, 46, -22, -40, -26, -62, -30, 123, -91, 93, -95, -9, -125, 2, -82, 27, -38, -31, 82, -124, -62, -88, -22, 42, -114, -11, 52, 80, -33, -19, 107, -118, 11, -38, -118, 101, 82, -34, 24, -94, -67, 91, 33, -122, -99, 89, 71, -98, 92, 100, -19, -44, 1, -110, -83, 22, 126, -123, 108, -113, 34, -108, -20, 123, -127, 29, 85, 123, -2, 79, 45, -76, -18, -107, -49, -79, -68, 55, -112, -90, 98, 33, -123, 16, 69, 78, -26, 7, -55, 56, 69, -65, -126, -51, 117, 91, 31, 0, 10, 9, -29, -74, -34, 84, -120, 42, 87, 79, 0, 110, -80, 3, -81, 29, 33, 104, -121, -10, 75, 8, -27, -77, -121, -50, 56, 26, -27, -12, 16, 111, 63, 36, 5, -12, -108, 81, 109, -69, 82, 91, -70, -108, -54, 111, -88, -111, -40, -125, -97, -29, 11, 67, -58, -45, 4, 120, 36, 20, 114, -28, 106, -87, 73, -115, 126, 51, 42, 23, -38, -126, -71, 105, -60, 74, 37, 125, 106, -102, -107, 109, 114, -76, 63, 95, 15, 63, 85, 16, -88, -65, -128, 117, 32, 101, -80, 33, -93, -104, 67, -62, 7, -113, 117, 97, 91, 52, -37, 107, -74, -46, 115, -1, 70, -78, -19, 20, -75, -114, -80, -25, 63, 99, -42, 96, -88, 50, -36, -61, 53, 24, 120, -70, -23, 42, -5, 59, 99, -103, -72, -106, 53, 107, 117, 4, -48, -70, -30, -69, -61, -98, -66, 21, -39, -20, -119, -89, 1, 45, 98, 62, -27, 40, 60, 63, 78, 1, -47, 42, -43, -31, 38, 94, 126, -27, 53, 51, -8, -104, -86, 107, 109, 77, 1, 122, -22, 96, -53, 31, -88, -103, 45, -39, 10, 44, 90, -76, 52, 2, 10, -59, -5, 40, 0, -85, 74, -21, 112, -36, 106, 47, 34, 1, -96, -7, 96, 42, -110, -11, -128, 80, 51, -2, 50, -71, 27, -23, 116, -109, 8, 5, -70, 22, 33, 102, 17, 99, 50, -15, 127, -21, 37, 4, 19, 96, 87, 39, 55, -73, -102, 71, 7, -3, 11, 59, 68, -57, 50, 2, -33, 20, 73, 14, 70, -56, 99, -48, -26, 3, -110, 67, -27, 27, -99, -13, 106, -38, 123, 24, -71, -87, -42, -52, 58, -45, -97, -70, 123, 108, 102, -42, -107, 70, -44, -126, 121, -59, 58, 59, 56, -80, 56, 82, -86, -27, 72, 78, -11, -74, -39, 122, -16, -79, 42, -27, -86, 58, 25, 67, -61, 54, 22, -121, -38, -37, -44, -112, 22, 58, -36, -94, 88, 17, 12, -73, 31, 68, -80, -43, -116, -10, -13, -121, -12, -58, 24, 104, 60, 58, 18, -43, -25, -28, 65, -117, -42, -95, 30, 75, -116, 22, 24, 106, -100, 102, 99, -26, -2, -127, -85, -74, -108, 101, -79, -2, 112, 88, 124, -48, 42, 3, 88, -111, 25, 53, -31, -78, -107, 21, -33, -76, -3, 123, -122, -120, -107, -70, -37, -17, -108, -62, -14, -74, 17, -61, 62, 67, 88, -126, -82, -8, 64, -55, 93, -116, 2, 9, 120, 119, 73, 63, 78, 62, 80, 16, -61, 38, -118, -8, 63, -80, 73, -48, 98, -103, 23, -81, 74, 80, 6, -37, -38, 65, -90, -110, 60, -93, 28, 78, 64, 104, 96, -66, 112, 28, 92, 112, -19, -105, 106, 44, -11, -118, -111, -102, -63, 40, -27, -108, 40, 48, 34, -65, -109, -10, -79, -64, -24, -11, 33, 78, -104, -42, -40, 35, -43, -8, 114, 109, 127, -125, 55, -81, -78, 62, -102, -96, 7, -31, -84, 122, -43, 92, -53, -120, 72, 6, -59, 52, -7, 113, 21, -48, -58, -112, 0, 102, -28, -122, -12, 67, -74, 16, 12, -109, 59, 96, 111, 34, 81, -22, 126, -29, -19, 44, 41, -42, -91, 121, 55, -101, 60, -46, -110, 80, 80, -36, -4, -3, 121, 30, -80, -120, 62, 22, 61, -12, -97, 99, 1, 66, 63, -36, 115, -66, 85, 14, 53, 23, -103, -126, 35, -83, 46, -21, 102, 54, -116, 21, -41, -17, 102, 112, 100, 64, 57, -104, -5, -106, -7, 8, 38, -86, -82, 55, 119, -96, -27, 14, -122, -115, -54, 93, 46, -57, -115, -61, 35, 10, -4, 13, -115, 71, 56, -90, 108, -38, 111, -57, 36, -89, 100, -78, -12, 49, -113, -33, -45, -69, -119, -92, -52, -47, 44, 29, -106, 6, -28, -27, 71, 56, -23, 106, 37, 106, -32, -111, 67, -75, -24, 45, -24, -68, 1, -113, -109, 16, 121, 11, -106, -48, -25, 0, 47, 70, 50, -28, -32, -12, -86, -61, -125, -18, 39, 48, -101, -123, -116, -77, -72, 126, 8, -69, 20, 88, -35, 18, -53, -85, 113, 22, -71, 113, 9, 9, 77, 52, 18, 74, 24, -80, 76, 60, -69, 41, 91, -76, -104, -119, 82, -68, 85, 115, 5, -31, 83, -27, 37, -48, -31, -78, -11, 74, -79, -109, 8, 2, -4, 56, -80, -12, 44, -125, -121, 78, 58, -99, -45, 65, 10, 19, 54, 2, -27, 27, 110, 20, -121, 114, -36, 119, 29, -100, -32, 1, -34, -120, -93, 14, -27, 91, 22, 28, -78, -124, 10, 85, -9, 123, -90, 102, -15, -24, -73, -72, -12, 113, -30, 12, 43, 1, -33, -9, 76, -106, 14, 5, -55, -61, 45, -85, -126, -56, 13, 28, -72, -13, -43, 112, -90, -81, -95, 127, 70, 43, 33, 121, 61, -125, -88, 102, -109, -52, -70, 6, -114, -3, 74, -48, 88, -77, 102, 103, -63, -27, 58, 116, 122, 68, 5, 113, -15, -17, -99, 80, -69, -123, -118, -29, -32, 95, 32, -13, 69, -79, -86, 63, -114, 8, -98, -94, -93, -8, 38, -19, -78, 122, -121, -125, 11, -24, -5, 14, -81, -100, 115, 34, -14, -45, 113, -43, 87, 92, -116, 79, 126, -127, 31, -101, 100, 6, 82, 66, -24, -97, -119, 92, 98, 8, 112, 14, -34, 27, 58, 55, -21, 104, 54, 107, -89, -45, 15, 42, -124, 60, 8, 45, 94, -17, -103, 122, 60, -80, -103, 5, -48, -41, -71, -117, -108, 97, 67, 125, 52, 104, 5, 69, 6, 123, -38, -11, -9, 70, -11, -73, 10, 120, -110, 26, -94, 26, 66, 116, -58, -22, 2, 8, -1, -39, -95, 101, -105, -32, 101, 124, 96, 0, -2, -106, 25, 79, 23, 84, 118, -45, -67, 37, -91, 42, -80, -46, -71, 10, 74, 120, -124, 122, -99, -120, 79, 22, -125, -52, 56, -88, 61, -41, 33, 106, -106, 41, -64, -92, 31, -52, 117, 103, -28, 29, 8, 115, -81, 112, -1, 87, 69, 109, -41, 67, 68, -17, -127, 100, -70, -90, -26, -36, 43, -29, -90, 127, 13, -108, -87, -49, 56, -41, 31, 110, -85, 74, -63, 52, -108, 93, 59, -1, -62, -101, 95, 79, -58, -121, -58, 109, -39, 56, -35, 107, 119, -2, 118, -60, 2, -127, -127, 9, -10, -84, 49, -109, -15, -104, 0, -30, -128, -71, -2, 78, 56, -1, 102, -14, 77, 82, 35, 125, -66, -81, 45, -117, -105, -101, 50, -76, -24, -81, 75, -96, -78, 73, -71, 80, -94, 55, -42, -72, -78, 47, -48, -39, 36, 97, 44, 116, -29, -7, -90, 126, 54, -63, 82, 11, -53, 4, -108, -42, 0, 91, 81, -71, 93, 12, -27, -108, -34, -57, 61, 64, 57, -7, -11, 35, 37, 39, -105, -60, -62, -108, 105, -99, -52, -89, 105, -24, -110, -73, 61, -99, 38, -7, 74, -83, 103, -101, -14, 20, 98, 68, -47, -30, 84, -43, -37, -24, -104, -103, 61, -82, 4, 118, -68, -14, -109, -51, 10, 0, 65, 37, 12, -103, -80, -111, 26, -66, 9, 21, 125, -16, 127, 22, -99, 58, 118, 89, -15, 105, 107, 68, -37, -58, 4, -14, 122, 120, 6, -62, -12, -103, -52, -91, 59, 67, -86, 56, 29, 52, -119, -112, -121, -26, 87, -107, 67, -126, 55, -57, 43, -1, -85, 114, 116, 45, -109, -63, 89, 61, -24, -33, -5, 12, 121, -126, 13, 12, -16, -127, -105, 101, 83, 85, 37, -50, -91, 26, 74, -118, 26, -93, 105, -106, -27, -123, 121, 49, -116, 113, -100, -14, -30, 71, 0, 85, -16, 42, -73, 6, -120, 119, 86, 6, 104, -79, 11, -25, 37, -19, 109, 55, 3, -68, 66, -71, 127, -113, 107, -89, -3, -60, 125, 28, 49, 105, -25, -31, -69, 123, -20, -71, 117, -18, -9, -91, 51, -5, 42, 29, -73, -69, -41, -14, 104, -109, 117, 23, -113, -69, 32, 25, -49, 8, -39, -49, -124, 5, 76, -53, -51, -106, -25, 106, 74, -18, 80, 51, -66, 33, -50, -120, -76, 94, 109, 47, 13, 123, 70, 85, 34, 25, -38, 18, 65, -46, -120, 0, 116, 72, -99, -10, -98, -23, -88, -5, 100, 68, -54, 113, 75, 21, 29, 54, -34, 98, 28, -99, 57, 58, 31, -85, 11, 56, -17, -36, 42, 19, -50, -123, 53, 29, -78, -108, 57, -42, -36, -95, 15, -78, 21, -14, -126, 49, 13, -37, -108, 52, 55, 75, 13, -116, -30, -64, -18, -47, -22, -40, 50, -78, 61, 41, -76, -63, 22, -69, -92, -126, -3, -93, -88, -88, 34, -108, 69, 102, 20, -74, 70, -1, -89, -25, -103, -33, -38, -65, 112, -74, -67, -94, -3, 58, 6, 44, -8, -112, -46, -77, 14, 25, -74, -64, -40, 67, 110, -30, -88, 127, -75, 81, -67, -56, 88, -14, -66, -81, 77, -52, -23, -16, 100, -17, -104, -81, -54, -80, 107, -79, 82, 89, -120, -22, 40, 16, -79, 83, 41, -121, -57, 53, -64, -19, -125, 16, -82, 49, -92, -119, -65, 62, -41, 75, 81, -43, 87, 59, -86, -95, 112, 66, -104, 32, 27, -125, 88, 20, 44, 109, -95, -85, 118, 85, 89, 50, 88, -107, -2, 4, -116, -46, 82, -67, -125, 89, -17, 11, 27, 14, -74, -115, -96, -83, 83, -112, 53, -88, -65, 89, -18, 43, -114, -85, -34, -47, 32, -78, -47, 13, 95, -64, -60, 4, -20, -50, 45, 126, -105, 43, 75, 117, 25, 97, -92, -99, -90, 60, -89, -83, 98, -81, -72, 75, -116, -10, -90, -88, -72, 94, -112, 28, 86, 13, -99, -46, -53, 82, 23, -95, 77, 38, 58, 101, 12, 112, 87, 112, -105, -13, -98, -93, 68, 70, 113, -54, 57, 50, -86, -7, -98, 78, 56, 0, 117, 37, 49, -51, 52, -63, -90, 54, 20, 121, 114, 16, -22, -50, 29, -55, -2, 95, -49, -124, 77, 67, 110, -45, 64, 89, 30, 115, -33, 33, 23, -7, 87, -114, 95, 67, -17, 63, 36, -98, 63, 7, -67, 7, -90, -1, -28, -100, 115, -40, 47, 73, -60, 100, -122, 55, 108, 76, -40, -108, -79, 4, -18, 64, 63, -49, -111, -77, -65, 76, -93, -56, -98, -56, 80, 45, 70, 57, 2, 111, 107, 34, 26, -82, -103, 36, 82, 64, -100, -53, 94, 24, 65, -1, -25, 26, -10, -32, -19, -32, -111, -113, 27, -106, 87, -116, -53, -94, 22, 22, -101, 19, 16, -108, -30, 7, -97, 82, -29, -34, -90, -78, 89, 70, 26, -25, 68, -79, -10, 28, -56, -114, -94, -69, -7, -44, -65, -41, 119, -107, -83, -64, -96, 76, -88, 50, -94, 64, 94, -45, -28, 32, -62, 83, -47, 17, 78, 44, -42, -90, -94, -66, -47, 78, -114, 121, 16, 81, -6, 32, 43, -19, -34, 59, 13, 4, -2, -44, 72, 28, -88, 19, 87, -96, -117, -9, -32, -58, -35, -47, 15, 32, -38, 42, -101, -79, 104, -7, -2, -83, -116, -50, 8, 43, 69, -11, 87, -61, -85, 91, 102, -51, 21, 36, -25, -33, -82, 19, 61, 61, 115, -109, -74, 52, 4, 110, -98, 122, 52, 32, -54, 115, 114, -23, 60, 63, -48, -124, 115, 126, -106, -4, -73, -105, 110, 76, 85, 104, -50, 92, 18, 42, -96, 81, 44, 41, -96, -74, -93, 49, -87, 70, -5, -66, -11, -18, -73, 22, -26, 13, -41, -2, -77, 103, 124, 54, -128, -7, 126, 89, 68, 8, 100, 127, 9, 53, -16, -14, -37, 16, 36, -62, 67, -120, -36, -38, -80, 30, 70, 31, -17, -95, -30, -108, -37, 96, 114, 44, 76, 121, -26, 82, -122, 11, -60, -93, -58, -80, 49, -103, -57, -116, -25, -35, -23, -72, -63, -77, 53, 21, -27, 53, 102, -84, -13, -87, -89, -20, -89, -79, 98, 41, -6, 40, -5, -102, -48, 35, -99, -97, 44, 5, 73, 38, 89, 65, -105, -73, -106, -125, -7, -36, 112, -16, 1, 123, 33, -17, -108, -40, -34, -74, 90, -9, 18, -61, 79, -48, 28, 98, -62, 100, -8, 8, 119, 87, -17, -54, -108, 121, -120, -110, 41, 72, 8, 60, -100, 113, 37, -99, 97, 120, -92, 75, -17, 57, 15, -53, -1, -34, -112, -71, 35, 108, -112, -35, 84, -5, 108, -116, -11, 25, -66, 8, -18, 69, -19, 67, 82, 24, 4, 83, 9, 55, 31, -2, -119, -57, -49, 54, -76, -65, -4, 86, 33, 104, 35, 55, 111, 122, -9, 63, 21, 111, 26, -59, 9, -92, 62, 39, 36, -55, -32, -29, -18, 35, 10, -44, -80, -89, 107, -43, -111, 111, 101, 125, 116, -3, 76, 46, -4, -48, -125, 92, -70, 101, -62, -6, -34, -41, 65, 125, 90, -58, 74, -46, 90, -81, -42, -91, 108, -64, -109, 74, -97, 105, -26, -67, -70, -57, -102, 98, 69, 125, -34, 31, -128, 86, -5, 84, 110, 110, 1, -93, 89, 115, 63, 70, -81, -126, -110, 21, -118, -126, -64, -103, 3, -110, 29, -50, -79, 9, 19, -60, -18, 108, -86, 55, 50, -23, -77, 44, 23, 30, 8, -17, -20, -92, 3, -42, -118, 55, 21, 53, 45, -46, -125, -7, 37, 15, -88, -24, -6, 115, -103, 83, 35, -98, 88, -76, -40, 25, -61, -17, 72, -14, -118, 118, -30, 63, 23, 90, 61, 111, 15, 65, 59, -46, 43, -2, 65, 45, 97, -88, -123, -125, -126, 62, -104, -83, -65, -56, 17, 70, 51, -14, -35, -2, -108, 66, -105, -126, -14, -24, 25, 106, -33, 34, -102, -99, 122, -52, -26, -122, 6, 43, -53, 22, 31, -52, -118, 15, -123, 88, -96, -33, 3, -123, -71, -75, 11, -57, -41, -69, 77, 57, -21, -22, 13, 38, -46, -45, 8, -59, 29, 35, -8, -42, -14, -36, -22, 5, -123, -84, -79, 69, -1, 4, -21, -34, 11, 64, -120, -71, 102, -4, -87, 19, -23, 127, -118, -28, 63, -124, -110, 124, 54, 125, 126, -118, 28, -60, 8, 30, 44, 71, -45, 25, 75, -17, 12, -125, 102, 88, 70, 109, -44, 69, -75, 24, 127, -47, -125, 48, 112, 68, -21, 88, -3, -101, 88, 27, -76, 121, -47, -89, 32, -47, 63, 65, -11, 74, 112, -100, 47, 77, -101, 41, -109, -108, 81, -96, 98, 24, 113, 67, -108, 107, 73, -88, -84, -69, 103, -98, -53, 46, 27, 68, 79, -74, 36, -33, 18, 0, 40, 31, -84, 0, 115, -122, -77, -122, -83, 108, -12, -25, 8, 108, -41, 34, 125, -70, -80, 27, -52, -73, -8, -25, -122, 41, -84, -120, 82, 119, -7, 110, -125, 8, 97, 113, 49, 89, 101, 12, 75, 13, 20, 96, -48, 2, -89, 41, 105, 72, -77, -114, -3, -86, 110, 54, -7, 64, 42, -38, -10, 92, 95, 88, 30, -35, 77, -85, 83, -111, 102, 25, -23, -52, -112, 82, 54, 102, -8, -93, 41, 48, 69, -3, 98, -87, 82, -81, 92, -22, -93, -1, 11, -78, -3, 53, -24, 127, -115, 78, -98, -108, 60, 82, -108, 42, 59, 59, 57, 97, -27, 51, 12, 93, 123, 109, -71, -46, 17, -72, -58, -52, 29, 44, -46, 78, 95, 29, -45, -91, 88, 42, 57, 5, -104, 125, 103, -123, -63, -101, 65, 97, -37, 14, 106, 84, 26, 92, 86, -43, -69, 89, 42, 118, 61, -58, -34, -42, 98, 77, 66, -17, 26, -48, 66, 7, 119, -13, -107, 122, -31, -85, -74, 119, -80, 76, 10, -67, 38, 102, -69, -79, 7, -21, -51, -78, 27, -42, 35, 107, -49, 61, -16, 126, 86, -89, -76, -105, -70, 95, 19, -92, -76, 86, -68, 86, -52, 66, 53, 102, 16, -6, -90, -84, 98, 100, -14, 73, -23, 100, 9, -57, 21, -120, -109, -15, -121, 33, 10, -25, -10, -42, -7, -14, -87, 69, 54, -35, 38, 51, -88, 88, 25, -115, -105, -8, 48, -62, 42, 7, 107, -101, 88, -36, 94, -25, -66, -42, -28, -17, 103, 125, -62, 46, 60, -10, -114, 63, -14, -57, 12, 85, -47, -127, 116, -11, 118, 16, 125, 111, -81, 78, -19, 43, 95, -35, -20, -98, -38, 48, 117, -123, 109, 77, -40, -77, 36, 5, 93, -50, -41, 49, -44, -50, 97, 113, 30, -71, 84, -50, -30, 70, -59, -56, 82, 121, -88, -20, 81, 61, -17, 31, 58, -56, 99, -15, -15, -128, -79, 89, 77, -125, 98, 53, 80, 87, 94, -80, 77, -28, 90, 124, -80, 56, 113, 35, 17, -102, 4, 121, -73, 13, 72, 43, -3, -44, 111, 124, -83, -5, 30, -72, -28, -22, -109, -50, 74, 7, 34, 15, 58, 11, 31, 74, -62, -84, 113, -62, -44, -62, 82, 114, -99, -111, 7, -32, 15, -88, -21, 88, 20, -28, 91, -125, -89, -33, -36, 0, 72, -29, -35, -94, -24, -70, 115, 114, 101, -86, 23, 64, 15, 45, -73, 19, -6, -102, 119, -60, -99, 78, -86, -55, -46, 48, 54, -70, 16, -76, 33, -91, -84, -49, 11, -86, 3, -119, 18, -9, -73, 75, -69, -49, 30, -58, -91, -124, 70, 109, 124, 108, 120, 50, 24, 113, -123, -31, -118, 6, -65, 7, 32, -101, 51, 23, 48, -26, 78, 74, 2, -12, -120, 124, -68, -106, -3, -10, -26, 3, -22, -65, -17, 23, 68, -47, -22, 23, -27, 54, 23, 78, -29, 102, -38, -110, 108, -13, -19, -70, -19, 81, 111, -38, 86, 71, -36, -60, -27, -11, 3, -114, 12, 111, 68, -82, -127, -111, 127, 69, -36, -106, 13, -81, 31, 100, 69, 89, -6, 61, -45, 46, 76, -55, -57, -44, -24, 80, 51, -96, -27, -119, -35, -87, 33, 106, -87, -123, 24, -60, -74, 61, 98, 35, -61, -35, 3, 68, 12, -113, -100, 83, 52, -77, 72, 51, -111, -47, 49, 123, -90, -76, 67, 28, 22, -25, -19, 100, 34, 106, -4, -93, 72, 92, -87, 30, 84, 90, 31, 21, 1, -84, -51, 19, 91, 32, -37, -35, -92, 123, -6, -54, -108, -88, 69, 54, 70, -58, 71, 124, 77, 24, -116, -100, 11, -61, -19, 16, -102, 12, -117, 40, -2, -22, -6, -3, -19, -3, 97, 24, 10, 30, 83, -126, 74, 86, 104, -19, -37, 29, -92, 44, 67, -32, 42, 85, 50, 114, 42, 68, -10, -18, 30, 76, 121, -104, -19, 15, -36, 14, -78, 63, 0, -113, 33, -14, -54, -34, 114, 27, 19, 112, 95, 59, -39, -58, 7, -34, -24, 29, -96, -123, -47, 78, -95, -79, -71, 27, -111, 16, -41, -77, 58, 33, -53, 58, -4, -98, 41, 61, -107, 48, -117, 2, -12, 107, -39, 37, -3, -32, -123, 62, -16, 123, -16, 47, -118, 115, 14, 68, -100, -75, 72, 76, -109, -78, -91, -12, -112, 59, 54, -37, -61, -65, -32, 42, -109, 10, 60, -93, -5, 95, 100, 39, 26, 25, -30, 22, 114, -85, 2, -89, 116, 3, -94, -85, -16, 27, -127, 0, -70, 47, -119, 117, -70, -20, 95, 122, 44, -114, 20, -79, -41, -20, -45, 53, 74, -38, -23, 46, 11, 122, -48, 31, -3, -63, 55, -72, -81, 30, 15, 35, -8, -96, 37, -83, 79, 70, -13, 48, 11, -82, -37, -62, 23, -70, 31, 78, -6, 23, 14, -15, 110, -47, -61, 123, 104, -56, 51, -20, 3, 36, 101, 11, 82, -92, -113, 122, 17, 65, 27, 53, -48, 66, 97, 123, 80, 23, 18, 79, -121, -128, -27, -8, 63, -43, -88, -26, -15, 98, 2, 126, 97, -123, -107, -96, 14, 118, 38, -30, 125, -86, 77, 20, -116, 123, 90, 3, -8, 80, -92, -35, -22, 57, -52, -6, -22, -118, -94, -59, 60, -19, 42, 102, -62, 93, 4, -81, -87, 39, 106, -43, 54, 26, 96, 70, 112, 89, -53, -83, -123, 47, -37, 44, 67, 84, 38, 62, 72, 52, -125, 1, 18, -72, 12, 77, 70, -90, 36, 14, -40, -70, -42, -69, 61, 119, -51, -94, 99, 53, -14, -16, -6, -9, -79, -22, -22, -36, 62, -48, 127, -64, 69, -24, -39, 15, 110, 52, -128, -114, -113, 31, -107, 19, 76, 52, -123, 59, -91, -47, -105, -58, 54, 100, -95, 69, 64, 67, 47, 77, -76, -52, -96, -46, 8, -79, 69, 79, 39, -59, 125, -59, -123, 53, -108, -3, 117, 3, 111, -24, 84, 58, 118, 4, 40, 7, -81, -13, -53, -94, -71, -24, 59, 36, -105, 27, 110, 0, -27, -93, 58, -84, 103, 35, 62, 12, 35, 40, -16, 71, 118, 25, -32, 2, 45, 75, 92, -109, -34, -116, 15, 59, 54, 58, -85, 120, -51, -52, 113, -86, -60, -55, -109, 26, 0, 2, 87, -94, 113, 29, 15, 41, -98, -1, -33, -6, 62, -52, 19, -20, 87, 84, -75, 44, -107, -43, 42, 28, 102, 58, -127, 98, -58, -5, -52, 34, -43, 120, 11, 63, 98, 76, -15, -8, -115, -80, 106, -15, -25, -86, -1, 51, 100, 41, -42, -87, -41, -8, 112, -68, -82, 113, 117, 112, -73, -44, -45, 28, -34, 51, -66, -43, -87, -52, 19, -62, -115, 103, -11, -82, -123, -49, 47, -26, -125, 48, 7, -52, -124, -47, -71, -116, 102, 63, -88, 59, 98, 39, -49, -27, -33, 99, 115, 123, -20, -89, 70, -17, -102, -104, -72, -67, 11, -26, 52, -27, 74, 104, 14, -39, 65, 34, -31, -120, -111, 69, -34, -87, -55, 71, 75, -4, 66, 7, -77, -127, 96, 8, -23, -110, -127, 17, 33, -65, 53, 77, -31, -7, 83, -102, -88, -96, 51, 125, -115, 98, -103, -12, -90, -9, -33, -24, -118, 7, -80, -102, 119, 37, 117, -31, -102, -58, 84, -102, -15, 41, -120, -9, -71, -113, -9, 70, -24, -58, 22, 34, 53, -70, -75, 3, 44, 119, 51, 49, 110, -116, -62, 99, 54, 50, -116, -58, 123, -10, -106, -50, 16, -4, 119, 93, 85, -90, -64, -92, -77, -42, 89, 78, -59, -108, -48, 41, 1, 17, -94, -11, -64, -80, -29, -60, 95, -23, 107, 0, 13, 82, 77, 118, 33, 17, -4, 58, -97, 29, -16, 96, 84, -102, 30, 70, 94, -50, 84, -68, -125, 0, -95, -110, 62, 61, 112, -41, 29, 97, -52, -9, -48, 105, 8, 14, 74, 79, -13, -26, -40, -87, -16, 26, -76, 124, 22, -9, -24, 121, 109, -110, -51, 55, 57, 111, 15, 65, -26, -38, -39, 12, -21, -78, -114, -98, -83, 122, -50, 24, -78, 9, -52, -71, 115, -78, -20, 41, -57, 79, -110, -1, -117, 3, -125, -84, -100, 51, 75, 23, 79, 50, -126, 102, -33, -83, -23, -49, -122, -6, -81, -107, -71, 44, -5, 27, 110, -99, 15, -25, -100, -20, -118, -32, 122, 40, -115, 80, 13, -58, -8, -9, -47, -43, -83, 5, 104, -11, -74, -106, -6, 20, -2, -109, 28, -126, 77, 15, -99, -4, 5, -105, 49, 36, -93, -125, 98, 111, -116, 52, 39, -125, 45, -122, 32, 70, -51, -82, 5, 113, -114, 114, 77, -103, -76, -120, 116, 38, 88, -58, 44, 116, 79, 12, 70, 78, 69, -50, 54, 118, -59, 57, -47, 65, 8, -100, -54, 4, -57, -15, 100, 4, 127, -20, -6, -34, -100, 92, 65, 110, 82, -2, 51, -125, -110, 74, 43, -23, -95, 6, 39, -79, 28, -15, -27, -88, 123, 106, 61, -100, 26, 78, -96, -117, 76, -51, 102, -83, 102, 41, 76, -123, -43, -59, -22, 47, -1, -26, -20, 67, 114, -64, 57, 54, 109, -94, -12, -52, 102, 34, -58, -57, -80, -50, 5, 126, -4, -9, 82, 56, -82, -19, -18, -112, -120, 51, -27, -56, -11, -97, 79, 6, -27, 102, -76, -52, -118, -90, 5, 63, -94, 82, -83, -18, -84, -106, 79, 42, 100, 4, 39, 6, 33, 76, 80, 56, 73, 90, 18, -128, -59, -66, -59, 33, -1, 0, -119, -110, -11, 44, 41, -111, 70, 62, -43, -32, -15, -96, 24, 22, -102, 77, 120, 0, 35, -65, -39, 37, -43, 21, -50, -80, 4, 56, 114, -43, 49, 86, -89, -11, -14, 35, -81, 122, 45, -84, -14, 125, -109, -18, 85, 101, 34, 108, -42, 100, 77, 46, 12, -59, -111, -37, 45, 19, -8, 33, -117, -16, -49, -68, -106, -71, -51, 0, 6, -13, 6, 74, 17, 123, -1, 53, 49, -62, 51, 69, -122, -41, 107, 63, -112, -107, -31, -26, 79, -64, 23, -66, -77, 8, 53, -65, 48, 111, -60, 88, 97, -78, 53, -104, 40, -13, -116, 90, -64, -31, -39, -105, -107, 35, 62, -94, 103, -88, -13, -116, -54, 52, 127, -4, -110, -118, -63, -94, -53, 28, -95, 61, 3, -41, -107, 124, -59, 46, -93, 68, 104, -11, 43, 6, 100, -86, -123, 106, 82, 124, -33, -40, -68, -32, -115, -57, 63, 35, -46, 35, -69, 13, -17, 28, -50, -20, -87, -69, -67, -98, 103, -110, -21, -93, 5, 121, 46, 61, -30, -106, 34, 37, 32, 51, -44, -126, -33, 123, 124, 84, -56, -26, -118, -118, -84, 41, 7, 119, -53, -58, -87, -40, -92, 44, -119, 31, 45, 82, 78, 58, -29, 41, -40, 43, 91, -109, 22, -77, 14, -34, 25, 16, 4, -35, 73, 72, -36, 15, -52, -71, -12, 98, -86, 33, -114, -15, -114, 82, -123, 116, 86, -24, -116, -94, 116, -110, -83, 12, 34, 63, 119, -20, -27, -63, -57, 49, -38, 34, -73, 9, 21, 37, -10, 90, -60, 64, -52, 63, 90, 2, 70, -31, 41, 90, 95, 31, -120, -92, -121, 21, -46, -49, -78, 89, -20, 6, 73, 52, 52, 101, -95, 114, 81, 85, -29, -19, 6, 32, -100, 1, 45, -123, 38, -37, -24, -120, 110, -111, -114, -14, -72, 69, -4, -60, -115, 32, 69, 97, -54, 25, 53, 3, -43, 62, 8, 9, 29, 81, 73, 40, 65, 41, 99, 15, -105, 18, 127, 3, -59, -116, -70, 103, -108, 79, 118, -52, 89, -10, 51, -101, -64, -24, -70, -119, 78, 53, 92, 56, 14, -45, 86, 106, -9, -128, -124, 63, -113, -128, -5, 40, -18, -115, -18, 118, -119, -65, 115, -101, 70, 87, 94, 106, 21, -86, -119, -52, -99, 72, 15, -4, 4, 19, -72, 102, -41, -30, 8, -37, -92, 117, 65, -96, 89, 65, 7, -1, -23, -26, 43, -128, 69, -36, 16, 83, 56, 59, 56, -125, 25, 73, 68, -80, -60, -90, 100, -91, -67, 67, -122, -115, 73, 98, 98, 112, -35, 103, 96, -38, -123, -16, -4, -57, -11, -92, -31, -34, -92, -104, -64, -106, -83, 4, -125, 116, 100, 7, -87, 112, -38, -64, -30, 104, 121, -32, 9, -84, 44, -82, 51, 119, 56, -111, 26, 82, 51, -39, 51, -87, 37, 52, 38, -47, 126, 103, 38, 21, 88, -106, -75, 0, 28, -5, -122, -8, -75, -10, 86, -89, -35, 95, 0, -28, 117, 12, -4, 65, 78, 16, 13, -127, -60, 45, -105, -109, -42, 21, 27, 14, -26, -30, 18, -19, -61, -57, -43, -83, 86, 87, 123, 83, 1, -113, -27, 114, 80, 69, 24, 66, 60, 40, -11, -10, 57, -114, -26, 29, -95, 91, 112, -36, -88, -51, -76, -43, -121, -125, 24, -45, -27, -128, 0, 0, -15, 84, -117, 67, -122, 10, -55, 67, -34, 31, 53, -122, 14, 26, 92, 121, -71, 30, 42, 35, 93, -70, 102, 89, 111, 12, 52, 11, 28, 72, 93, -16, -68, 62, -58, 84, 57, 105, -10, -110, -63, -99, 97, -57, 94, 56, -78, -60, -40, 43, -122, -57, 8, 25, -84, 56, -2, -127, -39, 82, -121, 36, 42, -20, 18, 31, 1, 66, 83, 21, -99, 42, -19, 52, 41, 52, 30, 39, 104, 13, 95, -23, 107, 4, 97, 28, 6, 79, -32, 52, 46, 42, -5, -25, 77, -23, -72, -124, 106, -60, 33, 6, 26, -31, 5, -7, 68, 54, -96, -5, -42, 116, 1, 111, 49, -105, 118, -24, 6, -2, -54, 83, -36, 81, 83, 100, 106, -70, -30, 16, -94, -86, 52, -56, -25, -33, 20, 55, 65, 115, 81, -15, -16, -59, -32, 75, -111, -73, -33, -18, 60, 10, -58, -63, -40, 91, -104, 20, 51, 118, 64, -104, 6, 45, -91, 43, -2, -22, 58, -112, 114, 87, 15, -2, -80, -55, 44, -40, -45, 53, 87, 113, 56, -90, -8, -83, -23, 106, -37, 22, -120, 15, 34, -114, -64, -119, -39, -109, 64, 54, 23, 87, 87, 77, 123, 102, 44, 78, 111, -118, -46, -86, -16, -73, -81, -113, -122, -108, -50, -66, -42, -41, 8, 95, 113, 67, 90, -35, 34, 22, 118, 76, 79, 32, -117, 5, -24, 104, 85, 104, 77, -92, -15, -18, 20, 93, -17, -87, 50, -56, 115, -29, 31, -85, 56, 101, -98, -25, -16, -20, -71, 39, -6, 94, 22, 97, 100, 24, -13, 11, -47, 28, -19, -121, 46, -110, -92, -80, 6, 41, -125, 43, -91, -106, 60, -86, -13, 25, -118, -124, -119, -51, 1, 63, -16, 106, 74, -12, 92, 96, 46, 31, -41, -48, -120, -71, 107, 47, 116, 41, -31, -30, 86, 49, 4, -83, 9, -62, -77, 72, 84, -25, 13, 85, 109, -82, -44, 58, -41, 93, 68, -28, -85, 69, -8, 74, 124, 123, -79, 82, 3, 48, -111, 75, -128, 2, -6, 117, -89, -96, -58, -36, 40, -79, -17, 23, -74, 122, 119, -117, 18, -39, -107, 61, -7, 69, -65, -98, 24, -3, -12, -23, 94, 97, 18, -28, -121, -119, 124, 45, 77, 123, -54, -99, 50, -38, -21, 104, 90, 78, 91, 28, 41, -111, -17, -119, -120, 65, 5, -82, -115, 59, 51, -108, -81, -76, -61, 51, -121, 109, 116, -46, -111, 24, 18, 118, -15, -41, 49, 95, 11, -33, -91, 127, -2, -30, 27, 53, -45, 2, -90, -19, -45, -101, 59, 11, -36, 66, -128, 83, -119, 34, 54, 73, -8, -92, -51, -43, -83, 59, -50, -56, 58, -32, -26, -29, 61, -67, -81, -85, 11, 112, 41, -75, 61, 101, -51, -40, -12, 56, 6, -94, 3, 44, 3, -27, -53, -111, 24, 94, -125, 72, 8, -121, 67, 120, -10, 64, -32, 67, 34, -104, 82, 49, 83, -67, -77, -58, -65, 21, 57, -111, -34, -65, -79, 89, -114, 37, -119, 86, 6, 13, 117, -101, 99, -63, 26, 58, -18, -97, -91, 72, 42, 117, 31, 117, 18, 39, 25, 119, 34, -73, -48, -19, -12, 63, -11, 106, -66, -56, 60, -78, -127, 41, 15, -23, -9, -66, -100, 75, -112, 110, 37, -37, 74, -47, 120, 101, -119, 106, 80, -28, 36, -17, 52, -9, -89, -10, -50, -97, -103, 9, -54, -87, -125, -6, -98, 32, -22, 28, -37, -103, 23, 106, -57, -98, -110, 1, 102, -112, -48, -32, -104, 30, 49, -23, -63, 88, -122, -128, 28, -108, -69, -51, -15, -18, 109, -108, 82, -43, 40, 29, 99, -120, -87, 96, -39, 94, -92, 93, -29, -81, 117, 95, 14, -38, -124, 51, -86, 110, -25, 56, 95, -58, 54, 38, -93, -74, -51, 125, 115, -113, 70, -123, 54, 94, -78, -65, -85, 119, -50, 49, 115, -29, 31, 66, -58, 25, 91, 23, -46, 102, -22, -14, 109, 28, -115, -76, -119, -36, 42, -69, -28, 34, -11, -61, 7, -104, 93, -35, -41, 45, 44, 57, 43, -59, 24, 71, -56, 55, 55, -115, -17, -67, 72, 68, 48, 107, -22, 80, -26, -84, 74, -4, -33, -93, -16, -12, -104, 120, 23, -62, 102, 42, -86, -108, 104, 103, 108, -28, -9, 89, -107, 12, -26, -18, -35, 44, 43, -15, -67, 4, 108, 80, -83, -26, 58, -106, 76, -71, 41, 90, -39, -97, 33, -84, 6, 95, -48, 75, 66, -90, 113, 87, -113, 75, -49, -25, 12, 115, 116, 75, 98, 12, -6, 99, 126, -57, 108, 15, 115, 58, 12, -20, -47, 122, -8, 95, 67, 80, -60, 92, -10, -79, -61, -102, -120, 84, 76, 114, 67, -13, 63, 121, -14, -99, 115, -61, 96, 77, -80, -100, 52, -52, 39, -17, 0, 32, -2, 85, -96, 6, -62, 25, -92, 78, -71, -94, 91, -29, -50, 47, -110, 22, -23, 87, 35, -125, -43, -49, -44, 63, 32, -48, 113, 48, 78, 71, -57, 82, -41, 12, -115, 114, 69, 59, 126, -32, 15, -21, 107, -3, 85, 76, -1, 53, 27, -68, 39, -124, -1, -37, -115, 35, -42, -72, 28, 46, -124, -101, -22, -15, -120, 48, -104, 65, 28, 59, 105, -64, -97, -105, 54, -120, 13, 59, -85, 4, 72, 74, -16, 43, -22, 117, 104, 45, 67, 108, -118, 86, -60, 3, -8, 90, -94, 52, 18, 101, 57, -50, -45, 111, 6, -8, 67, -92, -91, -73, 115, 67, -46, -28, -81, -51, -90, 47, 47, -119, 38, 92, 115, 31, 62, 7, -53, 65, 122, 52, 100, 85, 117, 50, -30, 4, -95, -5, -5, 20, 32, 94, 69, -38, -14, -16, 57, -52, -10, 18, 74, -10, -50, -86, 90, -53, -62, 22, 105, 40, -16, -115, 46, 117, -95, -119, 82, -79, -109, 10, -99, 10, 121, 34, 70, 8, 115, -78, 25, 17, 87, 43, -33, -42, 35, -64, -103, 103, 66, -10, -20, 74, 38, 63, -3, 34, -48, 26, 33, -22, 37, -29, 103, 38, -27, -56, 13, -80, 9, 80, -54, 0, 14, 41, 54, 84, -76, 27, 33, -54, -30, 126, 44, -106, -81, 22, -24, -15, -8, -41, 96, -117, 59, 110, 70, -14, 121, 122, -46, 48, -43, 35, -36, -34, 2, 15, 49, 73, 11, -30, -50, 22, -99, -101, 29, 21, 118, -126, 2, -120, -105, 19, -68, -55, -94, -2, 92, 123, 73, -105, 83, 77, -28, 0, -26, 84, 31, 100, -47, -66, -58, -33, -14, -120, -59, -83, 74, -91, -81, 95, 16, 27, 127, 15, -85, 30, -49, -93, -56, 73, 35, -91, 13, 72, 127, -60, 114, -79, 19, -99, -63, 43, -20, -37, -111, -105, 102, -54, -34, -91, -10, 53, 26, 12, 60, -120, -65, 57, 21, 16, -5, -92, -106, 79, 114, -126, -95, -99, 73, 39, -26, -21, -19, -127, -49, -48, 33, 18, 21, 104, 32, 102, 86, -60, 63, 22, -111, 47, -114, 21, -67, -78, 89, 93, -7, 87, -10, 125, -26, 123, -125, 126, -14, -28, 63, 56, 124, 13, -7, 51, 12, -18, 109, -13, -126, -50, 116, -68, 76, 35, 110, -54, 2, -4, -75, -110, 92, 80, -2, 51, 114, 59, -10, 40, 56, -27, -19, -99, -104, 81, -72, 117, 122, 108, -62, -122, 63, -18, -105, -1, 23, -18, 48, -87, -77, 51, -110, -93, 61, -27, 51, -75, -82, 73, -108, 9, 88, -95, -18, 25, -23, -15, 113, -89, -120, 68, -94, -21, 107, -118, -46, 53, 21, -53, 18, -128, -15, 100, -90, -34, 3, 80, 91, 83, 40, -102, -105, -62, 41, -12, 64, 9, -9, 122, -87, -126, -70, -66, 23, 67, -103, -106, -127, -83, 40, -67, 81, 68, 30, 29, -49, 4, 52, 30, -122, 99, -68, -26, -118, 17, -64, 18, -101, 94, -3, 76, -55, 111, 103, 51, 75, -96, 119, -42, -43, 30, 0, -15, -6, -116, -35, 110, -21, 117, -40, 41, 2, 37, 61, 12, -101, 60, -107, 122, -10, -66, -92, 97, 98, -96, -73, 5, -118, 66, -83, 89, -31, -125, 79, -13, 40, -15, -18, 17, 121, 122, 8, 16, -18, -24, 52, -46, -72, 107, -117, 17, 46, 109, -97, -49, 29, -26, -20, -104, -25, -107, 81, 26, -57, 79, 117, -6, 106, 116, -18, 29, -5, 74, 8, -4, 79, -100, 42, -69, 88, -95, 80, 35, 118, 58, -89, 66, -71, -99, -111, 24, -27, -18, 117, -75, -125, -48, 52, -93, 34, -33, 71, 76, -18, 17, 62, -33, 125, 76, 66, 8, -86, -21, -38, 122, -115, -73, 116, -99, 59, 88, 122, 93, -21, 86, -109, -4, -12, 116, 45, 72, 87, 37, -95, 30, 7, 101, -48, 13, -67, -69, 25, 36, 21, -124, 29, -102, -14, 72, 17, -77, -88, -52, 62, 107, 3, 4, -21, 102, -128, -71, -121, 119, -10, -87, 61, -78, -105, 93, 106, -84, 47, -92, -105, 48, 76, -34, -77, 46, -66, -66, 60, -117, 67, 74, 108, 29, 23, 125, 123, -76, 67, 35, 25, -84, -41, 114, -84, -27, 16, -123, 92, -13, -6, 92, -117, -67, 37, 37, 9, -76, 94, -28, 5, 45, -70, -47, 108, 66, -46, 46, 20, -28, 28, 68, -47, 42, -9, 65, 71, 20, -17, -67, 60, -7, -76, 26, 45, 35, 99, 23, 116, -68, -100, -60, 73, 62, 115, -112, -19, -45, 115, 56, -50, -76, 75, 25, 77, 89, -109, 88, 100, -55, 88, 35, 94, 89, 8, -71, -103, 113, -89, -7, -23, 122, -120, 118, 39, 85, -9, 35, 25, 119, 20, -102, -60, -74, -50, 83, 114, 99, 107, -63, -65, 40, -99, 59, 75, -40, 95, -86, 34, 22, -24, 74, 106, 8, -109, -114, 104, 91, 57, -21, 70, 39, 74, 89, 4, -36, 66, -16, -40, -103, 113, 5, -47, 107, -30, 15, -63, 9, 20, -86, -109, -47, -76, -128, 120, -57, 63, 29, -8, 92, -7, 44, -5, -1, 109, 110, -127, -123, 75, 109, 76, -31, 72, -26, -11, 46, -59, -82, -10, 108, 73, 65, -122, 78, 76, 91, -78, -18, -112, 84, 23, -61, -58, 74, 70, 0, 78, -15, -50, 113, -112, -87, -39, -116, -103, -40, 113, -27, 20, -34, -86, -49, -20, -46, 114, 61, 21, -36, 30, -4, 62, -93, 96, -66, -76, -126, -37, 27, 36, 5, 109, 28, 103, 108, 54, -104, 55, 119, 63, -76, -68, 4, 60, 80, -33, 82, -13, 4, 70, -79, 73, -61, 107, -125, 116, 84, -101, 30, 75, -121, -97, 93, -58, -104, -112, 89, -127, -84, -11, -46, -96, -105, 20, -87, -11, 61, -29, -20, -67, 43, -54, -106, -39, 11, 117, -102, 63, -41, -19, 102, 29, 119, 13, 56, 126, 97, 111, 88, 83, 15, -104, -79, -115, -75, -50, -6, -32, 47, 51, 59, -25, -18, -78, -79, 121, -68, 65, 121, -58, 77, -7, -92, -31, 33, 43, 107, -90, 65, -28, -107, -66, -75, 64, 127, 57, 107, -18, -46, 19, 43, -80, -88, -73, 1, -25, 106, 30, -10, -102, -13, 38, -31, -88, -68, 111, -43, 30, -119, -14, 110, 22, -57, -106, -11, -91, 37, 56, 32, -92, -87, 68, 35, -115, -98, -77, 112, 62, -9, 66, -62, 43, -74, 50, 100, -89, 65, 116, 106, -100, -92, 47, -56, 64, -94, 9, 93, 40, -104, -44, -60, -73, -42, -6, -57, -80, 46, -126, -30, -85, 118, 41, -40, 28, 46, -68, 93, -75, 43, -43, 27, -20, -29, -103, 109, -43, 0, 37, -11, 14, -12, 32, 110, -88, -11, 90, 20, 51, -104, 101, 46, -89, 75, 23, -68, -37, -12, 8, 113, 28, 105, -69, 33, -61, 14, -70, 51, 23, -127, 111, -29, 26, 124, 8, -36, -97, 13, 54, -42, -27, 58, -116, -107, 64, 2, 32, -95, 2, -76, -34, 90, 1, 88, -51, -62, -66, 3, -42, 88, 62, -13, -81, 20, 83, -97, 55, -105, 127, -45, 24, -92, -62, 113, -9, -55, -41, -101, 10, -1, 47, 55, -20, 33, 42, -112, -5, -126, -62, 70, 82, 50, 95, -55, 46, 62, 115, -108, -63, 12, 63, 127, 31, -114, -89, -115, 35, -73, -8, 118, -23, 15, -86, -80, -45, -72, -59, 54, -51, 6, 43, -39, 21, -54, 48, 17, 123, 40, 120, -45, 66, 6, 73, -22, -74, 116, -93, 88, 64, -87, 81, 109, 57, -122, 40, 37, -46, -50, -38, 94, 108, -30, -89, 26, 82, 86, -46, -119, -75, 67, 66, 1, 34, 118, -66, -43, 118, -65, -3, -65, 83, 15, -54, 109, 58, -41, 60, 68, 111, -25, -82, -40, -19, -55, -114, 44, -87, -1, 60, -51, 88, 126, 17, 14, 91, -26, -68, -63, 34, -52, 8, -23, -89, -64, -119, -87, -110, -111, -17, -9, -47, -110, 42, 16, 121, -87, 4, 95, 41, 45, 72, 89, -19, -84, -58, -120, 78, -95, -68, 57, -47, 46, 93, 36, -52, 103, 42, 120, -75, -33, -24, 43, -15, -107, 127, 68, 15, 87, -85, -51, 118, -124, 37, -1, 16, 21, 77, 80, 77, -87, -8, -116, 27, -127, 42, 73, 63, 103, 17, -76, 24, 122, 112, -38, -89, 87, 7, 72, -102, 117, -39, 35, 36, -24, -90, 24, -86, -104, 126, -9, 83, 30, -95, -60, 16, -79, 51, -23, -89, -31, 49, 119, 107, 115, -96, -126, 52, -81, 87, 81, -56, 107, -15, 68, -90, -102, 97, 75, 76, 27, 84, -113, -76, -114, 47, -13, 7, -92, -45, -43, -118, 34, 27, -97, -11, -38, -93, -33, 9, -11, -22, -33, -71, 24, 115, -47, -66, 89, 79, -36, -115, -31, 107, 0, 27, 62, 38, 119, 73, 85, 99, -112, 59, -128, 93, -105, -28, 42, 18, -90, 45, 121, -43, 99, 27, 21, 8, -117, 110, -84, 32, -30, -44, 89, -66, -76, -77, 82, -54, -62, -88, 40, -62, 43, 5, 26, -14, -119, 126, -81, -35, 3, 86, -87, -2, 1, 29, 63, -40, -24, 90, 40, -25, -98, -52, 41, 65, -80, 43, 12, 115, -40, 81, 0, -66, -64, 119, -118, -58, 31, 43, 0, 123, 93, -15, -30, -76, -76, -71, 19, 97, -2, -32, -72, -49, -110, 70, 75, 67, -103, 15, -36, 124, -20, 110, -54, 29, 62, -41, -44, -117, 45, -3, -118, -72, -2, -14, -1, 122, 62, -85, 6, 64, -122, 71, 38, -42, -96, 89, -89, 75, 26, -3, -24, -85, -51, -117, 54, 114, -108, -28, 29, -46, -45, -33, -79, 60, 122, -43, -38, -124, -62, -64, 109, 107, 2, -4, -58, -127, 33, 30, -113, -83, -84, 45, -39, -78, 52, -34, 101, 99, 87, -56, -90, -103, 58, 103, 40, 94, -13, 29, -50, 21, -95, 30, -76, -99, 88, 116, 43, -58, 123, -77, -33, -123, 126, -120, 28, 101, 18, 4, 57, -106, -37, 103, -96, 123, -67, -97, 73, 30, 112, 1, 103, -33, 87, -64, -14, 23, 36, 29, -3, 2, -36, -91, -66, 82, 71, -41, 119, -41, 111, 65, 22, -109, -11, -50, 94, -2, 123, -14, -81, 110, 96, -54, -43, 64, -85, 45, -90, -127, -109, 23, -46, -66, -82, 119, -61, 83, 102, -117, -125, 57, 40, 68, -80, -11, -118, -40, 112, -19, 65, 72, 108, -48, 11, -11, -56, -60, -90, 97, -110, 85, -119, -7, -46, -118, 71, 119, 88, -57, -22, -8, 7, -106, 105, 95, 65, -20, 41, 31, 72, 97, 43, 29, 104, -93, 37, 3, 102, 16, 71, 23, 18, -2, -42, 86, 42, -64, 116, -123, -35, 9, -87, 96, -128, -41, -122, 53, 62, -12, -26, -107, 5, -23, 121, -77, 60, 109, 25, 116, -30, -56, 67, -88, 36, -65, -50, 104, 30, 70, -76, -99, -72, 8, -18, -80, 115, -28, -97, -94, -1, 65, 83, 53, -7, 86, 102, 123, 27, -105, -9, 32, -114, -5, 48, 120, 58, -77, -82, -97, -4, -88, -3, 69, 108, -112, 103, -55, -115, 112, 85, 63, -73, -82, 40, -7, 14, 76, 81, -128, 80, -3, 92, 5, 32, 51, -102, -107, 29, -38, -80, -13, -57, -92, -63, 84, 4, 14, -60, 17, -43, -43, -72, -22, 98, 69, 42, -128, -124, 116, -97, 104, -34, 22, 127, -9, -91, -12, -74, -101, -50, -13, -100, -11, -91, -87, -93, 50, -64, 6, -8, -72, -57, 111, 42, -19, 92, -101, -23, -128, 104, -126, 22, -75, 5, 54, 18, -97, 120, 7, 85, -54, -11, 71, 13, -1, -30, -72, 29, -3, -24, -107, -127, 4, -46, -120, 62, -107, 28, 8, 39, 20, -83, -50, 55, 4, 80, -5, -47, -4, 42, 89, -95, 31, 29, 113, 109, 77, -8, -14, -62, -52, -119, 119, 112, -68, -118, 101, -110, 59, -94, -67, -122, 36, -117, 2, 38, 120, 78, -124, -103, -7, -116, -8, 27, -38, -29, -116, -20, 50, 90, -48, -31, 121, 93, -55, 73, -76, -90, 103, 38, 41, -42, 84, -52, -36, 118, 105, 74, 80, 122, -71, 7, -43, -112, -25, 72, -125, -102, -42, 41, 19, 111, -30, -104, -15, 40, -82, -80, -31, -61, 60, -43, -52, -78, 72, 127, -84, -100, -11, -81, -82, -19, -48, 34, 41, -21, -41, -83, 69, -101, -117, -116, 39, 48, 63, 119, -66, 67, -17, -106, 124, -42, -107, 63, 101, -108, 81, 101, -60, 100, -123, 16, 91, -48, -105, -2, -2, 4, 80, 1, 16, 117, -62, 43, 120, 52, 23, 47, -108, 79, -11, -114, -38, -73, 119, -7, -65, 23, 118, -48, -123, 74, 113, 59, 21, 108, 48, 96, -30, -50, -45, 31, 32, -60, -69, 70, 16, -92, -97, 74, 51, -25, 56, -7, -25, -11, -60, -29, -68, 55, 65, 5, -24, -61, -89, -122, -128, -59, -91, 63, -8, -65, 105, -124, 4, -31, 4, 113, 7, 73, -93, 13, 47, -13, -124, -2, -35, -115, -26, -74, 12, -8, -119, 63, -80, -69, 108, -128, 96, -56, 127, -64, 68, 48, -94, -73, 15, -67, 68, 96, -63, 104, -123, 24, -49, 34, 110, 98, -127, 70, 125, -92, 126, -111, 23, 23, 68, 56, -65, 76, -106, 40, 98, 10, -64, 46, -96, 70, -83, 82, -47, 37, -20, 62, -18, -36, -19, 91, 32, -110, -50, -99, 115, -78, -4, -98, 90, 37, 79, -21, 67, 95, -32, -107, 124, 1, -19, -107, 76, 115, -26, -49, -4, 37, 19, -83, -57, -64, 73, 88, -2, 112, -16, 34, -62, -11, -111, -50, -33, -110, -53, 122, 115, 110, 2, 44, 126, 36, 22, 83, -72, -59, -33, -114, -77, 116, -2, 82, 75, -88, -48, -68, 21, -98, 14, 86, -19, 97, -96, 13, 77, 2, -15, 82, -82, -96, 32, 125, 104, 111, -83, -36, 103, 77, -32, -96, -34, 115, 1, -114, 95, 60, 85, -128, -4, 83, -72, 102, -80, 66, 19, 58, 75, -109, 74, -4, 124, 79, 98, -125, -116, -90, 121, -49, 66, 13, 107, -55, 60, 44, 79, -60, 2, 38, -5, -52, 79, -118, -7, -124, -102, -102, 84, 3, -76, -21, -43, 104, -37, 82, 54, 84, 80, -25, -86, 59, -42, -93, -11, 12, 88, 74, -49, -65, -65, 11, -113, 39, 107, 100, -17, -13, -113, 36, 96, 12, 101, 76, 81, 83, -123, 119, -10, 10, -42, 48, 37, 99, 39, -28, -33, 55, 71, 121, 84, -64, -106, 11, -19, 104, 108, -41, -16, 78, 86, -83, 77, 47, -51, 120, -28, -101, 17, -123, 3, -95, 21, 108, 105, -7, -12, 87, -65, -112, -74, -47, 76, 80, -43, 71, 77, 121, 31, -17, 18, 25, -61, -107, 9, 83, -6, 84, 75, -51, 93, 63, -74, 60, 37, -105, -99, -62, -14, 30, -119, 26, -20, -86, 57, 40, 38, 5, -17, 0, 39, 91, 90, 2, 5, -14, -104, -94, 38, -97, 114, 35, -16, -51, -48, -28, -1, 122, 60, 19, 95, -85, 11, -68, -52, -114, 45, -117, 54, -32, 105, -110, -40, -57, -116, 36, 59, 51, -106, -69, -106, 77, -98, 111, 89, -100, 36, -76, 17, -90, -34, 88, 89, -105, 23, 98, 61, -32, -20, 12, 39, -81, -103, -91, -54, 7, 14, 2, 55, -57, -11, -46, 49, 24, -84, 58, -54, -11, 100, -40, -64, 0, -76, 74, -30, 86, -107, 63, -72, 68, -23, 87, -44, 88, -83, 60, 66, 116, -127, 104, 11, -22, -121, -57, 72, 36, -22, -75, 104, -84, 27, 2, -1, -79, -96, 5, 65, 114, -89, 83, -3, -61, 18, 107, -92, 81, 85, -64, 17, -108, -90, -27, -121, 52, 25, -118, 87, 94, 67, -103, 63, -57, -33, 113, -42, 49, 82, -123, -51, 51, -97, 36, 25, -5, 19, 122, 65, 7, -4, 115, -38, 123, 61, 14, 125, -82, -106, -49, 62, 113, -87, -93, 6, 40, -38, 15, -80, 60, 29, -36, -47, 19, 109, 48, -66, -11, -7, 40, 63, -127, -79, -121, 84, 32, -27, 94, -12, 19, -41, -93, -91, 29, 80, -1, 118, 58, 73, 88, 62, -6, -124, -39, 77, -80, -95, 81, 62, 95, 108, 39, 25, 55, -68, 53, 56, -25, -21, -47, 34, 107, -70, 47, -122, 81, -124, 126, -35, 60, -81, 16, -52, -61, 74, -121, -117, 112, -90, 67, -62, -56, 69, -1, 51, 52, -126, 111, -74, -64, 55, 41, -17, 77, 56, -38, 18, -64, 48, -80, 42, -115, 111, 23, 91, 1, -48, -21, 32, 86, 41, -57, 37, -116, 89, -121, -76, 92, 105, 35, 88, 1, -63, -6, 70, -95, 47, -19, 104, -86, 0, 80, 102, 50, -15, -57, -123, 123, -119, -107, 72, -62, -22, 28, 45, 1, -38, 106, 101, -4, -21, -45, 7, 124, 47, -126, 5, -71, 51, 41, 118, -95, 26, -58, -126, -37, -22, 99, -105, -128, 83, 84, 73, 54, 49, 75, 93, -53, -40, -53, -68, 71, 92, -63, 36, -120, 86, 117, -97, -22, 36, -103, 15, 10, -115, -18, 85, 73, -38, -97, -28, 21, 103, 127, -36, 93, -57, 89, -51, 116, -81, 9, -5, -25, 98, -119, -77, 92, -7, 101, 28, 7, 106, -43, 10, -76, 38, -78, -127, 33, -113, 79, -107, -50, -49, 61, -29, 75, 67, 51, 116, -124, 16, 93, -33, -71, 100, 46, 10, -104, -27, -10, -55, -55, -4, -22, -80, 100, -15, 84, -54, 67, 36, -59, -102, -83, -67, -90, 95, 27, -103, -11, 98, 39, -57, -80, -44, 103, 79, -33, 97, 102, -119, -71, -82, -8, 23, -14, -9, 65, 78, 98, -30, 57, 124, -93, -24, -66, 32, -40, 66, -104, -108, 45, -95, -115, 10, 86, 116, 124, -84, 66, 96, 60, 4, 69, 2, 17, 3, -124, -40, -80, 74, 72, -87, 122, 48, 116, -46, -107, 78, 64, -12, -85, -77, 102, -29, 84, -30, 23, -124, -48, -22, 4, 97, 110, -112, 114, 10, 3, -98, 62, -95, -105, 43, -9, -93, -102, -3, -95, -60, 15, -44, 89, -112, -101, 119, -31, 67, -19, -47, 66, 63, -28, -115, 117, 107, 20, 45, -56, -26, -11, -3, -4, 23, -44, -39, 125, -93, 127, 38, -12, -59, -31, 65, 35, -2, 49, 7, -44, -120, 98, -114, -67, 12, -35, -117, 51, -16, 121, 34, -7, -57, -4, -39, -31, -9, -104, 66, -101, -27, 24, 62, -8, 99, -25, 110, -69, -54, -45, 90, -79, 55, 102, -45, -12, 126, -17, -104, -9, -85, 74, -74, 13, -64, 85, 103, -34, 19, -108, -1, -33, -122, 5, 39, 125, -33, 51, 12, 104, -78, -76, 105, 40, -118, -96, -6, 52, 115, 111, 23, -87, -68, 5, -11, -111, -3, 116, -83, -48, -98, 82, -29, 7, 32, 18, -45, 51, 12, -128, -23, 36, -16, -27, -81, -65, -78, -63, -16, -86, -127, 48, 9, 12, 25, -45, 0, 61, -95, -34, -65, -69, -86, 56, -88, 127, 126, 29, 75, 53, -73, 23, -82, 81, -111, 44, -54, 66, -63, -33, -24, 15, 114, -69, -102, 25, -92, 1, 119, 66, 74, -60, -127, 66, 40, -25, -100, 63, -86, 103, 127, 107, 104, 84, 124, 16, -83, 61, 90, 26, 111, 68, -82, 24, 60, 35, -25, 37, 25, 81, -87, -18, -21, 34, -6, -29, -67, 33, 48, 0, -92, -55, -8, 70, 56, 124, -76, 84, 93, 43, -102, 8, -80, -76, 100, -61, 105, -10, 66, 66, 14, -71, 53, -28, -107, -75, 36, 70, -109, -77, 24, 92, 70, 56, -41, -82, 7, -73, 126, -65, -95, 89, 77, -57, -34, 98, 71, 87, 37, -92, 116, -50, 116, 15, -125, 124, 36, -106, 78, 20, 30, 60, -64, -29, 1, 37, 85, -95, 109, -117, 55, 63, 78, 13, -21, 46, -21, 122, 60, -62, -56, -32, 117, -15, -15, 86, 124, -56, 5, -93, 25, 99, -70, 118, 62, -109, 38, -57, 85, 111, -87, 103, 25, 84, 124, -3, -41, 114, 93, 9, -60, 111, -107, -51, -26, -115, 66, -78, 70, 86, 57, 57, 117, 88, 24, 64, -55, -104, -42, -88, -52, -37, 88, 123, -114, -127, -125, -72, -59, -72, -26, -46, -114, -121, -41, 102, -116, 92, -48, 39, -79, -81, 42, 27, -70, 72, -87, 14, -83, 101, 26, 3, 42, -60, -71, -98, -29, 89, 45, -66, 57, 0, -3, 8, -92, -128, -43, 74, 88, 87, 62, 48, -29, 116, -22, 31, 84, -94, 36, 104, 101, -23, 97, 68, 51, -74, -98, 123, 19, -107, -77, 108, -107, -81, -113, -43, -79, 85, 74, 111, 93, 105, -108, 117, -75, 41, 2, -59, 109, -66, -78, 106, 87, 21, 28, -10, 2, 12, 125, -56, -50, 80, -76, 104, 48, -89, -108, -91, 122, 42, -127, -17, -117, 73, -6, 100, -56, -99, -124, -44, 121, 99, -53, 102, 65, -35, 57, -3, -27, -75, -117, -35, 117, -79, 32, -110, -31, -45, 24, 73, -47, 95, -55, 41, 1, -87, -50, 114, 32, 81, -92, 1, -27, -3, -94, 40, 2, -21, -66, 96, -31, 69, -74, 4, 21, 46, 12, 64, 53, 61, -5, 1, -2, -60, 52, 69, 59, -13, 96, 60, 45, -108, -56, 73, -89, 16, 14, -85, -61, -65, -104, 42, 5, 67, -98, 115, -124, -39, -3, -73, 53, -118, -12, -123, -13, -31, 36, 44, -18, -53, 121, -20, 89, 54, -34, 46, 109, -123, -53, -88, 53, 56, 16, -21, -20, -85, 113, 21, 121, 71, -5, 11, 57, 17, -69, 24, -13, -111, 29, 125, 47, -31, -65, 86, -71, -6, 68, 44, -103, -118, 127, 26, 51, -110, 121, 64, 114, 5, -31, -68, -40, 101, -79, 25, -118, -24, -38, -4, -67, 15, 110, -37, -95, -20, 34, -107, 100, 120, -105, 38, 21, -64, 57, -67, -71, 89, 44, -45, 38, 15, -26, -126, -80, -70, -21, -14, -54, -51, -29, 55, 42, 8, -121, 123, 67, -81, -76, 49, -115, 49, -35, 124, 102, 3, -90, -17, 117, -83, -10, 27, 95, 72, 40, 20, -73, 74, -17, -74, 15, 121, -76, -4, 70, 93, -59, 85, -99, 62, -99, 17, 69, -43, -12, 10, 15, 119, 84, -43, 8, -24, 23, -87, 87, 73, -120, 110, 104, 64, 28, -126, -89, -103, 34, 36, -61, 110, 18, 18, -4, 55, 45, -103, 2, -52, -101, -94, 46, -98, 43, -24, 29, -68, 28, -17, 124, 48, 28, 42, -123, -62, 82, -72, 3, -58, 91, 99, -77, 120, -68, 18, -11, 86, 27, 1, -1, -21, -114, -117, 38, 93, 37, 81, 94, -18, -24, -119, 71, 70, 76, -79, -36, -60, -45, -1, -4, -27, -19, -15, -16, 5, 127, 64, 63, 68, 62, -75, -14, 57, -117, -120, -93, 35, -29, -99, 124, -91, -93, -83, -92, 83, -95, 37, -15, -83, 121, -86, 2, -11, -27, -54, 117, 116, 45, 75, 25, -29, -117, 32, 74, -5, -46, -97, 52, 59, 43, 15, -1, 60, -17, 23, -12, 49, -126, 57, -4, 110, -7, 112, -48, -73, 0, 43, -103, -37, 13, -124, -99, -6, 115, 79, -127, 112, 91, 85, -64, 17, -37, -28, 47, 11, -37, -80, -87, 10, 111, -47, -110, -53, -94, 40, -95, -54, 127, 100, 15, -32, -53, 25, -109, -29, 50, -64, 78, -83, 45, -24, 104, -16, 115, -26, 76, 9, 87, -73, 2, -68, -101, -89, -37, -82, 113, 106, -97, -125, 7, -123, 90, -16, -11, -103, 2, 108, 78, -61, 96, -111, -13, 102, -76, 108, -112, -108, 120, -40, 35, -31, 12, 25, -31, 61, -106, 84, -110, -90, -112, -120, 19, -70, 67, 111, 61, -59, 111, -30, 14, 53, -3, 91, -111, 105, -56, 71, 84, 15, -35, -9, -74, 110, -43, 55, 106, 103, -58, -10, -72, -80, -63, -70, -1, 112, 72, -55, 18, -64, -58, 30, -62, -13, 79, -60, 105, 82, 32, -70, -103, -93, -67, 24, 101, -11, -7, 11, -73, 16, -3, -75, -14, -5, -124, -124, 72, 18, 106, 104, 42, -30, -78, -42, -65, -120, -72, -22, -27, 86, 122, 35, 115, 47, -118, -91, -92, 52, -28, 33, 22, 127, -57, -3, -7, -44, 49, -26, 107, -92, -10, 41, -30, -90, -36, -113, 36, -74, 29, -22, -73, -48, 119, 102, 54, 62, 57, -104, -23, 87, 70, 59, -96, -111, 120, -20, 127, -120, 4, -83, -109, -32, -85, 89, -32, 66, -15, -116, 76, 51, 12, -122, 15, -121, -97, -2, -76, -34, -53, -43, -107, -123, -24, 11, 92, -15, -20, -7, 42, -34, 68, 113, 15, -75, -34, 2, -57, 51, 4, 19, 79, -52, -78, 51, -26, 126, -111, 108, 82, 15, 12, -36, 40, -58, -61, 56, -21, 117, -5, -53, 118, -9, -92, 116, 114, 1, -56, 105, 125, -107, -13, 126, -57, 54, 58, -35, 66, 81, 71, -91, -87, 117, -79, -57, -50, -36, 33, 118, 76, 30, -25, 2, 85, 62, -79, -32, -104, 50, -104, 122, -107, -38, 89, -46, 125, -108, 118, -2, -30, -83, -93, -78, 74, -57, 38, 63, -45, -79, -40, -73, 11, -49, 112, 125, 41, 71, -108, 58, -15, -19, -64, -48, 122, -125, -94, 11, -123, 107, 62, 22, -33, 108, -35, -108, -13, -72, -9, 20, -35, -23, 93, -67, -61, 82, -16, -111, 78, 93, -63, -81, -115, 111, 68, -77, 110, 54, -124, -88, -25, 57, 51, 46, -11, -21, 81, 118, 93, 75, -88, 4, -54, -78, 111, -118, 116, 54, 34, -27, -100, -27, 90, -115, -73, -104, 104, 92, 109, -98, -112, 122, 89, 23, -120, -80, -112, 29, -66, 84, -120, 59, -23, 107, -74, -3, -101, -28, -121, 39, 22, 54, -78, 125, 19, -99, 123, 75, -83, 88, -45, -45, -44, -123, 85, 18, -77, 11, -108, -61, -6, 1, -115, -59, -95, -102, -121, 84, 65, -108, 92, -42, 2, -109, 118, -54, 89, -17, -71, -61, 54, -71, -2, 109, 56, 24, 54, 13, 44, 103, -108, -32, -4, -20, -82, 30, 123, -119, -81, 69, -56, 85, 69, 93, -25, 104, 5, -105, 20, -88, 4, -23, -96, -18, 77, 30, -109, 52, 2, -107, 97, 80, 85, -11, -4, 121, -87, -80, 8, 16, -111, -39, 29, -36, 54, -54, -90, -56, -87, 73, -27, 115, 42, 64, -102, -116, -76, 113, 91, 79, 35, -8, -86, 36, 24, -100, -108, 7, -1, -113, -94, 94, 105, -43, 124, -70, -30, 41, -101, -67, 90, -68, 86, 6, 124, -119, 67, -24, -85, 107, 105, 29, -89, -2, 18, -16, -32, 80, 78, -74, -67, 47, -41, 107, 67, -35, 34, -126, -112, -19, -52, 18, -92, -126, 1, 75, 10, -55, -80, -95, 16, 107, 49, -45, 54, 74, -54, 101, 3, 34, -84, -55, 73, -82, -95, 53, -21, 124, 11, -8, -2, -107, -108, -49, -59, 89, -70, 41, -52, 82, -109, 105, -97, 30, -77, -105, -91, 13, -15, 41, 3, -117, 5, -66, -124, -21, 42, 117, 91, -61, 105, 59, 60, -1, -98, 16, -12, -26, -115, 26, -124, -68, -76, 42, 112, -10, 60, 54, -80, -1, -51, -32, 32, -66, 61, 95, 79, -116, 61, 55, -106, 33, -7, -87, -124, 117, 79, -48, -70, -29, 108, -44, 107, 77, -87, 38, 49, -66, -78, -114, 18, -84, 113, -82, 102, -73, -82, -123, -89, 10, 56, 68, 85, -9, -10, 82, -28, 97, -98, 38, -26, -74, -96, -103, -8, 16, 3, -93, -85, 34, -1, 74, 92, 78, -54, -91, -100, 50, -109, 29, -28, 106, -119, 63, 92, -128, -9, 17, 10, 12, 14, -56, 10, 96, -26, -17, -87, -5, 28, -13, -42, -61, -30, 34, 34, 25, -39, 71, 23, 79, -104, -123, 1, 43, 23, -47, -79, 108, 122, 93, 29, 66, -23, -90, -114, -5, -51, 101, -25, 97, 119, 79, 42, 112, 69, 104, 13, 122, 78, -120, 98, 57, 116, -82, -82, -17, 119, -53, 94, -39, -65, 79, -77, -71, 8, -90, -82, -92, -67, 31, -114, -92, 46, 86, 47, 118, -13, 65, 30, 55, -40, -30, 99, 3, 77, -99, -115, 113, 8, -87, -26, -28, 117, -16, -99, -98, -80, -46, -70, -7, 101, -109, 87, 96, -46, 81, -71, 30, 9, -59, 95, -2, 79, 25, 81, -103, -102, -86, -20, 14, -87, -126, 106, -127, 88, 30, 83, -71, -77, -86, 107, 65, -114, 105, -71, 25, 98, 68, -57, -42, -79, 127, 123, -12, -39, -125, 108, -6, 123, -113, -36, -29, -27, 25, 7, 83, 59, -123, -119, 43, 71, 45, -103, 97, -79, 75, 124, -17, -84, -96, -51, -26, -83, -37, 61, -100, 73, 80, 75, 0, -74, 2, 99, 97, 98, 110, -33, 38, 122, -79, 12, 102, -34, 48, -30, -8, 23, 59, -30, 48, -62, 90, -48, 9, -103, 120, 126, -30, 21, 67, 121, 97, 91, -89, 48, 51, 0, 112, 96, -99, 85, -15, -14, 103, -17, 96, 49, -117, 78, -91, -15, 103, -16, -127, 89, -4, 45, -51, 57, -13, -2, -40, -31, -29, -83, -14, -107, 11, 65, 86, 17, 26, 16, 0, 62, -117, -21, -116, -106, -66, -25, -11, -81, 103, 117, -127, 6, 7, 29, -25, -58, -42, 120, -110, 45, -98, 124, 36, -116, 104, -119, 104, 106, -63, -116, -121, 67, -8, -113, 3, 103, 84, -120, 104, 76, 54, 91, 9, -38, -106, -28, -55, 24, 116, -43, 33, -100, -1, 34, -17, 45, -38, 82, 61, 110, -83, 109, 98, 77, 0, 36, 125, -68, -30, 57, 61, -49, 90, -60, -110, 101, 22, 28, 37, -72, 45, 10, 95, 39, 117, 8, 15, 5, -84, 10, 68, 49, 34, 92, -10, -75, -88, -86, -5, 42, -16, 5, 43, -31, -32, 0, -126, 39, -114, 88, -34, 124, -112, 1, -112, 22, 60, -126, -42, 90, -90, -3, 39, 115, -39, 112, -16, 62, -32, 117, -92, -80, -112, -98, 12, -112, -81, -10, -13, -3, 57, 67, -26, 12, 83, -22, -46, 110, 12, 49, -55, 75, -94, 119, 97, 0, -52, -107, -128, 118, -86, -120, 63, 44, -105, -114, -113, 40, -111, 113, -35, 47, -11, 16, 106, 124, 36, -94, 85, 3, -87, -95, -77, 2, 53, 1, -61, -24, -105, 5, -10, -55, -57, 72, -39, -85, -36, 66, -73, 127, -2, 72, -10, -120, -71, -43, 103, 122, -77, -126, 86, 77, 3, 89, 3, 18, -43, 122, 35, 9, -31, 2, 29, -56, -108, -82, 12, -86, -116, -35, 72, -57, -2, -113, -115, 19, -45, 43, -9, -118, 94, 84, 56, -26, -33, -119, -18, 67, 8, 18, -61, 19, -79, 118, -107, 6, -94, 59, -120, -21, -86, -27, -86, -52, -88, 3, 106, -29, -75, -81, -59, 36, -71, 98, 45, -109, -27, 76, 117, -69, -12, -93, -84, -127, 37, -35, 112, -87, 24, -32, -26, -121, 57, -123, -64, 63, 74, -82, -62, -81, -120, -123, 89, 50, 103, 65, 92, 0, 46, -105, 72, 17, 88, 66, 53, -128, -96, -29, -50, 12, 110, 120, -115, -80, 45, 64, 42, -10, -16, -63, -83, 117, -104, 111, -45, -63, -4, 56, -93, 9, -93, -80, -7, 113, -81, -78, -82, 119, -5, 33, 21, 122, 124, -103, 97, 71, 24, 25, -37, 29, -64, -33, 41, 75, -42, -57, -109, -120, -109, 111, 25, -127, -84, 51, 103, -123, 16, -25, -122, 76, -67, -4, -88, 93, 53, 105, 105, 57, 24, -75, -120, 7, -38, 8, -13, -106, -50, 88, -105, 34, -83, -120, -89, 1, 114, 93, -123, -107, -34, -63, 58, 62, 115, -61, -101, 101, -30, -50, 50, 50, -35, 32, -107, -77, -26, -33, 0, -5, -9, -76, 107, 29, -21, -6, -80, 40, 93, -5, 100, -57, -65, 50, -23, 89, 63, 95, -63, 13, -9, 117, -32, -80, 21, -103, -109, 18, 106, 27, 70, -36, -66, -91, -74, 43, -72, -96, 55, 81, -85, 96, -16, -123, -32, 92, -19, 125, -68, -97, 108, 74, -8, -84, 113, -15, 34, -32, 6, 13, -120, -52, 75, 62, 57, 90, 81, 39, 27, -89, 45, -30, -41, -40, 59, -11, -86, -19, 48, -53, -67, 87, 28, -75, 3, -92, 3, 61, -107, -45, -71, -113, -55, -97, 71, -27, -54, 118, 91, -66, -87, -57, -62, 37, -50, 78, -77, 15, 3, 60, 21, -117, 68, 98, -1, 56, -51, 60, 48, -62, 113, 108, 17, 4, -37, 118, 121, 8, 42, 105, -116, -23, -55, -64, -29, -121, 95, -4, -51, -89, 100, 77, -117, -124, -91, 124, -101, 81, -57, 21, -28, -81, 72, 90, 61, 109, 55, -36, 117, 54, -15, -102, -68, -6, 105, 77, 22, 81, -13, 51, -74, -123, 48, 100, -30, 47, 22, -102, -89, -33, -79, -71, -76, 8, 127, 117, -70, -2, 60, 27, 0, 107, 18, 15, -108, -37, 53, -61, -101, -56, 9, 59, 19, -62, -52, -98, -59, -65, 106, 65, -40, 68, -53, -107, 100, -102, 101, -124, 8, 62, -13, -29, 103, -100, -95, 108, 72, -80, -29, -61, 116, -55, 22, -62, 52, -33, 61, -124, -37, -112, 27, 58, -31, 26, -76, 79, 46, 81, -34, -19, -127, -77, -123, 123, -102, 108, -73, -88, 125, 114, -91, -80, -55, 24, -10, -58, 56, 92, -50, 9, -21, 27, -113, 109, -117, 62, -84, 119, -28, -13, -68, -46, -69, 116, 11, 107, -83, 52, 37, 29, 80, 59, -99, -35, 114, -92, -63, -64, 97, 60, 75, -101, 85, -5, 65, 8, -48, -22, 91, 7, -116, -31, 91, 105, 85, 62, -93, -127, -63, 59, 77, 90, -63, 113, -44, 1, 61, 18, -13, 10, 104, -41, 23, 10, -43, 124, 43, 28, -125, -78, -4, -119, 68, -33, -55, -108, -27, 112, 101, -95, 86, 81, -115, -106, 101, -53, 92, 112, 77, 13, -8, -100, 26, -78, 123, 56, -113, -85, 79, 112, -4, -116, -72, 62, -48, -6, -99, -83, 108, 108, -34, -85, -87, 110, 92, 11, -108, 29, -120, -108, -123, 81, -28, -102, -66, -15, 89, -55, 102, 23, 117, 107, 123, -56, -95, 72, -18, -35, -31, 108, -128, 81, -89, 90, 89, -113, 84, -48, -125, -79, 115, -23, -76, -105, 25, -28, -84, -107, -85, -56, -121, 80, -99, -86, 15, 102, 1, -8, -65, 13, -23, 28, 105, -39, -8, -81, 22, -35, -52, 74, 102, -56, 98, 30, 100, 121, 101, 79, -106, 103, -103, -114, -20, 107, -11, 127, -28, -63, -41, 124, 127, -105, 1, -13, -83, 33, 60, 13, 43, -7, -40, 49, -87, -94, -32, -41, -93, 70, 25, 76, -8, -23, -22, -8, -16, -39, 88, 93, -13, -27, 17, -20, 72, -81, 14, -117, -55, -48, 51, -66, -59, -36, -25, 58, 6, 99, -33, 98, -2, -81, 61, 23, 107, 127, -102, 94, -26, 101, 7, 55, 54, 119, 28, 19, -105, 29, -95, -53, 76, -107, 92, 33, -106, -104, -48, -106, -72, 101, -116, -79, 57, -43, -77, 19, 57, -42, 96, -126, -109, 86, -3, 86, -55, -97, -69, -17, -34, 19, -122, 85, 49, -96, -23, 40, 65, -10, 120, 97, 43, -86, -35, 44, 118, -32, 33, 100, -26, -50, 65, 56, -60, -41, -98, 127, -111, -40, 81, -67, -106, -7, 123, -35, 3, -121, 104, 22, 11, 31, -11, -84, 81, 104, -69, 35, 99, -4, -108, 2, 67, -116, -50, -19, 98, -6, -55, 33, -32, 5, -122, 7, -4, 95, 3, 73, 90, -81, -16, -122, -7, -12, -67, 65, 94, 43, -21, 49, 69, -84, 32, 126, -36, 106, 109, -89, -102, -68, 45, -50, -94, 3, 75, -8, -24, -79, 124, 88, 126, 93, -49, -95, 64, 115, 54, -89, 30, -76, 110, 81, 104, -11, 127, -123, 44, -128, 74, 62, -93, -70, -62, 63, 80, -119, -43, -27, -57, 63, 67, -19, -72, 0, -88, 100, -128, 41, -29, 42, -41, 86, 85, 108, 96, 89, 72, -122, -121, -10, -30, 57, -33, -125, 31, -100, -30, 37, -90, 94, 0, -16, -26, 103, 77, 6, 107, 104, -34, 61, 6, 60, 87, -65, -88, -37, 87, -20, -105, -3, 8, -11, -49, -26, 1, 46, -17, 13, 49, 93, 62, -50, 70, 72, -34, -7, -18, 88, -126, -49, -108, 113, 122, 19, -29, 97, -32, 29, -2, -119, 90, 22, 37, -9, -28, 62, 30, 63, -97, -118, -12, 48, 50, -71, 46, -115, -123, 83, 63, -79, -50, 75, -56, 94, -30, -76, 34, 96, 89, 30, -71, -59, -50, -51, 45, 76, -100, 46, 122, -40, 39, 71, -103, 36, -121, 78, 112, 9, 108, -90, 81, -116, -63, 52, 119, 32, -51, 35, -110, -22, 65, -125, -89, 14, -4, -52, -28, 117, -116, 87, -106, -92, 71, -21, 26, 93, -103, -40, -71, -4, 41, -55, -97, 23, 1, -90, 123, -57, -11, -89, 36, -82, -31, -38, 127, 109, -45, 46, 114, 115, -89, -32, -3, -112, -65, 73, 51, -77, 60, 99, -118, -111, -88, -58, -88, -73, -16, -71, -79, -54, -63, -126, 50, 20, 96, 69, -60, 31, 81, 84, -70, 25, 7, 121, 82, 73, -65, -9, -120, 95, -106, -8, -18, -5, 41, 51, -72, -108, -88, -36, 107, 99, -24, -122, 109, 125, -105, 73, -96, -95, -125, -44, -119, 83, -10, 50, -82, 13, 42, -76, -2, -40, -37, 100, -66, -46, -123, -22, 60, 74, 97, -107, 88, 87, 13, 11, -90, 75, 46, 77, -100, 115, -13, 84, 114, -99, -54, 127, 41, -68, -35, -43, 83, -27, 80, -92, 51, 68, 84, 77, -76, 36, 30, -83, 17, -123, -109, 14, -31, 70, 94, -46, -112, -68, 63, 48, -4, 107, 26, -16, -39, -48, 118, -36, 61, 65, 24, 7, 26, 14, 12, -51, -76, -27, 36, 87, -46, -30, -13, -67, 121, -69, 29, 40, -13, -19, -72, 32, -61, 19, -71, -52, 1, 89, 51, -78, -48, -19, 76, 7, -73, -112, 117, -98, -101, 118, 78, 9, -125, 59, -93, -101, -92, -105, -91, -65, -24, 62, -26, 8, -94, -17, 105, -57, -50, -77, -118, 117, -14, -118, 110, -124, 95, -88, -41, -104, -101, 7, -41, 2, -24, -106, -126, 36, 82, -97, -81, -26, -32, -34, 115, 16, 15, -37, 13, 3, 79, 104, 75, -32, 79, 127, -100, 22, -58, -48, -60, 88, 28, 41, 26, 116, 15, -108, -55, -59, -9, 96, -58, -61, -40, 111, -103, -22, 34, -53, -42, -126, -87, 25, -73, 106, 102, -89, 77, -54, -72, 76, 67, 24, 67, 122, -23, -40, 9, -41, -42, 93, 109, 32, -30, -92, -23, -77, -82, 17, 2, 114, -122, 28, 102, -39, 49, 114, 49, 109, -28, 118, -8, 19, -12, 121, 101, 66, -98, -30, 86, -3, -39, -82, 126, 12, -5, -13, -5, -38, -12, -120, -75, 36, -118, -25, -43, -84, -83, -77, 57, 92, -8, 27, 102, -61, -109, 39, 85, 50, 122, 9, 102, -109, 73, 38, 90, -82, -94, 98, 28, 59, 106, -33, 98, 53, 107, 75, -125, 12, -48, -53, 16, 48, -110, 74, 122, -23, -114, -125, -5, 113, -114, -69, 33, 71, 108, 107, -104, -51, -111, 66, 28, 124, 114, 17, -46, -1, 67, 106, -27, 49, -22, 103, 15, -76, 17, 76, 84, 85, 60, 61, -123, 45, -32, -60, -21, 2, -128, 81, -19, 17, -111, -120, 22, 65, 112, 74, -102, 63, -81, 24, -47, 123, 99, -123, -4, -118, 11, 106, -94, 114, 54, -14, 60, 30, 54, 34, -70, -8, -82, -92, 63, -93, -34, -72, -86, -10, 69, -103, -72, 104, 84, -105, 83, 26, 122, 28, -127, -49, 52, 115, 42, 30, 23, 78, -36, -32, 42, -5, 123, -47, 92, -83, -92, -118, 57, 18, -31, -78, -33, 62, -23, -8, -33, -75, 89, 106, -74, -101, -61, 13, -126, -66, -106, -119, -114, -75, -50, 105, -70, 40, -51, 74, -4, 31, -4, -33, -54, -18, 1, 5, -35, 24, 52, 113, -123, 6, 95, -35, -89, -82, -54, -81, 87, 16, 107, 72, 13, 4, -121, -4, -87, 53, 48, -104, -85, -67, 22, 43, 72, 72, -34, 51, 49, -1, 105, -103, -126, 53, -50, -34, 17, -93, 53, 13, -112, 39, -44, -55, 117, -110, -108, 122, -124, 47, -82, -109, -113, -15, -54, -73, 105, -115, 40, 61, 23, -82, 103, -37, -50, -75, 20, -50, -27, -106, -89, 26, -96, -46, 9, -83, -25, -78, 127, -34, -81, 62, 114, 85, 92, 98, 93, -55, -125, -29, -104, -44, 117, 48, -95, 56, 87, -98, -62, 50, 120, -36, 57, 96, -125, -15, 24, 0, 100, 61, -13, -110, 43, -52, -10, 66, 18, -90, 48, -110, 97, 58, -116, 2, 103, 74, 66, -84, 44, 17, -111, 116, 71, -104, -12, -53, -121, 83, -44, 96, 39, 63, -30, -56, 103, 54, -108, -50, -51, 105, 86, -41, 46, 52, 55, 83, 26, -108, 48, -25, -11, -68, 63, 16, -125, 38, -49, 45, -28, -119, -68, 61, 108, -88, -21, 33, -117, 77, 57, -10, 69, 55, -128, 41, -95, -117, 83, -123, 56, -102, -48, 15, 113, -42, 40, 120, 100, -89, 43, -41, -112, -87, -124, -67, -48, 75, -27, -119, -42, -68, -44, 11, -82, -55, 79, 37, -80, -28, 58, 23, -74, 9, 13, -94, 118, 13, 80, 102, 86, -14, -78, -110, 61, 116, -104, -81, 37, 103, -118, -78, -65, 73, 122, -63, 116, -86, 120, -17, 82, 69, -125, 97, 11, 41, 62, 61, 13, -81, -9, -62, -101, 35, 67, 119, 22, 5, 127, 68, 18, -79, 49, -50, -31, 40, 120, 66, -46, 117, -24, 122, -48, -116, 74, 120, -106, -96, 6, 53, -74, 80, 36, -35, 29, 12, 6, 111, -87, 31, -26, -42, -60, -66, 124, 0, -57, 69, 97, 126, -63, -92, -106, -92, -29, 71, 82, -39, 80, 86, 122, -9, 15, 114, -53, -61, 19, 88, 15, 42, 110, 11, -96, -68, -116, 34, -20, -52, 104, 22, -102, 85, -125, -16, -107, -79, 62, -96, -70, -38, -82, -51, 33, 47, -84, 26, 112, -97, 81, 85, -128, 40, 69, -55, 104, 116, 41, 105, -83, -79, -66, 50, 46, 106, -118, 99, -31, 55, -123, 107, -20, -48, -44, 117, -81, 30, -92, -97, -102, -114, 38, 40, 27, -115, 15, -18, -42, -55, -20, 49, -14, -94, 2, -5, -114, 111, -128, -17, -108, 61, -58, 79, 32, 79, -126, -20, -34, 51, 35, 89, -97, -121, -25, 88, -116, -30, -13, -14, -62, 42, 77, 99, -94, 71, -1, -113, 99, -7, 10, -20, 20, -65, -5, -79, 114, -86, -5, -122, 117, -23, -5, 96, 127, -126, -119, -31, 8, 12, 80, -47, -41, -77, -37, -43, 107, -9, -38, 80, 43, -127, 15, 92, -76, -49, -15, 83, -47, -70, -88, 5, -35, -104, -10, 126, -56, 117, 24, 30, 1, 41, -83, 122, -13, -42, 60, -87, -34, 81, 90, -55, 3, -43, -128, -8, -76, -7, 7, -17, -77, 57, -20, -81, 74, 16, -88, 87, -36, 8, -31, -49, 114, -81, 16, -28, 110, -13, -18, -9, 4, 34, -70, -31, -79, 80, 30, -28, -80, 83, -106, 38, -71, 28, -117, -128, 109, -19, 121, -124, -5, 55, -6, -92, 115, -123, 29, -31, 96, -82, 124, -98, -4, 96, 9, -81, -67, 100, 55, -32, -18, 122, -9, 0, 30, -44, 55, 56, 29, 70, 6, -91, -83, 54, 84, 38, -102, 90, -91, 122, -24, -65, -72, -102, 39, -41, 98, 32, -33, 13, -3, 8, -127, -66, -94, -95, -53, -72, -50, 6, -90, -28, -89, -124, 71, -90, 93, -6, -74, 2, -114, -128, 4, -57, 6, -53, -122, 93, -36, -117, -73, 76, -44, -56, -68, -105, 123, 8, 33, -48, -43, 11, -100, 41, 3, -127, -23, -121, -96, 71, -127, -12, -82, 74, -50, 43, -25, 83, 79, -9, -41, -128, -58, -96, -21, 1, -49, -40, 4, -125, -120, -81, 29, -105, 2, 65, -105, 112, 46, 117, 53, 102, -124, 39, -109, -60, -39, -104, -95, 79, -108, -96, 117, 50, 118, -63, 16, -31, -26, -101, -39, 95, -50, -8, 90, 77, -18, 92, 114, -102, -60, -24, 57, -60, -8, -67, 78, 66, 122, 62, 49, 104, -76, -38, 97, -59, -87, -73, 60, 26, 19, -15, 68, -36, 6, 13, -22, -57, -1, -123, -106, 106, 59, -127, -88, 41, 21, 80, -62, -107, -54, -106, 99, 64, 50, 8, -8, 13, -83, 76, 75, -75, -99, 44, -96, 38, -81, 84, 46, 86, 70, 92, -10, -42, 14, -70, 0, -112, 8, 115, -20, 4, -121, 20, 9, -3, -76, 10, -14, 103, -38, -2, -66, -43, -53, 37, -2, 32, -3, 51, 53, 41, -119, 122, 113, -98, -73, 83, 16, -10, 73, -105, -53, 41, -54, 63, 108, 20, -51, 81, 17, 21, 45, 125, 81, 59, -58, -99, -1, 109, -70, -103, -107, 70, -85, -37, -117, 98, -10, 10, 44, 76, 116, 72, -84, -38, -84, -47, -106, 70, -103, -84, 98, -75, -67, 26, 75, -94, 16, -65, 44, 30, -7, 113, -64, -53, -31, -126, 106, -93, -93, -109, 100, 67, -13, -127, 9, -45, -109, 8, -11, -21, -29, 56, -113, 76, 105, -41, -104, -55, 3, 1, 89, 102, 69, -101, 68, -68, -100, -8, -25, 8, -15, 7, 78, 4, 107, 89, 42, 31, -93, 17, 118, 102, 44, -59, 55, -111, 7, -114, 5, -23, 27, -128, -78, -123, 64, 45, -15, 42, -34, -64, 122, -39, -14, -94, -2, -37, 18, -41, 37, -80, -47, 23, -117, 82, -125, 59, 102, -121, 100, -124, -109, 24, -104, 102, 71, -79, 47, 102, -79, 73, -86, -90, 58, 41, -78, 112, 86, -58, -69, -17, 110, 29, 26, -61, -121, 67, 35, 93, 72, 7, 19, -116, 20, -69, 119, -44, -55, -61, -58, -66, 94, -124, 110, 25, -100, 105, -97, -77, 16, 89, -12, 111, -29, -25, 88, -23, -56, 14, -47, 39, -101, 3, -28, -2, -116, 59, 54, 99, -35, -32, 23, 60, 67, 123, 76, -126, -42, -118, 115, -90, 110, 86, 46, -128, -77, 71, -115, -85, -23, 2, 60, 88, -18, 44, 43, 27, -117, -32, 74, -126, 26, 63, -22, -109, 84, 94, 112, -110, 7, -55, -4, 46, 83, 98, -6, 98, -38, 8, -30, -44, 55, -80, 80, 90, 27, -80, 6, 41, 71, -93, 55, -114, -41, -105, 51, -9, -3, 107, -67, -29, -48, 61, 74, -71, -128, -31, 12, 72, 29, 94, 18, 124, -128, -128, 115, 68, 31, -57, 84, 56, 55, 44, 68, -54, -25, -50, 24, -122, -95, -86, 18, 70, -115, -52, 3, -73, 74, 55, 37, 122, -70, 113, 40, -2, 82, -64, 80, -85, -108, -5, -94, -118, -3, 84, 88, -29, -83, 58, 0, -103, -6, -107, -22, -63, -94, -34, -127, 26, 45, -107, -116, 15, 30, 123, -89, 74, 110, 127, 11, 93, -119, -2, 64, -24, 69, 80, 23, 122, 114, 46, -50, 31, -9, -68, 40, 86, 84, -36, 114, 92, 81, -124, -35, 31, 54, -110, 47, 21, -46, 74, -94, 65, -116, -2, 46, -68, 50, -119, -105, -34, -60, -57, 65, -23, -82, 20, -21, 106, 90, -40, -38, -76, 37, 118, -41, 114, -91, -34, -6, 105, 51, -17, 11, -4, 30, 79, 44, 95, -126, 83, -48, -80, -115, 47, 69, -20, -119, 57, 126, -73, 82, 3, -107, 38, 53, -12, 122, -113, -56, 126, -82, -109, 1, -10, 0, 54, 119, 26, -34, 84, -6, -41, 98, -70, -34, 59, -122, -98, -33, -3, -82, 43, -71, -104, 38, -8, -85, -32, 29, -3, 17, -40, -60, 55, 84, -73, -9, 91, 21, -23, 72, 117, -3, 119, 13, 62, 62, 64, -64, 18, -44, -42, 94, -121, -37, 15, 74, -94, -24, 107, 82, -22, -33, -77, -61, 84, 0, -95, 125, 121, 77, 125, 77, 13, -26, 24, -103, -88, -18, 70, 13, 84, -82, 33, 110, 123, -8, -90, -94, -15, -34, 39, -47, -57, -107, 103, 85, 20, 48, -22, -55, -45, -51, 22, 76, -37, 89, -127, 109, -69, -73, 52, 65, -29, 50, 1, 16, -80, 109, 116, -45, -38, 19, 127, -76, 81, -120, 74, 31, -27, -39, -48, -39, -124, -40, 31, -92, 31, 115, -111, -9, 26, 34, -94, 87, -90, 105, -46, 74, 25, 22, 40, 89, 1, -3, 59, 6, -56, 80, -1, -109, -87, 47, 60, -45, 35, 72, -29, 32, -4, -44, -11, 69, -69, -125, 32, 26, -1, -79, -40, 74, 108, -50, -79, 83, 11, -14, 110, -127, 36, 50, -60, -109, -39, 102, 112, 4, 115, 19, 99, -29, 2, 17, -89, 29, 77, -112, 58, 116, 94, -123, -14, -38, 105, -10, -6, -99, 109, -61, -53, 45, 51, 66, 113, -99, 70, 23, 103, 13, 102, 122, -66, 86, 74, 120, -79, -16, -48, 106, 123, 92, 57, 71, 87, -92, -96, 18, 121, -80, 95, -12, -12, -54, -35, 10, 34, 116, -74, 5, -15, 100, 89, 68, -66, 106, 1, 85, -106, -51, -121, 117, 120, -123, -32, -87, 67, 44, 9, -30, 62, -18, -118, 18, -50, -76, 103, 10, -72, 20, -28, -73, -115, 96, -33, 120, 37, 58, 95, 117, -64, -56, -53, -16, -104, -71, 44, 113, -20, -115, 119, 98, -55, -78, -6, 30, 97, 8, 100, -30, 80, 15, -105, 116, 31, 45, -40, 80, 32, -12, 61, 81, 103, 77, 120, -115, -10, -77, 115, 23, -71, 0, 30, -7, -66, 104, -38, 69, 11, -30, 54, 117, -13, -7, -47, 82, -103, -37, -89, 90, -53, 108, -31, -68, 65, -32, -23, -26, -120, -57, -26, 87, 99, 86, 111, -103, 102, -38, -126, 35, -26, 13, -17, 99, 42, -41, 28, 12, -73, -109, -53, 73, -2, -32, -69, 25, -102, -25, 7, -119, 121, -87, -125, -63, 3, 60, 116, 125, -128, 46, -58, -67, -7, 108, -22, 50, 104, 83, 76, -30, -105, -70, 64, -112, 99, -85, 97, -16, -52, 34, -51, -97, 40, -51, -14, -50, 49, -120, 85, -119, -25, 45, 15, 43, -116, 88, -46, 83, -38, -29, -88, 127, 19, -29, -1, 99, 91, 41, -113, 9, -46, -96, 88, -54, 71, -1, 43, 87, 54, -67, -45, -106, 76, 69, -83, 33, 113, 36, -80, -92, 67, 10, 87, -128, 114, -83, 95, 100, -111, -34, 75, 36, -11, -93, -105, 22, -84, -71, 3, -50, -84, -93, -28, -108, -117, -1, -127, 70, -34, -35, 1, -85, -18, -63, -6, -30, -114, 51, -10, 109, -73, -23, -117, -105, 113, 75, -34, 94, -37, -77, 18, 56, 51, 86, -36, -94, 83, 31, 10, -76, 43, -39, -127, -119, -27, 42, -11, 50, -10, 123, 93, -109, 52, 81, 90, -7, 100, -107, -34, -68, -38, -109, 53, 61, 60, 127, 9, -111, 39, -49, -14, -86, 108, -115, 47, -4, 12, 82, 126, -33, 93, 114, 103, -56, -17, 29, 79, 31, 8, -82, 127, 9, -1, 39, 117, -122, 96, -105, -41, -75, -21, -68, -102, 35, -67, -71, 49, -20, 79, 32, 110, -63, 5, -22, 21, -96, 32, -114, -106, 79, 69, -102, 15, 98, -1, 115, 51, -81, 17, -127, 90, -65, 13, 127, -108, 95, 72, 33, -8, -72, 100, -74, -52, -73, 23, -93, 34, -102, 84, 118, 19, -54, -57, -97, 99, 92, 41, 92, -37, 43, -119, 122, 120, -122, 126, -26, -32, -43, -105, -36, -37, -74, -8, -40, 97, -15, -60, 59, -118, -106, -43, 124, -97, 48, 90, -58, -107, -7, -103, 113, -103, -18, 71, 48, 27, -128, 15, -99, -79, 70, 46, -100, 66, -61, 122, -15, 122, -45, -103, -6, 91, -24, -117, -5, -51, 118, 31, 44, 85, -91, 44, 109, -23, 117, -39, -27, 52, -91, 120, 12, 9, 4, -101, 14, -2, 84, 24, -65, 19, 31, -41, -86, -27, -72, 47, 84, -15, -30, 38, 111, 42, 62, -30, 93, 123, -72, -89, 0, -97, 124, 36, -47, -97, -87, -2, -85, 109, -14, -54, 14, -37, -64, -27, 111, -42, -8, 124, 41, -33, -43, -23, 65, -95, -22, 114, -50, 6, -84, 3, 76, -123, 62, 111, -55, -51, -35, -4, 74, 17, -116, 13, 108, 43, -82, 30, -2, -116, -65, -92, -45, -98, 89, 71, -9, -39, -107, 91, -48, 90, -69, 45, -92, -78, -88, 120, 127, 33, 30, 48, -126, 105, -114, 78, -86, -28, 107, 76, 113, -20, 15, -69, 52, -32, 99, -73, 52, -3, 113, -64, -63, 12, -35, 35, 33, 70, 68, -91, -105, -110, 77, -62, -23, -12, -112, -52, 53, 102, 58, -122, 50, -110, -125, -38, -65, -98, 41, -96, -103, -28, -97, -22, -6, 101, 14, 127, -81, -6, -122, -3, 19, -98, -25, 74, 51, 96, -101, 62, 114, -98, -83, -58, -93, -32, 49, 5, -68, -102, 1, 114, 31, -108, -121, -80, 7, 126, 43, 51, 110, -40, -49, -113, -55, -32, -85, -42, -43, 76, 105, 71, 53, 116, 25, 55, -84, 18, 73, -4, 21, 124, -23, 49, -5, 108, 113, -91, -128, -78, -31, -74, 14, -86, -58, -106, -47, -22, 117, -117, -59, -101, 5, -121, 14, -98, 111, -39, -22, 83, -48, -92, -96, 84, -44, -55, -88, 46, 125, 99, -41, -85, 43, -128, 68, 38, 36, -91, -116, -63, -44, 83, -114, -111, -49, -102, -109, 92, -82, -120, 26, 69, 34, -10, 58, 43, 124, 97, 61, -1, -88, -54, 112, 58, 29, 90, -14, -44, -65, 96, -53, -18, 107, 47, -125, 86, 2, -76, 72, 28, -107, -61, 57, 115, -116, -72, -13, 109, 38, 60, 41, -32, 110, 94, -23, -24, 64, -83, -127, 45, 112, 49, -89, -104, -92, 1, 89, -19, 118, 19, 16, -68, -34, 119, 66, 111, -24, 94, 21, 49, -29, -25, 66, 117, -98, 81, 10, -94, 89, -48, 55, -125, -61, -37, -124, -56, -57, 22, 60, -39, -43, 69, -2, 18, -115, 79, 106, -86, 33, -123, 87, -58, -70, -7, -26, 30, 121, 103, 36, 77, -61, 101, 104, -127, 28, 5, 120, 35, -67, 43, 120, 5, 80, 113, 51, 73, 60, -31, 73, -97, -33, 91, -106, -98, 10, 35, 90, -37, 17, 4, -45, 18, 101, 106, 17, -13, -76, -93, 19, 122, -47, -58, -39, -20, -20, 96, -78, -118, -6, -93, -38, -85, 15, -57, 32, -90, 83, 8, -6, -53, -96, 21, -12, -32, -12, 64, 100, 87, 96, 9, 76, 19, -85, 67, 75, 56, -119, -2, -117, 53, 22, -73, 7, 24, 55, 37, -86, -7, -49, -73, -64, -88, -73, -35, -78, -73, 41, 88, -118, 76, 106, 81, 101, 5, 0, 93, 63, -50, -8, -23, -68, -120, 64, -69, -6, -17, 19, -25, -30, -21, -11, -61, 28, 16, -88, 108, -37, 25, -122, 82, -122, 19, -48, 29, -31, -118, -84, -119, -15, 116, 119, -15, -106, -92, 67, 124, -42, -87, 2, -113, -3, -116, 39, -120, -17, -7, 45, -119, 98, -103, -34, 38, -89, 74, -24, -127, 51, 84, -96, -108, 16, 101, -34, -117, 11, 4, -40, 23, 1, 7, 74, -37, -65, 4, 41, 66, -67, -62, 112, 108, 113, 20, 80, -123, 106, 112, -120, 31, 7, 118, -112, 8, -122, -84, 103, 32, -104, -13, -14, 113, -7, 100, -87, -84, 8, -104, -33, -46, 28, 4, -31, -105, 61, -37, 119, -104, 46, -21, 16, 102, -117, 1, 12, -102, -97, -2, -60, -78, 66, -27, -42, 24, 30, -68, 67, -48, 22, 68, 31, 59, 16, -72, -8, -57, -77, 121, -77, -91, -76, 70, 4, -52, 122, 49, 3, -76, -112, 94, 24, -88, -102, -108, 106, -28, 108, -12, 14, 125, -114, -59, 60, 35, -107, 4, 12, -37, -58, 122, 16, 51, 119, -119, 86, 58, 75, 115, 72, -36, 5, 28, 120, 59, -111, -119, -34, -117, -102, -46, 36, -74, -62, -63, 99, -64, -108, 34, 5, -53, -82, -38, -22, -55, -1, 92, -69, 13, -11, -79, -66, -17, -77, 13, 5, 103, -102, 112, 51, 99, -24, 21, 0, 127, -25, -87, -72, -26, -96, -66, -124, 110, -121, 119, -40, 84, 63, -62, 117, 72, -64, -68, -100, -18, 81, 126, 76, 106, -53, 81, -77, 50, -112, 81, -71, -123, 77, -67, 109, 18, -18, -8, 102, -106, 88, -83, -105, 70, 52, -96, 4, 58, 34, -86, -87, 69, 49, 90, -114, -112, 85, -17, 27, 24, 78, 67, -46, 116, -54, 76, -76, 120, -74, -73, -15, -87, -112, -112, -87, -2, 72, -108, 44, -79, 96, -56, -29, 90, 113, -10, -65, 92, 3, -53, 51, 48, 105, 67, -51, -123, -109, 23, -128, -114, 98, 60, 46, -95, -107, -97, -64, -121, 45, 61, 119, -52, 10, -74, -99, -127, 123, -29, -72, 91, 76, -32, -7, -100, -40, 78, -128, 109, 74, -114, 115, -35, 61, 104, 17, -49, 95, 54, 100, -42, 48, 122, 6, 77, 42, 78, -82, -45, -102, -41, 94, -75, 102, -71, -107, -101, 21, -2, -55, 12, -90, -75, 90, -124, -120, -34, -24, -56, 9, 101, 8, 42, -112, 48, 62, 6, -74, -68, 60, -75, -50, 98, 88, 41, 92, 98, 3, 87, -117, 26, -57, 42, 15, -113, 6, 83, -65, -66, -62, -30, 94, 31, -102, -102, 108, -107, 73, -18, -63, 6, -53, -125, -96, -12, 32, -109, -48, -24, 81, 17, 67, 123, 25, -53, -20, 70, 67, 58, 103, -101, 91, -16, 14, -32, 60, 20, 53, -69, -118, -8, -14, -13, 19, 110, -55, -36, 20, -9, -52, -32, -99, 44, 50, 57, -26, 67, 62, 40, 45, 51, -8, -118, -48, 64, 17, 98, 8, -61, 94, -102, 53, -9, -22, 117, -68, -21, -79, 88, 14, 95, -69, -49, -68, 94, -13, -35, 40, 47, -119, -53, 95, -87, 108, -16, 26, -118, 111, 0, 124, -66, 3, -76, 94, -93, 5, 30, 26, -50, 93, -105, -4, -101, -42, -115, 114, 96, -44, -64, 93, -20, -42, 9, -1, 90, -88, -1, -102, 103, -44, -115, -52, -26, -79, -98, 25, 107, 66, -17, -106, -111, -30, -63, -91, -121, -97, 107, -117, 97, 48, -48, 60, -13, 4, -67, -55, -17, 84, 89, -115, 69, -120, -7, -125, 52, -112, 38, -100, -98, 49, 112, 66, 69, 100, 84, -64, -52, -63, 127, -106, 101, 64, 83, -33, 116, 122, -69, 105, -54, 107, -25, -12, 1, 88, -116, 114, -92, 11, -65, 80, -34, -100, -118, 85, -25, -83, 105, -6, 35, -25, -10, 107, 62, 115, -20, -64, 67, 94, -18, -101, -95, 6, 119, 125, 109, -58, 96, 51, 35, 92, -118, 7, -12, 84, -85, -73, 127, -101, -9, 114, -109, -97, 29, 41, 83, -115, -79, -109, -63, 106, 65, 34, -77, 64, 78, 102, 66, -68, -73, -63, 99, 2, -81, 125, 17, 13, -8, -87, -75, -92, -125, -111, -115, -69, -116, -54, -110, 28, -36, -80, 54, -20, 49, 7, 103, -104, -26, -52, -2, 126, 95, 21, -96, 23, 74, -111, 36, -50, 108, -90, -25, -106, 82, 25, 86, -39, 113, 64, -19, 95, 54, 38, -53, -77, -63, -13, -15, -77, 24, 16, -54, 94, 15, 71, 61, 88, 75, 35, 57, -70, -3, -52, 94, -5, 84, -111, -76, -48, -73, 54, 34, -117, 46, 36, -92, -45, -11, 123, -94, -47, -82, 7, -126, 99, -62, -10, -17, -108, 23, 45, 86, -107, 55, 9, -43, 15, 18, 0, -77 );
    signal scenario_output : scenario_type :=( -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 88, 5, -128, -128, -128, -128, 47, 43, 26, 127, -128, 15, 127, -128, -114, -90, -128, -128, -128, -128, -128, -128, -128, -128, 37, 127, 127, 127, -103, 127, -72, -128, -117, -83, 127, 127, 127, 127, 127, -128, -15, 123, 57, 127, 10, 127, -128, -65, -128, -119, -128, 112, 127, 127, 127, 127, -73, -54, 127, 80, 127, 127, -74, 127, -128, 127, 71, -128, 127, 48, 127, 127, 127, 82, -128, -26, -46, 127, -82, -19, 42, -128, -41, -128, -75, 127, -128, 127, -128, 127, -87, 127, 127, -128, 127, -128, 127, 69, 127, 76, 127, -128, 127, -128, 127, 30, -60, 127, -128, 127, 13, 127, 127, 127, 127, 127, -128, -31, -128, 127, 63, 127, 127, -128, 127, -128, 127, -128, 30, -128, 28, 71, 127, 127, -110, 127, -128, 127, -128, -12, -46, -128, 127, -128, -96, -12, 10, -128, 120, -56, -9, -30, -128, -94, -128, -30, 90, -75, -128, -128, -128, -128, 9, 127, -128, 127, -40, 127, 80, 127, 127, 127, -48, -47, -128, -128, -128, -128, 127, -119, 127, -128, -85, -128, -18, -128, 86, 127, -128, -54, -128, -128, -128, 127, 119, 127, -28, 80, -23, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 53, 54, -128, -96, -128, 70, 58, 127, 127, 127, -116, -128, 127, -128, -46, -128, -24, -114, 108, 127, -86, 127, -128, 102, -128, -108, 127, 47, -25, 127, 11, 127, -128, 106, -128, -128, -128, -123, 127, -128, 73, -128, -128, -128, -128, 81, 54, 127, 63, 127, -52, -124, 127, -128, 127, -128, 127, -128, -128, 90, -70, -15, 127, -128, 127, -128, 127, 24, 127, 127, 127, 49, 127, -40, -128, 55, -128, 127, -128, 127, -30, -112, 127, -25, -119, 102, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 102, 127, 127, 127, 127, 127, -54, 12, -128, -128, -128, -128, -128, 127, -128, 127, 98, -8, 127, -128, -77, -128, -15, -128, 91, -128, 24, -128, -128, -128, -128, -128, -128, -92, -30, 127, 127, 127, 127, -128, 90, 6, -128, 127, 127, 127, 127, 127, 110, 127, 127, -128, 127, -92, -128, 51, -68, 127, 40, 127, 127, 127, 127, 127, 127, 127, -93, 127, -128, -128, -128, -128, 127, -128, 127, -128, 98, -128, -128, -128, -128, 58, 127, -128, 127, -128, 127, -86, 127, 104, -128, 63, 18, 127, 127, 127, 99, -128, -128, -128, 127, 53, 127, 9, -123, -128, -128, -128, 117, -128, 127, -128, -34, -128, -128, -128, 123, 80, 127, -10, 127, 55, 51, 6, -4, -128, 127, 34, 127, 127, 127, 127, 22, 76, 127, -128, 127, 93, 127, 127, 127, 127, 53, -128, -128, -128, -128, -116, 127, 127, 127, 127, -128, 127, 127, -28, 127, 86, 127, 127, 127, 127, 127, 127, 51, 127, -128, 127, -128, 54, -47, 127, 127, 127, 127, 127, -18, 127, -21, -86, 35, -128, -54, 51, -34, 127, 127, 103, 127, -128, 20, -128, -128, 20, -128, 127, 127, 127, 127, 127, -72, -128, -128, -128, -128, -44, 127, -112, 127, -128, -124, -128, 127, 122, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -22, -122, -128, -79, -128, -128, -128, -112, -128, -110, 86, 127, 127, 127, 127, 127, 127, 127, -36, 127, 127, 127, 127, -78, -128, -128, -128, -25, -53, 127, 127, -78, 127, 127, 127, 127, -128, -45, -128, -42, -128, -128, 103, -128, 127, -128, 127, -128, 127, 19, -128, -31, 121, -128, 56, -99, 127, -128, 127, -21, 39, -57, -128, 6, 114, -108, 109, -128, -93, -128, -128, -128, 127, 116, 127, 127, 89, 85, -128, -63, -128, -120, 127, 127, 127, -126, 127, 44, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 25, -105, 127, 59, 127, 127, 109, 26, 127, -80, 127, 52, -64, 35, -44, 127, 28, 127, -57, 127, -128, -128, -128, -128, -62, 127, 127, 127, 127, 124, 127, 127, 91, 127, -86, 127, 127, 127, 127, -128, 103, -128, -128, 19, -38, 8, -128, -128, 100, 127, 40, 127, 127, -128, 97, -49, -124, 27, -20, -77, 127, -128, 108, -128, -128, 113, -128, 127, 127, -8, -14, -128, -128, -35, -64, 127, 127, 89, 127, 127, -76, -128, -128, -128, -128, -35, 127, -128, 127, -128, -107, -128, 51, -128, 63, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 3, -102, -39, -128, -128, 92, 127, 127, -128, 127, -128, 127, 127, 127, 127, -113, 127, 100, 127, 127, 127, 127, -128, 66, 120, 7, 127, -39, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 1, 127, -128, -128, -128, -128, -128, -56, -128, 90, 127, -66, 127, -122, 127, -128, -128, 127, 48, 127, 127, 127, 127, 127, -105, 119, -68, -128, -128, -128, -128, -128, -128, 127, 48, 127, -128, 127, -128, -60, 127, 127, 127, -128, -48, -128, -128, -128, -128, -27, -36, 127, 127, 127, 127, 127, -77, 127, -128, 127, -106, 127, 127, 127, 127, 127, 127, 127, 127, 127, 18, -128, 127, -128, 127, -128, -128, 124, -128, 47, 127, 91, 127, -121, 127, -30, -128, -128, -128, -128, -128, 117, 127, 114, 127, 127, -15, 127, 96, -95, 127, -128, 59, -128, -46, 127, 127, 55, 27, -86, -128, -128, 127, -128, 127, -128, 75, -128, -128, 6, -128, -128, -71, -128, -128, -124, 105, 127, 127, 127, 127, 127, 127, -104, 36, -128, -128, -19, -128, -47, 127, -128, 127, -128, 127, -100, 127, 59, -128, -128, -128, -128, -1, 127, 127, 127, 127, 97, 127, 127, 127, 127, 36, -74, -128, -128, -128, -78, -128, -64, -128, -128, -128, 38, -128, 127, -14, 127, -26, 127, 30, -128, -128, -128, -128, -128, -128, -128, -128, -128, 74, 127, 98, 127, 127, 125, 127, -128, 127, -75, 127, 127, -128, 127, -128, -128, 14, -128, 127, -97, -4, -128, 75, -128, 64, -128, 127, -128, 127, -28, 127, -128, 113, -128, 56, 127, -128, -128, -128, -128, -128, -128, -70, 127, -3, 127, 127, 116, 127, 127, 127, -113, -66, 27, -128, 127, -128, 70, 13, -106, 127, -87, 127, -128, -10, -27, 96, 127, 127, 127, 127, -128, -77, -128, 123, -60, -128, -70, -128, -128, -128, -128, 102, 127, 127, 127, 127, 127, -17, 127, -55, 127, -3, -128, -125, -128, -128, -128, 29, 127, 127, 127, 127, 127, 127, -32, -128, -128, -128, -42, -128, -43, -44, 127, 127, 127, 127, -128, -9, 35, 7, 127, 127, 127, 63, 45, -38, -87, 47, -128, 14, -70, 14, -128, 127, -128, 127, -128, -128, -128, 38, -128, -128, -128, -128, -40, -38, 41, 127, -80, 127, 127, 28, 127, 102, 127, 124, -128, -128, -128, -128, 0, 110, 127, 127, 127, 28, -128, -128, -128, -128, -128, -128, -128, -42, 127, 63, 127, 127, 127, 127, -128, -128, -21, -128, 127, -105, 77, 127, -128, 27, -128, 58, -37, -54, -128, 127, -128, 127, -128, -98, 124, -47, 97, 127, 127, 127, -128, -18, -128, -128, 127, -128, 127, 10, 127, 127, -27, 127, -91, 115, 52, 96, 127, 127, 127, 42, 76, -77, 30, -128, -128, -128, -128, -70, -13, 28, -99, -89, -128, 127, -128, -128, -128, -128, -128, -120, 127, 1, 127, -128, -128, 91, -128, 127, -38, 26, 127, -83, 127, 87, -53, 127, -128, -2, -128, -128, -128, 127, -5, 127, 113, 127, 127, 127, 127, 127, 127, -53, 77, -128, -48, -128, -128, -82, -100, -128, -128, -128, -128, -94, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 47, -128, 127, 127, 127, 127, 127, 30, 127, -43, 127, -62, 28, -128, 60, -128, -128, 0, 127, 127, 127, 127, -128, -128, -128, -128, -34, -52, -122, -128, -128, 127, -128, 127, -80, 127, 127, -128, 127, -128, 127, -128, 87, -128, -128, 127, 127, 127, 1, 30, -128, 11, -43, -128, 127, -128, -61, -54, -128, -128, -128, -128, -128, 59, -128, 7, 127, -7, 127, -27, -128, -128, -128, -128, -99, -128, 37, 69, -128, 127, -91, 127, -128, -53, 5, -128, -71, -128, -128, -91, -128, -128, -128, -128, 46, 112, 127, 127, -128, 127, 97, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -121, -103, 99, -111, -127, -128, -128, -72, -128, -4, -128, -35, 109, -64, 127, -128, 127, -31, 127, 22, -128, -128, -128, -128, 127, -128, 127, -128, -30, -128, -30, -12, -128, 127, -128, 127, -107, 115, 127, -128, 127, -128, 127, 127, 69, 127, 127, 127, 97, 127, 127, 61, 127, -128, 21, -128, 127, 127, 127, 127, -128, -128, -128, -128, 46, -7, 127, -128, -5, -128, -128, -128, -128, 127, -128, 127, 121, 65, 127, 53, 127, -128, -128, -128, -128, -128, 75, 127, 6, 100, -128, 127, -128, -128, -128, -73, 127, 1, -128, 32, -128, -58, -128, -39, 127, -40, 127, 75, 127, 127, 127, 127, 127, 127, 36, -128, -128, -128, 127, -128, 127, -128, -76, -128, -128, 56, -98, 77, -128, -128, -128, -128, 127, 5, 127, 123, -111, -8, -107, -128, -128, 127, 127, 127, 127, 127, 127, -59, -128, 127, -128, -69, -37, -128, 14, -128, 109, -128, -128, -128, 127, 61, 127, 127, 102, -128, -128, -128, -53, 127, 127, 127, 127, 127, 60, -128, 95, -128, -8, -128, 2, 127, -12, 127, 127, -128, 104, -128, 127, 127, 5, 127, 127, 127, 127, -128, 127, -128, 127, 127, -64, 127, -7, -128, 64, 58, 13, 26, -28, -128, 114, 42, -128, 103, -128, 127, -43, -19, 93, -128, -128, -128, -128, 122, -128, -8, -128, -128, 127, -128, 35, 127, -9, -128, -128, -128, -128, -128, -128, -128, -13, -128, -75, -114, -128, -128, -128, -128, -128, -128, -128, 127, -128, 83, 76, 114, -128, -128, 74, -128, -128, -128, 80, -128, -128, -128, -128, 99, -128, -75, 127, -128, 127, -111, 127, 127, 38, 76, 127, -128, -128, -128, 68, 31, -128, -128, -88, -128, -31, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, 106, -48, 127, -128, 127, -128, 127, 127, 15, 127, 127, 127, -123, 127, 127, 127, 127, 127, 71, -128, 54, -128, 127, 127, 127, 127, 127, 127, 127, 127, 24, -128, -128, -128, 127, 45, 20, -64, -128, 21, -128, 127, 127, 106, 127, -128, 45, -128, 127, 127, 127, -89, 42, -128, -128, -128, -128, 90, 8, 127, 127, 127, 127, 127, 127, 61, 98, 127, -24, 127, 72, -108, -128, -23, -128, -128, -128, 54, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 78, -57, -128, 127, 127, 127, 127, 127, 127, 127, 28, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 122, 58, -60, 127, 123, 127, 69, 92, -128, -128, -128, -128, -32, -128, 127, 127, -114, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -62, -128, -121, -128, -128, 127, -128, 127, -128, 48, 127, -128, 0, -128, -73, -128, 72, -128, -128, -128, -128, 80, 127, 127, 5, 127, -9, -128, 127, -128, -128, -128, -128, -128, -128, -122, -128, -128, -128, 32, -119, 12, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, -80, 127, 127, 127, -128, 127, -128, -128, -86, -128, 127, 19, 127, 127, 127, 127, 42, 122, 52, 97, 127, 27, 127, 43, 96, 19, 21, 110, 56, -128, -128, -128, -128, 127, -128, -111, 46, -128, 7, 127, -112, 4, -90, 73, 2, 72, 127, -128, 91, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -116, -19, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -27, 127, 127, 18, 127, 4, 127, 127, 18, 127, -128, -128, -12, -128, 127, 0, 127, 37, 7, -128, -25, -128, -89, -128, 127, 127, 127, 127, -128, -113, -128, -128, -128, -128, 28, -128, -128, -128, -128, -128, -128, -128, -49, 59, -128, -128, -128, -128, -128, 74, 17, 127, 127, -128, 57, 125, -128, 127, -51, 127, 127, -45, -128, -128, -128, -128, -96, 25, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, 89, 27, 127, -128, -128, -128, -128, -128, -128, -128, -128, 56, -128, 127, -128, -68, 127, 127, 127, 127, 22, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 37, -78, 127, -128, -82, 78, -128, 127, -120, 127, 27, 127, 127, -76, 65, 127, -38, 127, 127, -128, -60, -72, -20, 127, 8, 127, 96, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 94, -128, 102, -128, 63, -128, -128, -128, -128, -128, 85, 127, 127, -36, -128, 127, -128, 127, -128, 127, -113, -48, -48, 119, -47, -128, 2, -86, -61, 58, 127, 127, 114, -122, 127, -128, 127, 99, 127, 127, -38, -128, -62, -89, 127, 127, 127, -81, -128, -128, -128, 127, 127, 127, 127, 127, 127, 104, 127, 127, -128, -128, -128, -128, -128, -128, -126, 127, -128, 127, -128, 127, -128, 17, -59, -128, 127, -128, 127, -128, 127, -18, 127, 127, -86, -128, -128, -128, 44, 127, -128, 127, -128, -97, -128, -41, 127, 127, 127, -39, -1, 90, -128, 127, -128, -128, -128, -128, 127, -128, 127, 36, 127, 127, -40, 127, -128, -128, -128, -10, -128, -102, -128, 2, -128, -128, 127, 127, 127, 93, 34, -128, -128, -128, -128, -119, 127, 53, 127, -128, 127, -128, 14, -18, 127, -51, 9, 127, 66, 127, 127, 127, 120, 127, 99, -128, 105, -88, 127, 127, 127, 93, 127, 106, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -126, -128, -128, -128, -128, 65, -128, 127, -20, -128, 127, -42, 49, 127, -57, -55, -128, -116, -128, 127, -128, 127, 127, -122, 127, -128, -128, -128, -128, 113, 127, 127, 127, 127, 114, -51, 127, -128, 127, -128, 76, -128, 47, -128, 27, 127, 127, 127, 127, 127, 127, -10, 127, 127, -56, 77, -128, -128, -128, 74, -65, -104, 127, 76, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -117, -128, 127, -128, 127, 39, -43, -128, -128, -128, 64, -128, 17, -128, 41, -37, -128, 47, -128, -77, -47, -27, 109, 127, -128, 26, -26, -128, -37, -21, 106, 127, -55, -128, 127, -17, 127, 127, -29, 127, 127, -128, 127, -109, -128, 127, -2, 127, 127, -128, -85, -128, 127, -77, 127, -128, 54, -128, -34, -128, 127, 124, 127, -128, 64, -128, 48, -116, -46, 127, -100, 127, -69, 127, -128, 127, -128, 127, -80, 127, 127, -128, -63, -128, -128, -128, -128, -42, -128, -109, -128, -128, -128, -128, 127, 121, -58, 127, -128, 127, -128, 40, 127, -11, -128, 127, -128, -128, -128, 127, 88, 127, 127, 127, 127, -128, 127, 10, 3, -39, -128, -128, -128, 127, -15, 127, 127, 127, 110, 82, -128, 127, -128, 127, -128, 90, -128, -128, -128, -128, -128, -128, -128, -128, -78, 86, 127, 127, 127, -93, 127, -96, -108, 127, 9, 127, -58, -128, -128, -128, -37, 127, 127, 106, 51, -128, -128, -128, -128, 127, 127, 127, 127, -5, -128, -128, -123, 107, -6, 127, 127, -121, 127, 49, 127, -128, 30, -128, -128, -119, -3, 127, 127, 127, -81, 127, -128, 127, -128, 127, -60, 127, 127, 127, 127, 127, 87, -128, -128, -128, -128, -92, 127, 91, -79, -128, -128, -128, -43, -128, -76, -128, -128, 73, 127, -29, 127, -128, 127, 127, 127, 127, 20, 127, 127, -46, 91, 18, 127, 127, -21, 127, -128, 127, 96, 100, 127, -128, -83, -128, -128, -96, -128, 127, -128, -86, -128, -128, 127, -99, 127, 127, 64, 127, -128, 6, -128, -128, -20, -128, 127, 95, 127, 127, 127, 127, 52, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 0, 127, -42, 4, 26, 127, 12, 127, -128, 127, -128, -128, 121, 127, 127, 127, 48, -14, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -97, -128, -128, 127, -128, 127, 55, 13, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 66, 42, -25, 54, -73, 127, 127, 127, 127, -3, 75, -128, -128, -128, 127, 92, 127, 127, 82, 127, -51, -43, -128, -128, -128, -128, -128, 127, 127, 127, 127, 110, 127, -128, 77, -128, -128, -128, -128, 40, -128, -128, 127, -128, 127, -128, 127, -128, -117, -128, -128, -128, 127, 17, 127, 127, -123, 127, 46, 127, 127, 127, 127, 127, -40, -128, -128, -128, -120, -99, -12, 123, -34, -68, -128, -128, -128, -128, -128, -128, -128, -125, -128, -83, -128, 89, -128, -19, 90, 36, 127, 127, 127, 127, 105, -128, -128, -128, -128, -71, -91, 102, -95, 127, 35, 127, 89, 127, 127, 127, 127, 127, 127, 49, 41, -128, -128, -128, -128, -124, 31, -128, -128, 127, -128, 127, -45, 127, 17, -128, -128, -128, -128, -128, -54, 81, -128, 102, -128, -128, -28, -128, 127, -128, 127, -119, 127, 39, 8, 127, -128, -54, -117, -123, -28, -3, -78, -128, -128, -76, -128, -128, 127, 127, 127, 127, 61, 12, 58, -128, -81, -128, -128, -128, -128, -128, 32, -128, 127, 127, 127, -87, 99, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -56, -128, -128, -128, -56, 127, 27, -128, -47, -128, -128, -128, -128, 127, -61, 127, 127, 127, 127, 127, 92, -47, -63, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 51, -128, 127, -128, 15, -128, -128, -128, -128, 127, 127, -15, 127, -128, 127, 0, 127, 127, -45, -128, -128, -94, 112, 127, 41, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -87, -128, 127, -128, 127, -128, -128, 127, -128, 75, -128, -128, -128, -128, 51, -87, 121, 127, 127, 127, 127, -15, -128, 108, -73, 127, 127, 127, 127, 127, -20, -85, -128, 127, -78, 127, -128, -12, -128, -128, -128, -128, -128, -128, -128, -34, -18, 55, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 93, -128, -128, -128, -128, -128, -128, 42, -128, 71, -128, -128, 127, -128, 127, -128, 102, -128, -128, -128, -128, -128, -128, -44, -128, 127, 127, 127, 103, -128, -128, 127, -128, 127, -128, 97, -128, -128, 64, -128, -96, 127, -128, 127, 82, -128, -95, -128, 39, 127, 77, 127, 95, 32, 127, 127, 24, 127, 127, -128, -128, -128, -91, -128, -128, 127, -128, 115, -128, -56, 111, -128, -94, -128, 127, -128, 127, -128, 127, -128, -128, 25, -128, -128, -128, -128, -59, 66, 127, 127, 27, 127, 127, 34, 127, 127, 127, 127, -27, 127, -128, 127, -128, -48, -128, 127, -126, 37, -128, -128, -42, -26, 95, 127, -128, 127, -128, 127, 75, 63, -44, 52, -64, -128, 127, -128, 127, -128, -110, -128, -128, 127, 127, 127, 127, 26, 127, -126, -52, -128, -128, 127, 127, 127, 127, 76, -128, 93, -81, 127, 127, 127, 127, 127, 127, 127, 127, 127, 74, 127, -107, 127, 127, -128, 127, -72, -128, -128, 11, -128, -128, -128, -128, -128, -128, -128, 21, 5, -128, 127, -100, 127, 18, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -27, 127, -128, 127, -128, -128, -102, -128, 64, 127, 127, 127, 127, 127, 43, 127, -121, 127, 127, 127, 127, 127, 47, -96, -128, -128, -128, 127, -128, 127, -128, 74, -128, -128, -128, -128, -128, -90, 47, 127, 127, 127, 127, -128, 121, 127, 109, 127, 127, -128, 111, -128, 127, -128, 127, 127, 127, 127, 40, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -25, -128, -128, -128, -128, -128, -128, -128, -128, -128, 88, -128, 127, 127, -97, -82, -128, -78, -128, 54, 57, 127, -14, -85, 114, 127, -25, -128, -90, -40, -128, 3, 127, 127, 127, 115, 127, -93, -128, -128, -128, 4, 127, 127, 127, 127, 127, 127, 127, 61, 1, -75, -128, -32, -128, 78, 127, 127, 127, 35, 63, 44, 127, -128, 127, -128, -4, -128, -128, 127, 11, 127, -128, 127, -128, -128, -128, 15, -117, 127, 0, 127, 127, -128, 127, -11, -21, -59, -128, 5, -128, 127, -128, 61, -96, 74, -128, 59, -43, 127, 127, 104, 127, -115, 127, 127, 127, 127, 127, 127, -128, -79, -32, -128, 2, 127, -128, 127, -128, -98, 127, 68, 127, -128, 127, 90, -128, 127, -128, 41, -128, -128, -128, -128, -124, -124, 127, 26, -66, 127, -128, 127, -128, 127, -128, 127, -128, 127, 41, -49, 127, -128, 127, 127, -128, 127, 127, 127, 127, -42, 127, 78, 127, 43, -128, 127, -128, 127, 74, 127, 127, 127, 127, 66, 4, 47, 127, -125, 127, 77, 127, 127, -128, 127, -95, -93, -28, 127, 127, 127, -128, 127, 127, -128, 127, -36, 127, 127, 87, 127, 127, 127, -90, -47, -38, -30, 2, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -97, -128, -128, 127, 73, 127, 127, 127, 127, -36, 127, -128, -62, -22, -69, -59, 127, -128, 39, -128, 17, -6, 117, 127, -128, -128, -128, -128, -128, 14, 69, 100, 127, -128, 9, -128, 79, -128, 127, 127, -128, -128, -128, -61, 107, 127, -81, -35, -128, -128, 127, -49, 127, 115, 127, 127, -6, 68, 28, 127, 68, -128, -128, -91, -128, -128, -127, 127, 54, 127, -9, 127, -128, 127, -128, 127, 44, 127, 127, -128, -27, -71, -128, -128, 2, 80, 127, -116, 127, 127, 127, 127, 127, 127, 127, 127, 127, 80, -128, -128, -128, -128, 22, 127, 127, 127, 127, 127, -83, 127, -87, 127, 70, -52, 127, -128, 127, -128, 127, 127, 127, 127, -128, 94, -55, -128, -20, -69, 0, 57, -128, 127, 14, 127, -119, 127, 125, 81, 127, 127, -14, -128, 2, -128, -128, -128, -68, 127, 127, 19, 127, -128, -128, -128, -128, -128, -128, -120, -21, 127, 127, 127, 127, -128, -85, 18, -71, 127, -128, -94, -128, -128, 127, -128, 127, -128, -53, -128, -128, -60, 127, 127, 127, 127, 127, 107, -62, -128, -128, -128, -43, -128, -80, 127, 127, 127, 127, 127, 127, 127, -128, 127, -68, 127, 127, -58, 127, 127, 127, 127, 127, 127, -128, 55, 115, -113, 127, -128, -128, -128, -128, -126, 127, -43, 93, 127, -122, -128, -128, -98, -128, 127, 127, 127, 106, 127, 113, -35, -128, -128, 5, 66, -128, -18, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 4, 127, 127, 127, 127, 127, 127, 127, -97, 127, -128, -4, -113, 15, 127, -128, 88, 127, 51, 127, 127, 127, 80, -128, -128, -128, -128, -12, -106, 127, -128, 99, -128, 127, 127, 127, 19, 127, 11, 127, 127, -128, -19, -128, -128, -43, -128, 127, -15, 127, 127, -3, 76, -128, -128, -128, -128, 96, -128, 9, -128, -127, -128, -128, -128, -128, 26, 127, 127, 127, 127, -89, -44, 9, -5, -29, -128, 127, -128, 63, 77, 55, -17, 73, -128, 127, 127, 127, 127, 80, -32, 127, 127, 127, 127, 127, -128, -85, -128, 127, -53, -128, 127, -128, 70, 54, 45, 127, 127, 127, 127, 127, -128, -108, -128, -128, -128, 127, 60, 127, 127, 127, -25, 127, -18, 127, 127, 127, 127, 127, 60, 70, -128, -87, -128, -128, -128, -128, -128, -128, -72, -128, 81, 127, 127, 127, -120, 127, -128, 57, -3, -91, 113, -79, -128, -128, -128, -128, -128, 127, -99, 127, -128, -57, 127, -128, 127, -99, -68, 127, -128, 127, 124, 127, 127, -106, 127, -128, 127, 127, 127, 127, -10, -128, 32, -128, -11, -109, -82, -128, 55, -128, 127, 127, -128, 127, -128, -54, -128, -48, -128, -128, -128, -128, 60, -128, -128, 92, -128, 127, 127, -128, 116, -128, 127, 63, 127, -104, -128, -128, -128, 127, 127, 108, 1, -112, -95, 127, 127, 127, 127, 71, -128, -128, -128, 127, 127, 127, 127, -85, -128, -128, -128, -128, -128, -128, 105, 0, 127, -128, 127, -128, -128, -45, -128, 127, -128, 127, -128, 127, 127, 127, 127, 62, -128, -128, -128, -128, -75, -128, -92, -87, 127, 98, 85, 127, -128, -26, -128, -8, 127, 127, 2, 81, -128, -128, 82, -128, 105, -128, -128, 51, -29, 127, 127, 60, 127, 127, 55, 127, -128, 127, -128, 127, -68, -128, -128, -128, -128, 127, 77, 127, 127, -128, 127, -128, 89, -128, -14, 127, 127, 127, 127, 127, 127, -37, 127, 55, -128, 127, 75, 127, -75, 127, -128, -128, -19, -93, 127, 62, 127, 17, 127, -128, 11, -71, -128, -128, 127, -128, 32, 127, -49, 127, -128, -69, 88, -80, 127, 127, 127, 127, 127, 127, 0, 127, -128, 94, 109, -128, 127, -128, 86, -109, -128, 43, -128, -36, -128, -128, -128, -128, 18, -128, -128, 127, 127, 127, 127, 127, 127, -128, -22, -128, 127, -109, 119, -10, 127, -128, -128, -128, -124, -128, -62, 127, 127, 127, -74, 127, 127, 127, 127, 82, 127, 127, -109, 127, -46, 127, -128, 127, 41, 127, 127, 117, -89, -23, -128, -128, -66, 127, 127, 127, 127, 81, -119, -128, -128, -128, -91, -128, 127, 49, 127, -73, -128, 127, -128, 127, -117, 72, -6, -128, -128, -128, -128, 56, -128, 42, 127, 53, 127, 127, 5, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 74, -128, -128, 127, -128, 115, 127, 61, 127, 28, 127, 73, -128, -2, 104, -128, -106, -128, 92, -128, 127, -128, 127, -128, 14, -114, -128, -39, -128, -128, 127, -119, -69, -128, -128, -128, -128, 77, 127, 127, 127, 127, -40, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -78, -128, -21, 97, -128, -63, -128, -128, -128, -128, -128, 113, -30, 127, 100, -128, 127, -128, -47, -128, 28, 127, -128, 127, 127, 127, 127, 127, 127, 127, 32, 127, 100, -128, 28, -128, -128, 127, 100, 127, -88, 127, -128, -128, 4, -128, 127, -110, 127, -76, -128, -128, -62, -90, -128, -128, 109, -128, 127, -113, -96, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 80, 127, 127, 127, 58, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -108, 127, -128, 25, 98, -128, -57, -128, -128, -128, -128, -128, -128, -128, -128, -128, -105, -128, 26, -128, 127, 89, 127, 127, -60, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 113, 17, 127, 127, 127, 127, -128, -128, -128, -128, 0, -128, -128, -128, -128, -51, -128, -128, -128, -128, -128, -128, -86, 127, -28, 127, -88, -2, -128, -128, -128, -128, 127, -128, 127, -128, 22, 37, -128, 7, 127, -128, 127, -128, 127, -128, 127, -128, -128, 35, 69, 127, 127, 127, -9, 127, -128, -128, -128, -128, -17, -69, -21, 127, 127, 127, 127, 48, 127, 127, 127, 30, 127, -128, 127, -106, -49, -128, -128, -128, -128, -1, 58, 127, 127, 96, 127, -124, 74, -128, -128, -128, -128, -128, -128, -128, -128, 43, -87, 127, -128, -128, -99, -128, 127, 127, 127, 106, -128, -128, -128, -128, -128, -128, 127, -128, -59, 127, 74, 127, 127, 127, 59, 127, 127, 11, -38, 12, -128, -24, -128, -70, 127, -128, -99, 122, -128, 127, 127, 127, 98, -128, 127, 127, 127, 127, 70, -103, 127, 20, 127, 127, 127, 127, 103, 127, 127, 43, 127, -128, -128, -128, -128, 76, 127, 94, 127, -128, -128, -128, -128, 127, -117, 5, -128, -128, -128, -95, -26, 127, 127, 44, 127, -128, 127, -128, 127, -110, 127, 14, -128, 127, -128, -3, -128, 127, -75, 127, 127, 127, -49, 127, -128, -115, -128, -128, -128, 9, -128, -62, -128, -128, -128, 127, 127, 51, 25, -128, -128, -128, -128, 11, -41, 10, 127, -128, 127, -128, 127, 79, 127, 127, 107, -128, 51, -128, 127, 127, 127, 127, -128, 62, -128, -128, -6, -128, -128, 76, -128, 127, -128, 127, -128, 127, -128, -117, -128, -128, -128, -128, -128, -128, 18, 127, 127, 127, 127, 127, 127, -128, -74, -128, -128, -4, -62, -58, 127, -128, 127, 42, 127, 124, 24, -128, -122, -128, -128, -128, 127, 127, 94, 127, 29, 62, -12, -122, 127, 0, 123, -128, 13, -128, 127, 108, 127, 127, -128, -128, -128, 127, 43, 127, 127, -23, -124, -128, -128, 127, -128, -45, 27, -128, 127, -119, 127, 36, 100, -128, -45, 105, -128, 127, -9, 127, 127, -128, 127, -30, -123, 127, -7, 127, 127, -6, 127, 127, -128, 127, 127, -88, 127, 127, 127, 127, 127, 127, 127, -57, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 65, -106, 127, 127, 127, 24, 127, 103, 127, -128, 127, -128, -128, -128, -128, -128, -128, 75, 127, 127, -104, -66, -128, -128, -91, -128, -128, 127, -128, 127, 18, 127, 1, -128, -128, -128, -128, 127, 127, 127, 127, 22, 127, 127, -128, 127, -128, -20, -83, -128, 127, 127, 127, -18, -128, -128, -128, -128, 127, -128, 127, 13, 23, -24, 123, 25, -128, 127, -86, 127, -60, 62, -40, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -10, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 2, 127, 75, 23, 127, -128, 127, -128, -111, 85, -128, -51, 127, -128, 127, 127, 127, 127, 127, 77, 79, 6, 78, -128, -128, -128, -128, -128, 79, -128, 127, -128, 72, -128, -128, -128, -128, -128, -128, 119, -128, 127, 127, 127, 127, -128, 59, -128, -128, -128, -128, 28, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 43, 19, 127, 106, 127, 127, -6, 100, -55, -17, -128, -128, -128, -5, -128, -66, -128, -128, -123, -128, 127, -128, 32, 127, -128, 127, -5, 127, 77, -80, 127, 92, 127, 127, 48, 127, -128, 127, -128, -128, 127, -128, 127, -128, -76, -128, -128, 127, 127, 127, -77, -8, -128, 127, 7, 127, 127, -128, 127, 87, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -56, 113, -128, 127, -128, 127, -128, 55, 1, 17, 127, 85, 127, -24, 104, 127, -128, 23, -128, -128, 127, -104, 127, -82, -34, -128, 127, -128, 127, 127, 127, 127, 127, -13, 0, -128, -128, -128, -128, 115, -128, 127, 127, 127, 127, -128, -40, -29, -29, 127, -55, 120, -128, -128, -128, -128, -128, 127, 127, 127, 77, 127, -128, -128, -128, -128, 127, -53, 127, 127, 127, -128, -128, -128, -128, -108, -128, 45, 51, -22, 127, -128, 75, -90, -9, -128, 9, -128, 127, -28, -128, 127, -128, -24, -128, -128, 24, -128, 127, -96, -125, 127, -128, 127, -128, -76, -128, 23, 127, 127, -128, -48, -128, -128, -22, 17, 85, -128, -80, -78, 34, 127, 127, 127, -85, -60, -128, 18, -128, 127, 53, 127, -128, 113, -128, 49, 127, 42, 127, 127, 127, 43, -21, -128, -128, -128, -128, -64, 127, -128, 127, -128, -128, 97, -73, 127, -116, 127, -45, -94, 85, 127, 93, -128, 0, -69, -128, -128, -2, -128, 127, -63, 127, 93, 127, -128, -91, -128, -128, -128, -106, -91, 127, -66, 127, 34, 95, 127, -57, -128, 127, -128, 1, 21, 127, 127, 127, 54, 127, 117, 127, 127, -56, 127, 25, 127, -128, 15, -128, -128, 127, 127, 127, 127, 127, -65, -128, -128, -128, -128, 127, 0, 115, 127, -44, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -40, 1, -128, 127, -128, -128, -128, -128, -128, -43, -68, -66, -109, -56, -128, 127, 127, 127, 59, 127, 127, -32, 7, 127, 80, 121, -128, -128, -51, 76, -99, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -96, 127, 35, 127, -128, -128, -128, -128, -23, 127, 127, 127, 127, 127, 127, 127, 70, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -93, -128, 127, -128, 127, -128, -74, -128, -128, -128, -85, 127, -60, 127, 28, 127, 127, 127, 127, 127, 127, 127, -128, -10, -128, -128, -128, -128, -128, -128, 23, 127, -23, 127, 127, 53, 127, -128, 127, -128, 127, 125, 127, 127, -128, -62, -128, 25, -128, -128, -128, -128, 15, 32, 127, -128, -14, -128, 77, -89, 127, 127, 127, 127, 39, 55, -128, -43, -6, 127, 127, 127, 127, -128, 13, -49, -128, 127, -53, 127, 127, 54, 127, -128, -128, -128, -98, -128, 127, 127, 127, 127, -43, 127, -128, 127, 45, 127, 127, 127, 127, 25, -128, -128, -37, -128, 127, 127, 127, 127, -128, 15, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 112, 53, 127, -100, -91, 58, -128, 127, -128, -128, -128, -128, 127, 13, 127, -29, 127, -5, 120, -5, 127, -128, 127, -128, -128, -89, -128, 107, -128, 76, 127, 115, 127, -56, -128, 30, -108, 54, -48, -128, -128, 47, -128, 127, -128, -22, -128, -128, -128, -26, -128, 89, -77, 127, -95, 127, 57, 127, 78, -128, -17, -128, -128, -128, -128, -128, -55, -59, -128, -128, -108, -128, -128, -128, -128, -92, -128, 127, 127, 127, 127, -91, -128, -128, -128, 23, 127, 127, 127, -128, -68, -58, -128, 127, -128, -17, -35, -128, 25, -128, 127, 127, 5, 127, 125, -24, 127, 37, -10, -105, -74, 127, 9, 127, 127, 70, 127, -128, -115, -128, -128, -128, -128, 127, -78, 127, 1, 127, -17, 102, -128, -128, -128, -128, 127, 127, 127, 127, 127, 30, -97, -73, -123, 127, -128, 19, -128, -92, -128, 127, 44, 127, 23, 127, 127, 127, 127, -117, -26, -128, -128, 113, -128, 127, 127, 2, 127, -128, 127, -106, 127, 127, 127, 3, 127, 52, 127, 70, 127, -66, -128, -128, -128, -128, -128, -128, -128, -39, -95, 127, 127, 127, -128, -128, -7, -128, -18, -128, 127, -128, -8, 127, -128, 127, 64, -54, 127, 65, 127, 81, -128, -128, -128, -128, 109, 127, 127, 127, -103, -128, -128, -128, -128, 127, -128, 104, -128, -128, -128, 111, 127, 127, 127, 127, 127, -28, 74, -128, -45, -128, -11, 29, 127, -128, 36, -128, -128, -128, -128, -128, -128, -128, 43, 68, 127, 127, 21, 127, -128, 127, -128, -79, -128, -128, -106, -128, 127, -70, 20, -128, -62, -128, -128, -128, 68, 127, 127, 127, 127, 127, 34, -128, -17, -128, -128, 0, 60, 127, 127, 127, 127, 127, -128, 127, 63, -128, 127, -128, 127, -66, -46, 127, 18, 127, 127, -128, 109, -128, -128, -98, -128, 92, -128, -128, 102, -128, -91, -128, 127, 127, 127, 127, 127, -41, -128, 91, -128, 127, -7, 127, 127, 6, 127, 127, -94, 127, -9, 127, -56, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 125, 127, 127, -128, -46, -74, -128, 94, -128, 76, -128, 73, 127, -116, 127, -13, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 4, -51, -128, -128, -128, -128, -128, -128, -128, 108, -24, 127, -128, -128, 127, -128, 127, 127, 127, -82, -128, -128, -128, -128, -128, -66, -128, -128, 72, -81, 127, 127, 127, 127, -128, -98, -128, -128, 127, -128, 127, 127, 34, 127, 127, 127, 127, 127, 127, 127, 127, 2, 19, -128, -128, 48, -128, -1, -128, 127, -128, 127, 39, 102, 127, 78, 104, 127, -128, 127, -128, 121, -83, -34, -30, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 97, -128, -128, -128, -128, 0, 3, -128, 127, 20, -128, 127, 127, -128, 127, -32, 127, 30, 127, 127, 127, 127, 127, 127, 127, 127, 75, 127, -96, 127, -128, 127, 127, -128, 127, -35, -72, -64, -128, 30, -128, -26, -128, -128, -128, -128, 26, 58, 25, 127, -128, 127, -128, -128, -128, -128, 110, 127, 127, 127, 127, 127, 88, 127, 127, 127, 127, 127, -124, 73, -128, -128, 127, -128, 127, -75, -128, -128, -128, -128, -128, 127, 127, 127, -20, -128, -128, -128, -128, -106, 45, -74, 127, 32, 127, 98, 23, 127, -95, 127, 85, 127, -128, 127, -128, -119, -18, -18, 127, 127, 127, 123, 127, -128, 127, -128, -128, -128, -128, -81, 109, 127, 127, 127, 127, 127, 127, -23, 10, 94, 87, 127, 127, -38, 127, 127, -52, 127, -66, 127, -128, -128, -128, -128, -128, 127, -128, -116, -54, -128, -128, -1, 63, 127, 38, -128, -52, -128, 127, 121, 127, 127, -128, 71, -128, 127, 93, 3, -128, -128, -128, -75, 29, 127, 127, 127, 127, 127, 127, -63, -128, -102, -128, 109, 37, 127, 107, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 97, 127, 127, 127, 107, 127, -128, -51, -128, -128, -128, -128, 64, -128, 127, 127, 127, 63, 87, -31, 127, -128, 96, -128, -69, 59, -128, -30, -128, -8, -124, 127, 127, 127, 114, 95, -128, 114, 127, -79, 127, -8, 127, -128, 9, -128, -128, -72, -128, 127, -58, 127, 127, 18, 127, -128, -128, -128, -128, -128, -128, 12, -128, 127, -128, 127, -45, 103, -13, -128, 127, -128, 127, 59, 127, -128, -85, 127, 127, 127, 127, 127, 127, 127, 127, -10, -128, -128, -128, -128, 127, 127, 127, 106, -128, 112, -128, 127, -78, -128, -128, -128, -128, 127, -85, -128, 127, -128, 127, 127, 127, 127, 127, -64, -49, -128, -96, -128, -128, 127, -128, -128, -128, -128, 83, 127, 127, 14, -52, -47, -128, 127, -128, 96, -128, -128, -128, -128, 127, 3, 127, -75, 127, 88, 127, 127, 127, 127, 44, 126, 127, 127, 127, 109, 52, 127, -44, 127, -128, 8, -128, -128, -128, 68, 96, 79, 127, 60, 127, -89, -128, 24, -128, 127, -128, -39, -62, -128, 127, 127, 127, 94, 127, -128, -83, -128, -128, -52, -23, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 48, -128, -128, 19, -128, 127, 127, 127, 127, 127, 127, 28, -128, -87, -128, 127, -128, 127, 42, 127, -60, 127, -128, 127, -128, -55, -128, -128, -111, -27, -128, 127, -98, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 11, 127, 46, -124, 127, -121, 127, 66, 21, -128, 22, -41, -73, -128, 127, -128, -5, -128, 127, -68, 127, 86, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -40, -128, -128, 127, -128, 127, -128, -51, -56, -128, -128, -75, 10, -127, 109, -116, 8, -128, -128, 8, -75, 127, -128, 125, -128, 127, 127, 127, 127, -128, -75, -128, 127, -128, -128, -64, -128, 37, -128, -70, 127, -63, 127, 127, 127, 127, 127, 127, -128, 14, -128, 91, -128, 127, 87, -128, -128, 44, -128, 127, -21, -9, -55, -128, 127, 127, 38, 127, 36, 40, 88, 127, 127, 62, 127, 127, -128, 18, -128, 70, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 4, -128, -127, -128, -128, -128, -128, -85, -128, -128, -128, -128, -128, 108, -76, 127, -128, -128, -54, -128, -128, -51, -128, 127, -117, 115, 127, -30, 127, -21, 127, -123, 127, 127, 54, 127, -128, 62, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -121, 127, 127, 127, 127, -128, -128, -119, -22, 79, 127, -128, 32, -35, -128, -125, -79, 26, -9, 127, 35, 127, -73, -106, 127, -21, 127, -128, 127, -128, 127, -114, 98, -128, -128, -128, 97, -128, -128, -128, -128, -42, 127, 120, 127, 100, -128, 48, -128, 127, -48, 17, 127, 127, 127, 22, 127, -128, -128, -128, -128, -128, 57, -124, 127, 127, 127, 127, 19, -128, -128, -17, -128, 127, -128, -128, -28, -128, -103, 79, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 12, 127, 127, 127, 127, 127, 127, 127, 125, -128, 127, -119, 77, 127, 127, 127, 127, 127, 127, 127, 127, 47, -128, 24, -128, -3, -25, 127, 17, 127, -128, -128, -73, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -58, 127, 127, 45, 96, -128, -128, 82, -128, 127, -128, -128, -128, -128, -128, -49, -128, -128, 127, 57, 127, 127, 39, -128, -128, -78, 8, 127, 24, -128, -128, -90, 109, 127, 127, 127, 127, 120, -2, 127, 75, 127, -128, -44, -128, -8, -128, 127, -19, 127, -13, -97, 127, -128, 127, -128, 97, 127, -128, 127, -128, 127, 112, -128, -128, -128, -128, 14, -128, 24, 29, -128, 47, -128, 127, -8, 127, 127, -128, 127, -128, -128, -128, -128, 127, 81, 127, 127, -128, 46, -128, 127, 127, -9, 127, -128, -128, 102, -113, -36, -128, -128, 127, -128, -75, -89, -128, -128, 127, 28, 127, 127, 127, 127, 127, 127, 127, 127, 76, 127, 90, 127, 5, 127, 127, 127, 37, -128, -128, -128, -128, -128, 127, -128, 127, 123, -5, 127, -106, 127, 36, 127, -128, 111, -71, 127, -12, 127, 127, 127, 102, 38, 127, -128, 108, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -28, 127, -115, -128, -128, -128, -128, -128, -128, -44, 18, 127, 127, 127, 127, -8, -73, -128, -128, -88, -31, 79, 127, 127, -81, -98, -128, -128, -128, -128, -128, -79, 71, -93, 127, -128, 127, -42, -128, -128, -128, 100, -128, 127, 127, 127, 127, -128, 35, 48, 2, 127, 127, 81, 127, 127, -128, 75, -128, -128, -128, -3, -128, -128, 127, 75, 127, 127, 127, 127, 127, -128, 127, -128, -128, -99, -128, 127, 127, 127, 127, -2, 127, 127, 36, 127, -128, 127, -128, 127, -128, 5, 114, 127, 127, 127, 127, -15, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 34, -128, -112, -128, 127, 77, -97, -83, -128, -128, -128, 127, -66, -128, -112, -128, 108, 55, -119, 22, 127, -14, 127, 127, -24, 127, 0, 127, 127, 127, 127, 71, 127, -128, 127, -73, -114, 74, -128, 127, -128, 95, -99, -128, 4, 1, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -125, 49, 127, -128, -55, -128, 83, -64, -46, 127, 120, 127, -128, -81, -57, -128, 127, -128, 127, -79, -128, 127, -128, 127, 6, 127, 13, 4, -17, -128, -125, -128, -128, 127, 42, -128, 90, -128, -13, -128, 46, -128, 127, -128, 19, -128, -128, -29, -128, 12, -74, 74, 127, -83, 127, -31, 26, -128, -128, 127, -128, 127, 127, -128, 95, -128, -128, 34, -128, -125, 78, -128, 68, 127, 127, 127, -128, 24, -128, -128, -128, 5, 96, 100, -11, 91, -128, 127, -128, 127, -44, 127, 127, 61, 127, 127, 124, -128, -128, -128, -128, -112, -128, -128, -94, -128, 119, -128, 14, 127, 127, -9, 127, 12, 95, -128, 29, -128, -90, -11, 98, 127, 127, 127, -105, -128, -128, -107, -128, -75, 91, 127, 127, 116, 127, 113, -87, -128, 127, -128, 127, -83, 127, -128, 127, -128, -128, -128, -128, -128, -28, 75, 127, 127, 127, 127, 127, 127, 25, -128, -3, -60, 127, 127, 127, 95, -128, -20, -128, -128, -128, -128, -128, -128, -128, 59, -108, 89, 104, 38, 127, 104, 127, 127, 127, 25, 39, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 1, 127, 127, 127, -6, 127, -99, 27, 0, 69, 127, 127, 127, 78, 127, 127, -128, -128, -128, -128, 7, 127, 65, 127, -128, -43, -128, 64, -128, -111, 127, 41, 127, 127, 127, -12, -121, 92, -128, 127, -90, 15, 127, -128, -128, -128, -128, -128, -83, 127, 127, 127, 127, 97, -128, 127, -128, 127, 93, 83, 127, -128, 127, -24, 127, 127, -128, -128, -26, -109, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -113, -128, -128, -128, -128, 117, 127, 127, 127, 127, 127, 127, 127, 127, 127, -124, -128, -121, -32, 127, 127, 127, 127, 127, 54, -128, -58, -60, 127, 127, 127, 127, 127, 127, -87, 127, -128, 18, -128, 9, -68, 127, 127, 60, 127, -15, 112, -128, 127, -128, -32, -49, 21, 127, 127, 109, 127, 32, 127, -128, 127, -128, -32, 26, -65, -128, -128, -128, -128, 127, -128, 127, -97, -72, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 32, 127, 127, -97, 127, 26, 127, 127, 127, 2, -128, -128, -35, -23, 73, 127, 22, 127, 115, -17, 90, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -45, 66, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -98, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 13, 127, -128, 127, -95, 86, -128, 127, 127, -125, 68, 104, -70, -128, 72, -105, 21, -128, -128, 127, 74, 59, 127, -128, -18, -128, -128, -128, -128, 13, -117, -7, -59, 127, 75, -23, -112, 127, -128, 7, -128, -128, -128, -128, -122, -128, -102, 95, 14, 127, 127, 127, 127, -128, -109, -128, -128, -128, -128, 89, -128, 127, -68, 127, 127, -93, 127, 62, 127, -128, -51, -128, -128, -128, -128, -18, 127, 85, 127, 127, 127, 127, -1, 95, -128, 127, -128, 127, -128, -97, -128, -128, -128, -48, 100, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 0, 127, 127, 127, -128, 3, -128, -115, -128, 116, 12, 121, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -7, -125, 63, 127, 127, 127, 127, 127, 127, 127, 43, 127, -15, 52, 36, -114, -128, -128, -128, -128, -128, -128, 0, -30, 127, 35, -128, 25, -128, -128, -128, -128, 79, 12, 63, 76, -128, -128, -77, -128, 127, 127, 127, 127, 127, 127, -128, -41, -128, 12, -128, -128, -70, -128, -45, 127, 127, -128, 127, -128, 56, -83, -128, 127, 127, 34, 127, -128, -128, -128, -128, 0, -113, -10, -104, -128, -91, -62, 124, -128, 127, 127, 127, 127, 127, 127, -72, 127, -128, 127, -128, 57, 109, -34, 127, -128, 24, -128, -128, 127, 88, -22, 127, 127, -66, 60, -128, -64, -128, 91, -56, 127, -128, 127, 127, 7, 127, -72, 127, 127, -89, 127, -128, 60, -128, -128, -128, -128, 29, 127, -128, 127, -128, -95, 11, -82, 127, 127, 127, 127, 11, -128, -128, -128, -128, 127, -128, 66, -45, 45, -42, 63, -128, -128, -128, -128, -6, -128, 85, -128, -128, -128, -128, 49, -19, 114, -43, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -103, -22, 98, -128, -128, 15, -128, 127, 127, 127, 127, 127, -121, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -31, 72, -80, -128, -128, -46, 127, 127, 127, 34, -128, -128, -128, -128, -128, -128, 68, -128, -128, -128, -128, -128, -41, 77, 127, 49, 127, -37, -68, -104, 85, -128, 77, 127, 36, 127, 127, 41, 127, 127, 127, 127, 107, 10, 41, 127, -3, 127, -54, -128, -128, -128, -128, 127, 127, 127, 22, 127, 115, -104, -128, 21, -128, 12, -128, -99, -128, -128, -44, -128, -54, 127, 0, -128, -128, -128, -128, -26, -128, -6, 127, 40, 2, 127, 127, -6, 127, 127, 11, 127, 1, 127, 127, -128, 127, -128, -58, -128, -128, -128, -128, -85, 56, 127, 127, -128, -73, -128, -87, 127, 127, 127, 127, -128, 127, -128, 28, -128, -23, 108, 127, 115, 127, -128, 104, -78, -92, -63, -128, 29, -128, -51, -128, -128, -128, -77, -128, -65, -5, 53, -25, -128, -72, -128, 127, -120, 127, 127, 127, 44, -46, -128, -128, -128, -128, -128, -27, -128, 59, -128, 127, -107, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 112, -106, -128, -22, -128, -128, -128, -128, -128, 53, 127, 127, 6, 53, -128, -128, -61, -128, -128, -128, -128, -49, -128, -19, 127, -14, -128, -128, -128, 104, -128, -117, 10, -128, -82, 97, 78, 107, 127, 12, 127, -34, 127, -34, 109, 127, -128, 107, 119, -128, 127, -20, 127, -128, -128, -128, -43, 127, 127, 127, 127, -117, 127, 26, 127, 127, 127, 127, -69, 127, -128, -92, -128, 58, 39, 127, -75, 127, 61, 78, 55, -99, -128, -37, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -52, 127, -128, 127, -128, 81, 23, 23, -21, -128, -128, 127, -128, 127, 17, 127, -122, 40, -128, -107, -25, -128, -128, 78, -31, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -37, -128, -108, -128, -128, -22, -128, 127, -25, 127, 127, 127, -128, 75, -128, 127, -128, -128, -38, -126, -128, 66, 127, -128, 127, -128, -128, 2, -128, 127, 127, 127, 127, 32, 127, 70, 14, 127, 91, 127, 39, 127, 127, 127, 25, 91, -128, -52, -128, -128, -128, 127, -128, -128, 127, -26, 58, -117, -128, 2, -128, -128, 127, 92, 127, -97, 41, 88, -128, 127, -128, 127, -128, 127, -128, -90, 1, -128, 56, -128, -100, 120, 127, 127, 14, 127, 127, 127, -79, -128, -128, -128, -128, -128, -128, -2, -128, -128, 7, -128, -128, -128, -60, 47, 102, 127, 127, 127, 127, 127, 127, 77, 127, 38, -128, -128, -128, -128, -128, -128, -100, -128, 73, -128, 96, -128, 127, -128, -13, 127, -128, 97, -128, -3, -128, -7, 35, 127, 127, 127, 127, 102, -128, 127, -128, 127, -29, 127, -32, -128, -77, -128, -128, 127, 20, 127, 127, 124, -22, -128, -107, -128, -17, 73, 127, 127, 127, 38, 122, -76, -117, -128, -128, -128, -128, -122, -128, -128, 127, -128, 26, -128, -61, -128, -114, 52, 127, -128, 127, -128, 127, -128, 127, -99, 127, 127, 9, -96, -128, -128, -128, -128, -128, -128, 66, -53, 127, -128, -128, -92, -128, 127, 45, 127, 127, -128, -128, -128, -128, -128, 83, 75, 127, 127, 127, 64, 127, -128, 127, 127, 127, 127, 127, 127, -31, 127, -128, -39, 127, 127, 127, 71, -89, -128, -128, -128, 51, -128, 127, 45, 127, 82, -128, -128, -128, -128, -128, 127, -69, -32, 121, -128, 127, -128, 127, -20, 127, 127, -110, 127, -128, -27, -35, 106, 127, 51, -128, 68, 100, -128, 38, -128, -12, -128, 127, 127, 127, 127, -128, -128, -128, -77, -128, 20, -13, -128, 89, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -79, -128, 127, -78, 127, -9, 127, -55, -128, 127, -128, 127, 127, 127, -24, 68, -61, -52, -55, 127, -128, 127, -128, 127, -121, 127, 127, 127, -128, -39, 45, -128, 127, -100, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -93, -128, 127, 127, -108, 127, -128, 121, -128, -128, 17, -38, -128, -128, -83, -128, 28, -128, -128, -51, -128, 127, 127, 127, 127, 114, -128, -128, -128, -128, 121, 127, 127, 127, 127, 127, 127, 127, 127, -72, 90, -128, -108, -128, -56, 124, 12, 97, 0, -128, -128, -128, 127, -57, 127, 127, 127, 127, 127, 61, 127, 127, 114, -3, 127, -128, 127, 23, -128, 127, -117, 5, -108, 127, 30, -128, -128, -70, -128, -128, -128, -13, -128, -128, -128, -25, -128, -46, -128, 126, -128, -7, -119, -128, 127, 10, 127, -17, 127, -128, -128, -128, -128, -15, -128, -44, -48, 127, -127, 127, -128, -99, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 119, 127, -24, 127, -128, -128, -128, -128, -128, -128, 95, -128, 22, -128, -128, 98, -128, 127, 127, 74, -71, -128, -128, -128, -128, 34, -128, -61, 97, 21, 127, 127, 11, 111, -92, -128, 127, -128, 127, -128, -128, 10, -128, -51, -42, 127, -128, -40, -128, -128, -128, -128, 127, 127, -99, 127, -128, 59, -46, -128, 127, -21, -57, -128, -87, -128, -128, -128, -128, -128, -46, -128, -55, -128, -57, -128, 127, 127, 127, 95, 127, 2, -128, 125, -88, 10, 14, 46, -30, -128, 127, 127, -126, 127, -63, -40, 127, 127, 127, 127, -28, -57, -128, -128, -128, -85, -128, -128, -121, 127, -23, -42, 127, -128, -128, -128, -128, -128, -112, 9, -128, 127, -128, 127, -128, -128, -31, -128, -119, -128, -124, -4, -97, 127, -128, 60, -128, -74, -128, 127, 127, 127, 127, 127, 127, 122, 127, -60, -128, -128, -128, -128, 25, -128, 77, -128, -128, 127, -128, -128, -128, -128, -91, -128, 127, 8, 127, -128, -66, -128, -128, -128, 127, 27, 127, 127, 127, 127, 127, 127, 127, -11, -7, -128, -128, -128, 127, 127, 127, 127, -110, 119, -128, -39, 1, -128, 127, 127, 127, 127, 18, 127, -128, -48, -128, 127, 127, 127, 127, 38, 73, -128, -128, 43, -83, 70, -116, -31, 127, 127, 127, 127, 127, 127, 55, 127, 127, -128, 127, -128, 127, 127, -57, 127, -123, 127, 59, -128, -47, 8, -128, 26, -128, -128, 127, -128, 127, 127, -106, 127, -128, 87, 127, -128, 127, -128, 87, -128, -128, -128, 97, 127, 127, -128, -128, -128, -128, -128, -128, -128, 13, -128, 127, 127, 127, 127, 127, 127, 127, 52, -24, -128, -128, 78, 23, 36, 127, -77, 127, 63, 127, 127, -128, -9, -128, -128, -128, -128, -128, -128, -128, -128, -128, 34, -128, 127, -128, 127, -128, -90, -120, -128, -128, -53, -128, 22, 23, -128, 105, -128, 127, 127, 127, 127, -128, -70, -128, -43, -128, -128, -128, -128, -128, -128, -15, -43, -128, -128, -128, -19, -128, -14, 18, -128, 127, -128, 127, -128, 70, 65, -128, 14, 127, -61, 127, -128, -128, -128, -128, -128, -128, 100, 127, 127, 127, -128, 127, -128, 127, -89, 57, 75, 40, -68, 127, -27, -61, 90, -32, 39, -128, -128, -128, -128, -128, -128, -5, -99, -91, 127, -99, -128, -35, -128, 127, -128, -128, -88, -128, -128, -7, 127, 127, 127, -49, 93, -128, 127, 81, 127, 127, 18, -128, -86, -73, -43, 127, 127, 127, 32, -128, 127, -128, 127, 127, 26, 127, -128, 127, 76, 127, 127, 127, -59, -128, 127, -4, 127, -128, -102, -128, -128, 127, 127, 127, 127, 127, 111, 127, -128, 127, -78, 127, -128, -43, -128, -128, -128, 127, -128, 127, -128, -6, -128, -128, -8, -28, -128, 18, -128, 127, 127, 127, -6, 127, 32, 127, 127, 127, 127, 127, 127, 127, 127, 1, -128, 52, -128, 122, -128, -128, -128, -128, 41, -128, 127, 127, -29, 22, -128, -128, -128, -73, 127, 127, 127, 127, 127, -36, -74, -81, -128, -99, -128, -68, -128, -128, -128, -128, -128, -128, -109, -128, -128, -128, -99, -112, 127, 127, 127, 81, -128, -128, -128, -128, -128, -128, -74, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 70, 127, 127, 82, 120, -128, -128, -128, -128, -28, 80, 122, 127, 127, 127, -122, -128, -128, -128, -128, -128, 127, 127, -37, 127, -128, 127, -128, 127, -12, 127, 127, -7, 127, 80, -106, 25, -128, -128, -104, -128, 127, -74, 127, 127, 127, -128, 127, -87, 127, 127, -94, 127, 127, -128, 127, -128, -128, -128, -128, -27, -95, -42, 127, -5, 127, -128, 127, 127, -128, 127, -128, 127, 127, 5, 127, 127, 127, 127, 127, 127, 127, 96, 106, -128, -128, -128, -128, -128, 20, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -72, 127, -128, -24, -128, -102, 127, -128, 127, -128, -94, -128, 43, -74, -128, -124, -128, -128, 115, 14, 127, 127, 127, 127, 127, 127, 96, -128, -39, -128, -119, 88, -128, 127, -128, 127, -128, 127, 127, 127, 127, 123, -3, -128, 74, -128, 74, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -80, 127, 127, 127, 127, -128, 22, -128, 127, 127, 127, 83, 127, 112, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -47, -128, 96, -128, 72, -128, 30, 46, 127, 90, 27, 127, -128, 127, -14, 76, 0, 127, -128, -128, -128, -128, -128, -128, 127, 127, 20, 127, -128, -128, -128, -128, -128, 43, 7, -57, 3, 127, -128, 127, -128, 108, -64, -128, 127, -128, 13, 36, -26, -36, 127, 127, 30, 127, 127, 127, 127, 127, 57, 127, -114, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 27, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 66, -128, 122, 127, 34, -128, 37, -128, 55, -128, -128, 127, -128, 127, -73, 127, -81, -128, -128, -128, -128, -128, 127, -128, 51, -128, -128, -128, -128, -95, -128, 127, -38, 127, 9, 127, -83, -128, -61, -128, -74, -127, -5, 127, -128, -17, -128, -128, -128, -128, -128, -128, -120, -128, 127, -57, 127, -128, -112, -128, -64, -128, 24, -128, -79, 127, -128, -128, 127, -128, -13, -128, -11, 127, 127, 127, 127, -128, -128, -7, -128, 127, 30, 127, 127, 34, 127, -128, 51, 127, 0, 127, 127, 127, 48, -128, 127, -128, 127, -128, 61, 127, 90, 127, 127, 25, 40, -128, 66, 127, -128, 127, -39, -128, 127, -111, 46, 127, 127, 127, 127, 59, -41, 127, -128, -128, -103, -128, 127, -45, 127, 127, -128, 127, 20, 71, 4, -128, 72, -128, -128, 73, -128, 127, 23, 127, 127, -38, -74, 52, -128, 127, -128, 99, 30, -117, -93, -128, -128, -126, -128, 127, 127, 127, 127, -20, 127, 95, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -120, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -61, 127, -128, -128, 127, -96, 127, -99, 29, -128, -128, -128, 73, 127, 92, 127, 3, 0, 127, 127, 127, 127, 127, -68, 7, -128, -128, 127, -128, 127, -128, 127, -128, 90, 127, 45, 127, -128, 121, 87, 127, 127, 127, 56, -128, 127, -128, 127, -128, 21, -128, -128, 59, 127, -56, 127, 112, -128, 127, -128, 127, -105, 121, 127, 127, 114, 127, 127, 127, 127, 127, 127, 127, 127, 126, -128, -128, -128, -128, 36, -128, 127, 127, 127, 127, -128, 127, -71, 1, 127, -38, 127, 40, 2, 83, -128, -51, -112, -128, 127, 127, 127, 127, 127, 127, 127, 89, -30, 53, 127, 127, 127, 127, -128, -11, 2, 111, 127, 127, 127, -52, 32, 48, 127, -91, 127, -128, 11, -128, -128, 127, -128, 127, -89, 127, -128, 127, -71, -128, -128, -128, -128, -128, -93, -128, 127, 40, 127, 63, 127, 127, -104, 127, -128, -128, -128, -128, 12, -23, -52, -11, -97, -55, 73, 127, -49, 127, 39, 127, -128, -107, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -24, -44, 57, 127, 47, 127, 124, -58, -34, -77, -128, -60, -128, -128, 117, 127, 127, -17, 127, -58, 127, -128, 127, -128, -51, -128, 127, 127, 127, 127, 127, 30, -128, 21, -128, -66, -128, 127, -128, -4, -60, 127, 127, 127, 127, 31, 127, -76, 127, 127, -128, 127, -128, -128, -128, -128, 74, 127, 127, 125, 127, -128, 127, -21, -39, -9, 127, -128, 17, -128, 127, 127, 127, 127, 127, -128, -17, -128, 127, -128, 112, 127, 8, 127, 127, 127, -73, 127, 127, 127, -11, 88, 4, -128, 14, -128, -17, 124, 127, 127, 127, 127, 127, 127, 112, 23, 127, -128, 127, 127, 127, 127, -128, 127, 89, -128, 125, 40, 127, 127, -128, 127, 127, 109, 127, 36, -12, -103, -128, -128, -128, -128, -81, 127, 121, 127, 127, 55, 127, 39, 36, -31, -128, -46, -128, -128, 127, -128, 126, -128, -128, -128, -128, -128, 127, -116, 127, 127, 54, -39, -128, -128, -58, -128, 108, 127, -93, -128, -128, -128, 127, 127, 127, 127, 127, -85, 127, -128, 127, 26, -128, 109, -128, -49, 75, -128, 127, -128, -128, 127, -128, 127, -87, -28, -128, -128, -116, -128, -128, -128, -128, -128, -58, -128, 127, -128, 75, -34, -128, 12, -128, -128, 19, 108, 127, 127, 127, 127, 127, 25, -15, -128, -128, -128, -128, 127, -128, 127, -123, 125, 127, -25, 127, 127, 127, -128, 127, -128, -128, -29, -128, 127, -128, -127, 27, -128, -128, 36, 21, 11, 127, -89, 111, -85, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -110, 127, 127, 127, 127, 127, -128, -51, -128, -128, -128, 57, 98, 127, -128, -128, -128, -128, -128, 127, -35, 27, -128, -85, 49, 127, 127, 127, 127, -13, 127, -128, 127, -128, -128, -65, -128, 64, 114, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -46, 127, 127, 96, 117, -56, -59, -128, -99, -128, -107, -128, 78, 127, 127, -58, -128, 127, 23, -128, 127, -42, 127, -128, 65, 127, 24, 127, 127, 106, 127, -104, 58, 38, 35, 127, 127, 86, 127, 23, -128, -128, -124, 105, 79, 127, -91, 0, -128, -128, 36, -128, 35, -128, 95, 127, 127, 127, 127, 127, 4, 58, -128, -128, -128, -128, -128, 82, -128, -128, -38, -128, 127, -128, 127, -124, 69, 127, 127, 127, 127, 127, -25, 127, 127, 127, -102, 127, -128, -94, -128, -76, 127, 51, 127, 127, 127, 127, 127, 44, 127, -70, 127, 87, 127, 103, -128, 26, -128, 95, 52, -128, 115, -128, -15, -128, -128, 127, 127, 127, 127, 127, 127, 94, 77, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -102, -128, 127, -128, 127, 108, -5, 78, -25, -128, 8, 10, -128, -64, -85, -128, 127, -109, 127, -115, 39, -128, -82, -41, 127, 89, 127, -128, 127, -128, 127, -128, 127, -128, 45, -128, -128, -128, -128, -128, 58, -74, 127, -128, -37, -128, -128, -128, 14, -128, 127, -128, 127, 127, 127, 127, 127, 43, 55, -12, 122, -128, -71, 127, -128, 127, -128, 25, -128, -128, -128, -128, -120, -128, 127, -128, 127, -128, 127, -19, 127, -55, -128, -128, -128, 127, -80, 127, 127, 62, 115, 127, 30, 127, 127, -128, 127, -128, -111, -128, -128, 127, -65, -55, 127, -128, -105, 93, -78, 127, -19, 127, -104, -128, -128, -128, -128, 127, -4, 127, 36, 127, 127, -68, 52, 127, 52, 127, 127, 111, 127, 62, -128, 127, 127, 127, -114, 87, -128, 127, 127, 127, 127, -54, 127, 127, 127, 127, 127, 127, 0, -128, -128, -128, -98, -128, -53, 82, -128, 25, -89, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 77, -128, 127, -128, 127, 127, 34, 127, -128, -128, -128, 68, -128, 107, -128, -128, -128, -128, -128, -88, 127, 127, 127, 78, 4, 36, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -73, -94, -128, -78, -128, 127, 127, 45, 127, -74, -79, -128, -128, -128, -8, 60, 127, 102, 127, 127, -32, -29, 127, -128, -128, -128, -128, -25, -128, 127, 127, 108, 127, -128, 127, -128, 127, -38, -68, -128, -128, -128, -128, 111, 49, 127, -87, 48, -128, -128, -128, 63, -128, 127, 127, 127, 127, 127, 72, 127, -12, -128, -128, -128, -128, 0, 58, 127, 127, 127, 127, -128, -42, -128, 9, -128, -128, 127, 102, 127, 127, 112, 127, 117, 127, -128, 19, -128, -128, -128, -128, -112, -71, -62, 127, 127, 127, 127, -128, 107, -128, -128, 127, 55, 127, -21, 127, -38, 127, 127, 127, 127, 110, 127, 127, 127, 106, 127, -128, -128, -128, -128, 127, 59, 127, 114, -128, 127, -128, 127, -128, -128, -44, -128, -76, 127, -73, 127, 127, 61, 127, -128, 127, -128, -128, 83, -128, 127, -19, 64, 127, -70, 127, -128, -128, -126, -128, 127, 127, 127, 127, -120, -81, -63, -128, 127, -128, 127, 127, 127, 127, 127, 63, -9, -128, -128, -128, 24, -121, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -77, 127, 93, 127, 127, 127, 127, -128, -128, -128, 60, -128, -71, -128, -128, -128, -128, -128, -109, -29, -128, -128, -5, -128, -128, -91, -47, -51, -128, -128, -128, -128, -128, -128, 109, 127, 125, 127, 127, -125, 127, -23, 91, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -18, 123, 127, 127, 127, 127, 103, 127, 60, -128, -128, -128, -128, -128, -128, -128, 127, -31, 127, 127, 127, -128, -128, -117, -128, -87, -128, -21, -128, -128, -14, 127, 127, 127, 26, 87, -121, -128, -128, 85, -128, 127, 41, 3, -12, -128, 127, -128, -80, -128, -128, -128, -49, -128, 127, 127, 49, 127, -128, -128, -128, -62, -128, 122, -128, -128, -128, -128, 70, -71, 3, 113, 127, -72, -103, 4, -128, 127, 127, 127, 127, 127, 113, -106, -128, 127, -128, 34, 127, -128, -54, -128, -128, 23, -123, 127, 127, 127, 35, -62, -128, -128, -128, 123, 113, 127, -128, -128, -128, -128, -68, -3, -91, -128, -128, -128, 20, -110, 127, 127, 103, 127, 9, 127, 127, 127, 127, 102, -3, -128, -76, -78, 127, -128, 127, 20, 127, 127, 26, 127, -128, -121, -128, -128, -128, -128, 127, 127, 127, 127, -15, 127, -128, 57, 127, -128, 127, 127, 127, 37, 18, -128, -128, -128, -128, 96, 80, 127, 127, -36, 127, -26, 127, -36, 58, 127, 37, 127, 127, 1, 23, -128, -78, -128, -128, -128, -128, -128, -128, 19, 127, -128, 127, -128, 127, -128, 100, 38, -128, 127, -128, -29, -97, -128, -128, -128, -128, -128, 107, -128, 127, 127, 127, 127, -128, -128, -55, -128, -47, -128, -128, -128, -128, -128, -30, -111, 127, 127, 127, -76, -128, -48, -128, -128, -128, -128, 127, 122, 127, 91, -57, -128, 127, -128, -128, -128, -59, -56, 122, -128, -128, -128, -128, -128, -108, -128, -128, -43, -128, 127, -128, 7, -128, -128, -17, -115, -128, 127, -82, 119, 102, 100, 66, -128, -10, 15, -128, 127, -128, 127, -87, 19, 127, 79, 127, -128, 20, -128, -126, 127, 127, 127, 65, 127, 127, 127, 127, 127, 127, 127, 56, 127, -82, 127, 127, -128, 127, -128, -128, -128, -126, 126, 127, 127, 127, 127, -128, 105, -128, 127, 127, 127, 127, -56, -128, -128, -128, 68, -128, -42, 127, -128, -87, -128, 12, -69, -128, 127, 127, 127, 86, 127, -128, -128, -128, -128, 77, -128, 89, 127, -61, 127, -128, 81, -128, -81, -128, 127, 20, 85, 127, 76, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -124, -128, -128, -128, -128, -128, -128, -128, 127, -128, -110, 127, -128, 127, -128, -128, -128, -128, -110, 45, 43, -26, -22, -128, 99, -128, 127, 127, 127, 127, 19, 127, 106, 127, 127, 127, 127, 108, -128, -128, -128, -128, -128, 116, -81, -128, -128, -128, -73, -128, 127, 127, 14, 127, -128, -2, -128, -128, -128, 112, 24, 127, 127, -27, 127, -15, -128, 28, -128, -128, -19, -128, 127, 125, 127, 127, 48, 127, -128, -31, -47, -128, 127, -4, 127, -128, 127, -128, -65, 127, 127, 127, 127, 127, 127, 108, 127, -128, 73, -128, -128, -128, -56, 112, 44, -21, -128, -128, -128, -128, -128, -128, -128, -123, 109, 127, 127, 127, 127, 127, 127, -75, 127, -91, -35, -26, -128, 117, 89, -128, -128, -128, -128, -128, 88, 127, -128, 11, -128, 25, -39, 127, 127, 127, 127, 127, 127, -128, 65, -38, -128, 127, -128, 57, -105, -128, -65, -128, -128, -128, 127, 5, 90, -89, -128, 125, -128, 127, 26, 28, -128, -128, -128, -128, -128, 48, -27, -41, 80, -128, 103, -109, 34, -128, 127, -128, 127, 6, 127, 127, -128, 96, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 103, 70, 52, 83, -114, -128, 127, -128, -35, -128, -128, -128, -128, -128, -124, -106, -128, 127, -128, 127, 127, 127, 120, -128, -29, 125, 27, 127, -128, -128, 90, 127, 127, 127, 69, -128, -128, -128, -128, -4, 127, 127, 127, -128, -128, -128, -128, -128, 117, -69, 127, 127, 127, 127, 82, -35, 127, -128, 127, -128, -128, -34, -128, 127, -128, 127, 5, 127, 94, 127, -59, -68, -128, -128, -30, -15, -85, -128, -128, -128, -41, -128, 127, -110, 127, -128, 127, -128, -128, -128, -128, 127, -13, 127, 127, 76, -128, -113, -128, -15, -56, -92, 127, -128, 127, 43, 127, 127, 110, -103, 127, -128, 127, 19, 127, 127, 97, 127, 25, 23, -128, -128, -128, -128, -106, -128, 127, -111, 127, 106, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -25, -128, 20, -128, -85, -99, -128, 45, -128, -107, -128, 127, -128, -70, 89, -128, 69, -43, 127, 127, 127, 39, 121, -128, 127, 86, 108, 104, 127, 127, 127, 127, 127, 127, 30, 102, -38, 92, 46, -128, -128, -121, -128, -62, 127, 116, 127, -128, 127, 127, -128, 26, -128, -128, -128, -55, 127, 127, 127, 127, 98, 127, 120, 88, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -49, -128, 127, -114, 127, 127, 127, 127, -85, -128, -128, -128, -128, -51, 127, -18, 127, -30, -34, -55, 127, -128, 73, -128, 62, 69, 127, 78, 127, 127, -128, 127, -93, -128, -74, -121, -128, 127, -128, 127, 127, 127, 127, -61, -24, 127, -128, 24, -128, -128, -128, 117, -128, -8, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -104, -128, -128, -128, -128, -128, -128, -128, -128, -43, 88, 127, 127, 6, 127, -128, -128, -128, 127, 9, 127, 117, 73, -128, -128, 127, 31, 127, -20, 127, 96, 110, -17, 127, 0, 7, -128, 127, 41, 127, 127, 127, 127, 127, -128, -128, -128, 13, -128, -61, -128, -128, -65, -128, 127, -2, 7, 127, 23, 127, 127, 127, 127, 127, 107, -31, -128, -128, -128, -128, -128, -128, -3, -128, 120, 127, 66, -109, -128, -128, -128, -128, -128, -18, 127, 127, 127, 127, -112, -78, -91, 127, 127, 127, 127, 127, 127, 44, 127, -128, -128, -128, -128, 127, -91, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 5, -128, 127, -128, 127, -119, -128, 39, -128, 127, -128, 127, -128, 127, -128, 56, 127, 2, 127, 127, 86, 127, -128, 127, 127, 127, 127, 127, 127, 83, 127, 107, 127, 95, 127, -115, 22, 44, 127, 127, -108, 127, -128, -128, -128, -100, 127, -31, 127, -128, -21, -128, -128, -128, -128, -3, -128, 124, -128, -94, -128, -126, -128, -122, 20, 127, -128, 127, 127, 127, 127, 127, 36, -26, -77, 89, -10, 127, 127, 127, 127, 127, 127, 127, 127, 88, 127, -14, 127, -90, 127, 98, 94, 127, -94, 127, -12, -72, -128, -128, -120, -128, 127, -96, 127, -128, 127, -24, 127, -48, 127, -128, 9, 72, 40, 127, 32, 127, -128, 127, 89, -128, 127, -128, 127, 127, 127, 127, 127, 127, 3, -128, -128, -128, -128, -87, -128, -128, 127, -29, 127, 127, 127, 127, -17, -128, -128, -128, -128, -128, -128, 66, -128, 114, 51, -128, -30, -128, -128, 123, 113, 127, -82, 127, 18, -128, -78, -128, 59, 127, -128, 127, 127, 91, 127, -128, 127, -128, -128, -128, -79, 103, 127, 127, 127, 127, -128, -128, -128, -128, 127, -106, -100, 117, -128, -34, -128, -128, -128, -128, 57, -32, 127, 127, 127, 127, 127, 127, 127, 127, 127, 17, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 58, 127, 127, 127, 104, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 49, -128, 127, 89, -128, 113, -51, -17, 127, -128, 127, -128, 127, -128, -72, -128, -128, 37, 88, 127, 127, 127, 127, 127, 61, 49, -75, -128, -128, -38, -128, -128, -128, -128, 79, -128, 53, -128, -128, -63, -128, 83, -128, -128, -18, -128, -128, -128, -128, 43, 127, 127, 127, 127, 127, 127, 127, 71, 127, -128, -128, -128, -128, 127, 127, 127, 127, -62, 127, 25, 24, -20, -43, -128, -128, -128, 127, 127, 127, 127, 127, -27, 127, -128, 122, -42, 127, 127, -128, 86, -11, 127, 127, 127, 127, 127, 80, 52, -128, 98, -128, 11, -128, 127, -128, 91, -128, -71, -128, -103, 49, -128, 127, 76, 127, 127, -128, -119, -124, -128, 127, 54, -128, 127, -128, -32, -128, 41, 127, 127, 127, -35, -128, -128, -128, 127, 127, 127, 127, -124, -128, -128, -128, 112, 127, 127, 127, 127, 45, -128, -128, -128, -128, -128, -8, -128, -128, 124, -128, -128, -128, -128, -128, -128, 53, 127, 104, 127, -128, 127, 7, -24, 76, 127, 56, 127, -1, -24, 127, 8, -128, 127, -54, 127, -128, -128, -128, -128, -128, -69, -128, 28, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -104, 82, -128, 127, -128, -72, 97, -128, -128, -128, 37, -115, 127, 127, 127, 127, 37, -128, 99, 46, -128, 23, -47, -1, -20, -128, -113, -128, -128, -128, 127, 3, -58, 127, -128, 127, 127, 46, 127, 127, -128, 127, -117, 127, 127, -128, 127, -128, -128, -128, -128, 4, -128, -128, -93, -128, 66, -128, -128, 127, -128, 127, -128, 127, -54, -104, 127, -128, 127, -128, -99, -128, 75, 127, 127, 127, 127, 127, 106, 127, 0, 127, -128, -128, -128, -128, 127, 127, -11, 127, -128, -102, -128, -128, 36, -128, -128, -4, -128, -128, -20, 111, -70, 127, -128, 127, 127, -46, 127, 10, 127, 127, -128, 127, 34, -128, 52, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 111, -128, 11, -73, -128, -128, -105, -128, -62, -103, -128, -77, -128, 40, 94, -19, 26, -128, -128, -128, -128, -128, -128, 43, -128, 60, 127, 127, -103, 127, -128, 127, -128, 124, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 25, -60, 127, -128, 127, -46, 10, -17, -128, -27, 102, -60, 127, -24, 54, 106, -128, 127, -128, 66, -111, -128, 127, 79, 127, -2, 127, 127, -78, 127, 127, 77, 127, 126, 127, -7, 127, -128, -128, -128, -128, -128, -1, -61, 8, 55, -128, -128, -19, -128, -128, 127, -128, 127, 96, 127, 127, 82, -56, 127, 21, 32, 89, -128, -77, 66, -108, 127, 127, 127, 127, -128, 127, -128, 88, -128, -128, 1, -128, -51, -72, 113, 127, -23, 127, -128, -128, 127, 127, 127, 127, 127, -128, -23, -128, -128, 85, -128, 127, -4, 76, -70, 127, 127, 116, 119, 127, -128, -55, -128, -15, 127, -128, 127, -128, -128, -128, -128, -128, 127, 115, 127, 127, -12, 127, 127, -128, 124, -9, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -19, 127, -128, 127, -87, 127, 127, 127, 127, 45, 127, -128, -32, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 64, 64, -35, 127, 127, -108, 127, -128, -93, -128, -128, -74, 127, -128, 127, -54, 36, -37, -128, -32, -128, 109, -128, 127, -128, 127, -112, -128, 127, -128, -121, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 91, 127, -64, -1, -86, -128, 127, -54, 127, 127, 127, 52, 9, 127, -24, 127, 127, 127, 31, 127, 61, -128, -128, -128, -128, 36, -128, -85, -96, -128, 85, -128, -128, -128, -128, -128, -128, -47, 100, -128, 127, -44, 127, -128, -128, -128, -128, 0, -128, 127, -128, 127, 127, 69, 127, 127, 127, 127, 127, 127, 127, 127, -108, -128, 127, -128, 127, -128, 127, 38, 127, -103, 127, 13, 102, 18, 127, -42, 89, -128, -128, 107, -128, 127, -83, -40, -128, -128, -54, -128, 127, 13, 127, 127, 127, 127, 127, 127, 2, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 59, 127, 127, 127, 5, 22, -109, -128, 86, 0, 127, -106, 5, -83, -113, -128, -11, -93, 127, 34, 87, 65, 109, -128, -82, -128, -128, -128, -128, -128, 46, -128, 36, 127, 127, 127, 127, -58, 127, -112, 127, -128, 127, -34, -93, -128, -128, -72, 127, 127, 124, 127, 127, 127, 127, 127, -81, 93, -128, 127, -109, 127, 127, 38, 127, -128, -47, -128, -87, -128, 127, -71, 119, 127, 69, 127, 127, 127, -128, 36, -128, 127, 95, -89, -128, -119, -128, -128, -74, 127, -128, 27, 127, 68, 127, 116, 127, 127, 127, -24, 127, -12, -128, 127, -128, 127, 99, 127, 127, 49, -51, -128, -128, -128, -128, 127, -76, 93, 65, -128, -128, -128, -75, -128, -128, 105, 4, 127, 127, 127, 127, 9, 127, -128, 127, 93, 103, 127, 8, 98, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 26, -128, -128, -128, -128, 102, -128, 56, 100, 127, 127, 127, 127, 44, 41, -128, 127, -128, 79, -128, -128, -90, -128, -128, -128, -128, 127, -128, 127, 127, 127, -51, -128, -128, 127, -114, 41, -64, -128, -102, -90, -69, -128, -128, -128, -128, 127, -21, -11, -128, -128, -128, -58, -123, 127, 127, 127, 127, 127, 127, 7, -62, 19, -128, -69, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -53, 127, -128, 127, -128, 127, 127, 127, 127, 36, 127, 38, 86, 46, -128, -128, -56, -73, 117, 127, 127, -128, 127, -128, -128, -128, 17, 79, 127, 127, 127, 127, 127, 127, 127, -12, -128, -128, -128, -128, 55, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -35, -128, 0, -61, -128, -128, -128, -128, 127, -128, -128, 127, -128, -26, -98, -128, 127, -128, -20, 99, -128, 115, -55, -99, -128, -57, -128, -128, 127, -128, -89, 127, -128, -74, -124, -126, -128, 127, -128, 76, 127, 88, 127, 127, 19, -128, -128, -128, -128, 127, 127, 127, -57, 5, -128, -128, -128, -128, -128, 8, -128, -128, -128, -128, -2, 127, 127, 127, -43, 127, -8, -59, -29, -14, -25, -128, -128, -128, 75, -128, -77, -128, 127, -59, 127, -7, 127, 115, 127, 4, 127, 23, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -119, 127, -9, -128, -54, 25, -128, 127, -128, 127, -128, 61, -127, -128, -128, -128, -38, 127, -128, 127, -128, 127, -10, -128, 127, -43, 127, 127, 127, 127, 100, -7, -128, -113, 14, -128, 39, -57, -25, 127, -128, 127, -128, -3, -128, -128, -128, -128, -31, -128, 127, 97, 127, 127, 127, 127, 127, -32, 127, 127, -128, 127, -104, 127, -128, -128, 112, -128, 127, -30, 127, -99, 127, -128, -128, -128, -128, -105, -128, 127, -6, 127, -128, -128, -128, -128, -97, 82, 127, -102, 127, 96, 127, 127, 127, 127, 127, -52, 127, -128, -128, -128, -128, 127, -128, 127, -123, 127, 127, 111, 127, 103, -64, -128, -128, 127, 26, 127, 127, 127, -36, -44, 9, 72, -83, 127, -128, -6, -128, 127, -128, -21, -128, -128, -43, -128, 127, -128, -128, -128, -107, 49, 127, 127, 127, -17, -128, -128, -128, 42, -128, 127, -128, 87, -128, -128, 127, 110, -45, -59, -128, -128, 127, -128, 39, 20, -128, -128, -128, 127, -54, 127, 127, 103, 127, 127, 127, 127, 127, 127, 82, -128, 127, -128, -44, -110, -128, 127, -128, 9, 127, -128, 127, -128, -128, 127, -128, 127, 127, -31, 127, -128, 127, -128, 85, 127, 127, 127, 127, 32, -80, 127, 120, 9, 127, 127, 20, 127, -61, 92, -95, -128, -15, -128, 127, 127, 127, 127, 127, -56, -54, -128, 49, -22, 127, 127, 127, -128, 127, -128, 127, -52, 127, 15, 127, 121, 127, 127, 59, 127, -83, 127, 127, 81, 127, -128, -51, -128, -128, -77, -100, 127, -128, 127, 102, 127, -128, 127, 65, 127, -42, 93, -128, -128, -128, -123, 127, 127, 127, 127, 44, -128, -126, -128, -24, 127, -128, 127, 127, -128, 127, -58, 127, 127, -128, -72, -112, 24, 127, 127, 127, 127, 127, 127, 127, 127, 31, -40, -128, -128, 89, -128, 127, -73, 127, -108, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -53, 127, -128, 127, 127, -38, 127, 113, 127, -49, -113, -62, 127, 43, 127, 127, 14, 62, -128, 30, -128, -103, 127, 127, 127, 127, 127, 34, 127, -128, 127, -128, -59, -128, 127, -128, 127, 17, 127, 127, 127, 127, -128, -65, -128, -128, -128, -128, -128, -2, 40, 127, -91, 35, -128, -128, -102, 86, 127, 127, 81, 127, -63, -64, 0, 120, -128, -98, -128, -47, -128, 85, 127, 127, 127, 127, 127, 127, 37, 127, 120, 127, -128, 127, -120, -27, -28, 127, 127, 127, 127, -128, 127, -128, 51, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -111, -128, -128, -128, -4, -128, -128, -128, -128, -74, -126, 127, -128, 0, -51, -128, -128, -128, 120, -128, 123, 127, -120, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 69, -123, -128, -128, -128, -128, -128, -93, 127, 127, 127, 91, 48, -128, -119, -128, 98, 127, 74, 127, -117, 75, 34, -128, 108, 89, 53, 127, 127, -128, -71, -128, -68, -120, 127, 127, 127, 127, 127, -128, -47, -128, -128, -128, -128, -128, 127, 127, 127, -128, 35, -128, -128, -128, 3, -98, -49, -43, -128, 127, -128, 127, -128, -61, -128, -128, -128, -31, 127, -128, 80, -128, -128, -128, -128, -94, -115, -85, 127, 127, 127, -128, -128, 127, -128, 127, 92, 127, 127, -128, 127, -128, -117, -128, -88, 127, -128, 127, -128, -96, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 9, 127, 19, -128, 90, 87, -128, 127, -128, 45, -128, -10, -128, 127, -128, 127, -128, 104, 127, -20, 127, 119, 11, 127, -128, 127, 127, -128, 127, -128, 127, -64, -128, 73, -5, 64, 127, 127, 127, 127, -128, 2, -128, 127, -128, 127, -128, 127, 127, -85, 127, -128, -117, -8, -128, -21, -9, -22, -128, -128, -128, 127, -128, -40, 87, -128, 20, -128, 127, 127, 60, 95, -128, -128, -128, 127, 127, 127, -91, 127, -128, 7, -128, 97, 127, -128, 127, -128, 127, -128, 127, -107, -128, -24, -128, -128, 127, 56, 127, 127, -21, -35, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 112, -128, 127, 5, 127, 125, -128, -128, -128, -128, 127, -30, 127, -90, -128, -108, -128, -128, -128, -128, 18, 79, -49, 127, -128, 44, 108, 36, 127, 127, 127, 127, 127, -63, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -89, 127, -128, -82, -128, 127, 127, 87, 127, 72, 126, 116, 34, -13, -15, -128, -128, -127, 127, 127, 127, 91, 86, -109, 127, -128, -85, 127, -128, 127, 62, 127, 127, 86, 127, 127, -14, 127, -128, -128, -128, -128, -128, -128, 0, -128, 127, 125, 127, 127, 127, 127, 74, -128, -128, -128, -128, -85, -128, -64, -128, -128, -128, -128, -128, -128, -128, -128, -128, -14, 93, 127, 32, 127, -52, 127, 66, 127, 127, 18, -102, -128, -128, -128, -128, 70, -128, 127, -43, 127, 127, 125, 127, 127, 127, -41, 127, -128, 61, -128, 127, 82, 127, 127, -5, 127, -29, -128, 110, -128, -106, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 37, 127, 127, 98, 127, 14, 47, -104, 71, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 5, 127, -128, -128, -128, -128, -128, 42, -128, 127, 127, 127, 127, 127, -3, -128, -128, -126, 12, 127, -52, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 78, -128, 11, -128, -128, -128, -128, 7, -128, -128, -128, -128, -64, -108, -128, -90, -95, -15, 5, 100, 120, 127, 127, -128, -128, 72, -128, -1, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -106, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 76, -128, 127, -128, 82, -128, -128, -2, -128, -126, -128, -20, -128, 73, -27, 127, -128, 127, -128, -128, 17, -128, 127, -128, 112, -85, 127, -128, 127, 127, 96, 127, -107, -128, -72, -128, -128, 52, 127, 127, 127, 27, 127, -127, 127, -128, -36, -128, -104, -128, 127, -75, 127, 127, 127, -120, -128, -128, -128, -103, 0, 127, 64, -105, -128, -128, -105, 86, 127, 38, 127, -88, 112, -8, 127, 0, 127, -128, 127, -128, -128, -128, -128, -128, -128, -91, -128, -7, 127, 127, 127, 60, -66, -66, -128, 37, 127, -128, 81, -119, 56, -99, 127, -128, 26, -128, -128, -70, -128, 127, -69, -11, -34, -128, -128, -68, -52, 103, 127, -128, -128, -128, -128, 127, 127, 127, 112, -17, -128, -128, -128, -128, -128, -128, -128, -128, 90, -128, 127, 127, 127, 127, -45, -24, -128, -128, -111, 127, 127, 127, 127, -128, -68, -128, -112, -128, 57, -128, 127, 127, 127, 127, -59, -128, -128, 52, -128, 127, -128, 127, -115, 127, -6, -128, -128, 127, -128, -94, 127, -128, 127, 57, 127, 127, 127, 127, -128, 127, -128, 127, -112, 127, 54, -128, -128, -128, -51, 32, 127, 127, 127, 127, 14, 127, -128, -11, -128, -31, 40, 127, -4, 127, -88, 127, 11, -9, 86, -79, -128, -128, -128, -128, -128, -128, -128, -91, 71, -12, 127, -22, 127, -128, -96, 48, -128, 79, 117, -128, -79, -128, 127, 127, 127, 127, 15, 127, -128, -128, -128, -100, -128, -92, -10, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 112, 127, 127, 127, 127, 127, 127, -30, -30, 127, -36, 127, 125, 127, -128, 127, 5, 26, 127, -124, 47, -115, -128, 127, -128, -72, -128, -128, 127, -128, 127, -128, 73, -128, -128, 53, 27, 127, 77, 127, 22, 127, 127, -128, 70, -128, -128, 127, -128, 127, 99, -57, -6, -128, -128, -128, 44, 29, 21, -128, -128, 72, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 51, 127, -128, -128, -128, -128, -20, 92, 127, 127, 127, -128, 127, -128, 127, 114, -54, 127, -128, -124, -10, 127, 127, 127, 57, 89, 127, -128, 127, -128, -8, -128, -128, -128, -128, -128, -128, -128, -128, -11, 18, 92, 21, 127, -128, -128, -128, 49, -19, 127, 127, -88, 6, -128, -59, -80, -2, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 47, -128, 80, -128, 120, 122, 127, 57, 127, -128, -128, -95, -128, 97, -128, 127, -128, 127, 7, 127, 127, 127, -128, 127, -128, 127, -126, -60, 4, -128, -128, -128, -128, -128, -128, -128, -128, -128, 18, -60, -128, 127, -128, 127, -128, -126, 105, 77, 127, 127, -128, 127, -83, 83, 127, 124, 127, 127, 127, 127, 112, -128, -128, -128, 38, -2, 127, -52, 23, -128, -128, -128, 82, -128, -128, -128, 30, -64, 127, -22, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 25, 127, 127, 127, 127, 92, -3, -52, -128, 127, 41, 127, 127, -128, 127, -3, 127, 127, 127, 127, 127, -51, -128, -128, -128, -128, -128, -128, -128, 8, -120, 127, 127, 124, -128, -128, -128, -128, -128, -104, -128, -110, -27, -128, 127, -121, 124, -111, -128, -128, -128, -128, -19, -93, 32, 127, -128, -7, -128, -128, -128, -128, -14, -128, 127, 127, 127, 127, -128, 127, -128, 30, -24, -128, 127, -9, 127, 127, 127, -128, 127, 127, -128, 127, -128, -56, -83, -103, 56, 127, 127, 104, 127, 127, 127, 127, 100, 127, 127, -128, -128, -31, -128, 104, -128, -128, 127, 1, 127, -128, -25, 86, 127, 127, 127, 127, 127, 127, 36, 106, -128, -21, -128, -79, -29, 10, -112, -128, -128, 65, -99, 127, 127, 127, -11, -128, -65, -128, -128, 46, 7, 127, -54, -59, -128, -128, -128, -128, -128, -128, -119, 127, -128, 127, -128, -128, 127, -128, 127, 127, 56, 127, -128, 36, -128, -120, -128, -128, -128, -123, -128, -128, 125, -128, -128, 32, -128, 127, -128, 37, 127, -128, 127, -128, 127, -128, -128, -128, -64, 108, 127, -99, 119, -15, -128, 127, -123, 127, 127, 127, 5, 127, -128, 127, 127, -128, 127, -128, 127, -76, -47, 127, -128, 127, -128, 70, -13, -128, -128, 127, -128, 127, -128, 127, -128, 127, -116, 127, -122, -17, -128, -122, -128, -128, 100, -128, 127, -128, 127, 112, 127, 37, 127, -55, 47, 13, -128, -128, 127, -128, 127, -51, 127, 19, -128, -126, -128, -128, -5, -11, 127, 127, 127, 127, -128, -42, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 97, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, -85, 127, -54, 127, 127, -128, 127, -86, 127, -52, -128, -128, 127, 127, 127, 127, 127, -73, 127, -128, -27, 86, -128, -128, 119, 126, 127, 51, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -57, 125, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -105, 127, 43, 127, -128, 127, -128, 44, -128, -49, -92, -128, -128, -128, -128, -1, -128, 127, -128, 127, -128, 49, 127, 127, 127, 61, 127, -29, -128, -128, -128, -128, 127, 91, 127, 127, -123, -128, -128, -128, 45, 127, 127, 127, 127, -114, -81, -128, 127, 127, 127, 127, 45, 127, 5, -73, 127, -128, 127, -42, 127, 127, 127, -7, 127, 127, 127, 127, 127, -126, -128, -128, 73, 127, 127, 127, 127, 97, 29, 127, 97, 127, -128, 127, -2, -128, -58, -128, -128, 127, -56, 127, 127, 127, 96, -128, -128, -128, -128, -128, 76, 127, 127, 127, 127, 127, 127, 40, -22, -128, -128, -126, -56, 127, 127, 127, 127, 95, 127, 127, -115, 88, -128, -128, -128, -128, -128, -47, -46, -128, 77, -128, 127, 127, 19, 127, -22, 127, 127, 127, 127, 127, -122, -128, -128, -128, -97, 17, 88, 127, -128, 115, -128, -45, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -3, -117, 127, -128, 127, -128, -47, -128, 127, 123, -128, -89, -128, -128, -128, 127, -58, 127, -128, 111, -128, -128, 127, -128, 127, 47, 127, 127, 127, -114, 127, 64, -128, -128, -128, -128, -128, -128, -45, 127, 121, 112, -71, -128, 103, -128, 127, -128, -1, 114, -128, 127, -128, -128, 54, -128, 42, 127, -113, 127, -128, 127, -128, 127, -78, 127, -128, 127, -46, 127, -14, 127, -126, 105, -128, 127, -128, 20, -63, 127, 65, -124, 15, -128, 127, -128, -80, -128, 103, 78, 127, 127, -62, 127, -128, 127, 62, 127, 113, 127, -128, -113, -128, -128, -128, -128, -128, 127, -45, 127, 127, -12, 127, -128, 90, -128, 127, 127, -24, 127, -128, -128, -32, -128, 46, 127, -10, 127, 127, 127, 127, 127, 127, 127, 127, 127, -102, 127, -128, -128, 127, -128, 68, 43, -115, -87, -128, -62, 95, 79, -128, 127, -128, 127, 117, 113, 127, 36, 14, 2, -128, -2, -128, -128, -128, -128, 127, 79, 127, 27, -128, -110, -128, -123, -79, 127, 127, 127, 127, 127, 127, -63, -128, -128, -128, -128, -128, 39, 127, 127, 127, 127, 127, 102, 96, -6, -42, 127, -128, 88, 73, -112, 127, -64, -7, -65, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 79, -2, 127, -128, -128, 89, -128, 127, -39, 127, 127, 127, -128, 65, -128, -128, -35, -128, 127, -87, 127, -128, 127, -128, 127, 46, 127, 127, -72, -30, -128, -128, 127, -128, 127, 127, 127, 127, 46, -128, -99, -109, -88, 112, 127, -128, 127, -49, 127, 62, 127, -102, -128, -128, -128, -52, -128, 127, -128, -11, 127, -128, 127, 127, 127, 127, 2, 104, 22, -13, 113, 115, -128, -108, -110, -99, 127, 54, 127, -128, -128, -128, 36, -128, -128, 125, -128, 127, 127, 127, 127, 127, 127, 106, -100, -128, -128, -128, 97, 127, -77, 98, 127, -128, 127, -128, 1, -68, -128, -128, -23, -128, 127, 127, -91, 56, -117, -99, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 6, -21, -128, 127, 12, 127, 127, -52, 127, -117, -128, -10, -128, -89, -128, -18, -128, -128, 127, -128, 127, -128, 127, 127, 127, 34, 127, 109, -128, 127, -128, 127, 127, -65, -128, 54, -128, -128, -128, -85, -128, -72, -36, 127, 127, 27, 127, -128, 127, -128, -128, -128, -128, -128, -27, 127, -44, 127, 20, -128, -59, -11, -77, 30, 127, 127, 127, 25, -128, -128, -128, -128, 127, 114, 127, 127, 127, 127, 127, 61, 127, -128, -128, -66, -128, 99, -128, 32, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 17, 127, 127, 76, -128, -109, -128, -128, 2, -128, 127, 127, 127, 127, -128, 127, -128, 110, -128, -128, 127, -128, -4, 127, 97, 127, -128, -89, -128, 127, 49, 127, 127, 127, 114, 121, -128, 127, -128, -128, -128, 32, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -62, -12, 127, -128, 127, -111, 14, 127, 127, 127, 75, 127, -128, -128, -34, -128, 27, -56, 108, -112, 127, 127, 73, 127, -128, 127, -128, 31, 127, 127, 127, -128, -128, -128, -128, -128, -128, 81, -128, -115, 127, 127, 99, 127, -128, 27, -128, -128, -128, -23, -128, -128, 18, -128, 127, 17, 127, 127, 127, -128, 121, -128, 71, -128, 127, 39, 127, -25, 127, 91, -128, -128, -18, -128, -128, 127, -128, 127, -127, 127, -128, 26, -128, -128, -112, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, 89, -128, -128, -42, -58, 127, 127, 127, 88, -128, -128, -128, -128, 3, -28, 13, -128, -105, 19, -128, 127, -53, 127, -103, 106, -128, -126, -128, -102, -86, -128, -98, -128, -128, -128, -128, -128, -128, -128, -10, 102, -32, 127, -24, -128, -54, -128, -128, -128, -128, -128, -29, 127, 127, 127, 127, 127, 109, -128, -63, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 59, 4, -128, -126, -128, 64, 127, 127, 127, 105, -128, -103, -128, -126, 74, -121, 127, 127, 127, 127, 127, 127, 127, 127, -1, 127, 127, 127, 127, 127, -56, 125, 88, -66, 127, 127, 59, -79, 42, -128, 72, -128, 60, -126, 36, -65, 3, -128, -95, -128, 0, 127, 127, 127, 127, 121, 127, -128, 43, -128, -128, -128, 127, 114, 127, 127, -97, 127, -111, 40, -128, -128, -128, 37, -128, -128, -61, -3, 127, 122, 127, 127, -2, -128, -111, -128, -128, 127, -128, 127, -128, 93, 127, 127, 127, 127, 127, -95, 109, 127, -128, 127, -128, 127, 100, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 36, -56, 127, -128, 127, -128, 127, -4, 127, 127, 108, 127, -128, 110, -128, -91, 127, 127, 127, 73, -4, -80, 66, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 68, 127, 127, 5, 127, 127, 127, 127, 88, 127, 127, -128, -128, -128, 93, -128, 11, 127, 39, 127, 127, 127, 127, 127, 127, -26, -128, -128, -128, -128, -128, 127, 65, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 10, 105, 61, 127, -128, 127, -128, 30, -41, -77, 94, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 110, 127, 127, 127, 37, -128, -103, -128, -128, -44, 127, 127, 127, 127, 127, 127, 79, 127, -128, 127, -63, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 28, -128, -128, -128, -128, -128, 124, 127, 127, 127, 127, 127, 80, -128, 127, -128, 127, -128, 74, 74, -111, 127, 127, 127, 127, -18, 41, 127, 21, 127, -128, 127, -64, -12, 127, -128, -37, -128, -128, 127, -128, 0, -128, -128, 127, -128, 105, -128, -127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 40, -51, -128, 22, -128, 127, -128, 127, 106, 127, 127, -128, 127, -128, 126, 127, 127, 127, 127, -128, -98, -128, 74, -128, 28, -128, 127, 29, 113, -128, 127, -128, 127, -11, 127, 127, 127, 120, 127, -128, -22, -58, 127, 127, 127, 127, 127, 127, -128, 71, -128, -104, -128, -128, 86, -128, -128, -128, -128, 64, 97, 103, 127, -128, 62, -128, 127, -128, -64, -128, -128, -54, -128, 127, -120, 127, 117, 125, 127, 127, 70, 127, -15, 127, -53, -128, -128, 14, -128, 127, 28, 73, -60, -68, 127, 127, 127, 127, 9, 127, -72, -73, -64, -128, -128, -128, 127, 127, 34, 127, -28, -128, 11, -49, 127, -128, 14, -82, 78, 4, 127, 127, 45, 127, -8, 127, -128, -45, -128, -15, -112, -128, 0, -128, 5, -128, 127, -3, 121, -124, -106, -128, -128, 127, 127, 127, -126, 125, 124, -128, 25, -7, -128, 127, 51, 77, 127, -128, -128, -128, -128, -128, -128, -83, -128, -56, 26, 76, 53, 127, 127, -76, 97, -128, 11, -128, -128, 13, 127, 27, 127, -128, 127, -128, -127, -34, 110, 127, 42, 127, 127, 127, -89, -128, 0, -128, 127, -19, 112, 127, 127, -7, 127, 66, -36, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 34, 57, -128, -128, 127, -128, 127, 41, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -53, 127, -128, 30, -128, -128, -128, -128, -128, -128, -85, -74, 127, -128, 127, -56, 127, 127, 127, -88, 64, -128, -128, -30, -128, 25, 127, -128, 127, 14, 127, 126, -128, 127, -128, 127, -54, -52, -128, -128, -128, 36, 127, 127, 127, 127, -128, -128, -58, -91, 127, -55, 127, -128, -128, -128, -21, -88, -61, -47, -77, 107, 127, 127, 127, 127, 127, -52, 2, -128, -128, -128, -128, -128, -128, 115, -105, -3, -128, -128, 57, -128, -64, 104, -128, 127, -128, 127, 0, -128, 127, -128, 127, 127, 127, 127, 127, -80, -128, -90, -128, 63, -128, 89, -46, -81, 127, 127, 127, 72, 62, 45, 12, 12, -128, 20, -68, 127, 38, 127, -128, 127, -128, -28, -128, -128, -128, -128, -128, -128, 127, -57, 127, 127, 127, 127, -121, 127, -128, -31, -128, 127, -128, -128, -128, -128, -109, -38, -93, -128, -128, -128, -128, 127, -1, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 105, 127, -128, 127, -6, 127, 94, 127, -31, 127, -128, 108, -128, -128, -128, -128, -128, 106, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -116, 127, 127, 127, 6, 48, -128, 127, -128, -119, 127, -128, 127, -128, -31, 127, -128, 127, -128, 82, -80, -128, -128, -128, -128, -128, -105, 127, 127, 127, 127, 127, 83, 127, -128, 127, -128, 127, 112, -128, 127, -128, 127, -128, 37, -47, -128, -11, 127, 127, 127, -1, 114, -128, -128, -128, -128, -128, 127, 127, 127, 76, -104, -128, -128, -20, -73, -90, 127, 127, 127, 127, -128, -102, -128, -128, -128, 51, 127, 127, 10, 31, -128, -128, -55, -128, -128, -128, -128, -128, 124, 127, 127, 127, -20, -52, -128, -128, -128, -128, -128, -80, 127, 127, 127, 127, 127, 12, -128, -128, -128, -128, 127, 127, 127, 28, 127, -128, 127, -128, 127, 85, -80, 127, -128, 121, -128, -128, -128, -128, -128, 99, -128, 127, -128, 127, 127, 127, 127, 127, -53, -114, -37, 127, -15, 76, 109, -128, 127, -11, -7, 127, -128, -83, -128, -9, -128, 42, 127, -128, 127, -128, 127, -34, -128, -25, -128, -128, -128, -65, -128, -128, -128, -128, -128, -128, -68, 43, 127, 127, 21, 87, -83, 127, 127, 127, -66, -17, -128, -128, -128, 105, 127, -21, 127, -79, -128, 127, -128, 127, 127, -53, 127, -128, 127, -128, -128, -36, -128, 127, 93, 86, 127, -115, 127, 29, 51, 127, 127, 127, 127, 64, 51, 98, 106, 127, -90, 127, 127, -77, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 55, 43, 15, -128, -128, -128, -128, 72, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -73, -128, -128, -94, 127, 22, 127, -128, -128, -128, -128, -58, 127, 127, 127, 127, 127, -23, -128, 27, -128, 127, -128, -128, -128, -128, 123, -128, 127, 127, 26, 127, -128, -108, -128, -119, -128, -128, 127, -5, 51, -8, 4, -128, 48, -128, 31, 127, -41, -128, 24, -88, -128, 127, 127, 127, -87, -128, -56, -128, -71, 127, 127, 127, 127, 127, 127, 127, 127, -85, -128, -82, -128, 127, 127, 58, 127, -128, 127, -128, -128, -128, -128, -128, 127, -47, 127, 14, 127, -128, 127, -66, -102, -78, -128, -128, -128, 29, -102, 127, -128, 127, -128, 127, -128, -128, -128, -14, -128, 127, 61, 127, -100, 127, -107, 127, 127, -128, 127, -128, -128, 79, -128, -128, 127, -128, -21, -128, -128, -100, -128, -128, -128, -128, -128, -39, -128, 127, -4, 127, -80, -128, 127, -128, 127, -128, 127, -128, -25, -128, 75, 127, 127, 127, 127, 127, 127, 15, 96, -128, -128, -114, -128, 127, -34, -15, -91, -128, 127, -128, 127, 127, 127, 127, -92, 103, -128, -91, -128, -128, 54, -128, 121, -24, 18, 77, -128, 15, -128, 127, 127, 91, 127, -61, -57, -128, -128, -61, -128, -128, -128, 42, -128, -41, -78, -128, -128, -128, 69, 127, 127, 127, -128, -128, -128, -13, 61, 127, 127, 127, -123, -128, -128, -128, -128, -128, -128, -128, -128, 122, 98, 127, 127, 127, 127, -128, 59, -128, -128, 127, -21, 127, 127, -128, 127, -128, 127, -128, 127, 127, 4, 127, -128, -128, -117, 127, 127, 39, -55, -94, 36, 34, 127, 127, -128, -128, -128, -128, -128, -128, -128, -119, -128, 36, -66, -52, -119, -128, -128, -5, 127, 127, 127, 127, 127, 25, 127, 127, -128, 127, -128, -128, -128, -128, 127, 30, 127, 127, -128, -111, -128, -128, -128, -128, 52, 127, -45, 127, -128, 127, -128, 127, -128, 28, -128, -119, -128, 77, -64, 116, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, -104, -128, 127, 108, 127, 127, 62, 127, -128, 81, -128, 13, -128, -128, 127, -31, 114, -128, 127, -128, 22, 127, 127, 127, -128, 102, -111, -128, -128, -128, -128, -25, 31, 127, -128, 126, -128, -128, -128, 76, 127, 127, 127, 127, 19, 127, -60, 4, 127, -128, 7, -128, -128, -128, -128, -94, -128, -60, -128, 1, 127, 127, 127, 18, -128, -128, -128, -128, -103, -43, 127, -128, 127, -128, 127, -128, 71, 105, -128, 127, 19, 61, 9, 127, -127, -126, -20, -128, 8, -128, -87, -128, -128, 69, 105, 127, 127, 127, 127, -128, -38, -128, -32, -128, -51, 127, 127, 127, 127, 127, 127, -36, -128, -128, -128, -128, -46, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 48, 127, -47, 127, 127, -128, 127, -128, 3, -87, 127, 7, 127, -128, 53, -128, -128, -112, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 90, 127, -128, 127, -74, 127, 12, -128, 127, -128, 4, -128, -128, 127, -128, -128, 44, -128, -128, -128, -128, -17, -79, 127, 127, 114, 127, -128, 127, 85, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -96, -128, -34, 31, 15, 127, -128, 127, -128, 41, -128, 127, -39, 127, 127, -128, 127, -128, -1, -38, 79, 36, 127, -99, 127, -128, -124, 127, -128, 127, -128, 108, -128, 127, 127, 79, -1, -128, -128, -15, -128, 127, 127, -23, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 75, 99, 127, 127, -108, 127, -24, 111, 127, 127, 127, 127, 127, 4, 127, -8, 56, 127, -128, 103, 127, -128, 127, 40, 82, 99, 105, -128, 104, -128, 127, -90, 127, 112, 127, 127, 127, 127, 127, 127, -122, 127, 83, 127, 127, -13, 59, 127, -128, 127, 127, 19, 127, -128, -82, 42, -128, 127, -128, -10, 127, -23, -112, 127, -128, 120, -128, 24, -128, -128, -128, -128, -70, -35, 127, 127, 127, 127, 127, -128, -93, -128, -128, -128, -128, -128, -128, 37, 127, 109, 127, -114, 94, 52, -128, 114, -51, -128, -43, -66, -91, 127, -128, 127, -128, 127, 127, -128, 127, -128, -60, -128, -128, -71, -48, 127, 36, 127, 127, 127, 127, 20, 127, -115, -128, -128, -128, 6, -35, 127, 15, -69, 78, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 12, 127, 74, 80, 2, 5, 127, -56, 127, -57, 49, -128, 127, 103, -39, 127, -128, 83, 127, 127, 127, 127, 127, -128, 29, -128, 32, 127, 127, 127, 127, -128, -128, -128, -128, -128, 82, 127, 127, 73, -127, -128, -128, -128, -128, 53, -128, 127, -128, 127, -128, 127, -128, 127, -128, -89, 26, -128, 127, 127, 78, 127, 127, 127, -111, 127, -128, -85, -128, -128, -128, -128, -128, -128, 38, -128, 127, 127, 127, 127, 127, 75, 42, 102, 127, 52, 77, 127, -128, 127, -24, 127, -128, -107, -128, -128, -128, -39, -128, 127, -128, -128, -128, -128, -128, 57, 34, 127, -128, 127, 63, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 55, 42, -128, -128, -128, -128, -63, -128, 53, -128, -128, -128, -6, -49, 127, 127, 127, -128, 127, -128, -128, -1, 27, 127, 76, 69, 40, 127, 127, 127, 98, -17, 127, 29, 127, -96, 127, -128, -128, -128, -128, -128, -128, -128, -128, -64, -128, -128, -128, -128, -128, -57, -128, -128, 127, -85, 127, 127, -12, 127, -128, -128, -128, 127, -29, 127, -25, -128, -53, -128, 80, -128, 122, -128, -14, -128, -56, -128, -128, -128, 46, -116, 127, -112, -128, -128, -128, -51, 127, 0, 127, -128, 127, 73, -7, 97, -128, -128, -128, -128, -128, 127, -8, 127, -128, 39, -128, -128, -128, -57, -128, 127, -128, -95, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -95, 52, -113, 127, 98, 127, -128, -128, -128, -128, -128, 127, 127, 119, 56, -98, 90, -128, 127, 127, -128, -128, -128, 65, 103, -128, 127, -128, 127, -128, -128, -128, -128, -128, 103, -128, -105, -128, 82, -128, 127, 127, 127, 52, 127, 127, 127, 127, -128, 127, -128, -128, -44, -128, 127, -75, -114, -128, -128, -128, -128, -128, 5, -128, 127, -128, -95, 68, -128, 9, -128, 58, -128, -128, 127, -20, 127, 127, 127, 109, -104, -128, -128, -128, -128, -128, 11, -128, -128, -53, -128, -128, -128, -128, 49, -23, 127, 127, -112, -128, -128, -128, 127, 127, 41, 127, -128, -58, -128, -70, 127, -42, -107, -127, -128, -128, -100, -128, 8, -15, 13, 114, 52, 127, -128, 127, -115, -38, 127, 119, 127, 127, -128, 127, 22, 127, 127, 61, 127, -44, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -38, -128, -128, -128, -128, -102, -65, 127, 102, 102, 47, -27, -128, 127, 85, 87, 104, 127, -128, 127, -105, 119, 127, -25, 71, -128, 127, -128, -128, -128, -59, 127, 127, 127, 127, 127, 83, 62, -128, -128, -93, -128, 127, -128, -55, -128, -37, -128, -81, 69, 85, -41, -128, -22, -128, -128, 64, -128, -128, -128, -128, -128, -128, -128, 127, 95, 127, 7, -128, -128, -128, -128, -7, 86, -48, 127, -128, 127, -128, 127, 34, 120, 127, -39, 127, 127, -128, 127, 107, 127, 127, -25, 127, 127, 127, 127, 127, 127, 21, -128, -128, -128, -128, -18, -128, -128, 87, -128, 127, -128, -66, -128, -108, -128, -128, 127, -46, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 42, -128, -92, -128, 29, 127, 127, 127, 127, 14, -128, -62, -128, 77, 123, 127, 127, -80, -128, -128, -128, -128, -128, 63, 127, 127, 127, 127, 127, 103, -8, 127, 127, 34, -128, 15, -128, -128, -128, -128, -28, -128, 40, 86, -128, -128, -128, -128, 89, 69, 127, 62, 77, -69, -128, 127, -128, -128, 127, -128, 127, -128, 127, -77, -94, -128, 127, -128, -123, 127, -128, -128, 127, -128, 127, -128, 112, -128, -114, -128, 44, -128, 127, -124, 127, 127, 13, 127, -32, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -96, -128, -43, -128, -128, 91, 127, 127, 127, -12, 96, -95, -128, -41, -128, 90, -128, 127, -128, 127, -128, 34, -128, 29, 127, 127, 113, 127, -128, 127, -15, 127, 11, 1, -128, -128, -128, -128, 127, -93, 127, 127, 127, -74, 127, -128, 127, -128, 122, -128, -112, -78, 127, 127, 127, 127, 123, -128, -128, -128, 4, 127, 127, 127, -5, 127, -128, 127, -128, 127, 127, 94, 123, -77, 127, -77, 127, 127, -128, -32, -128, -128, -128, -122, 11, -128, 127, -110, 127, 127, 127, 117, -43, -128, -52, 21, 105, 127, 127, 64, 127, -128, -128, -128, 127, -128, 127, -128, 127, 22, -74, -4, 15, -128, -128, -128, -128, 90, -128, 127, 115, -74, 104, -55, -52, 127, 77, 4, -128, -128, -128, -65, -128, -41, -128, 127, -128, 113, 127, 127, 127, 127, 127, 13, 127, -128, -128, -128, -47, 127, -97, -36, -122, 127, -128, 127, -128, -42, -128, -128, 112, -128, -128, -128, -6, -128, -128, -128, -128, -128, -128, -128, -128, -15, -128, 127, -77, 127, 66, -18, -128, 127, 18, 127, -62, -126, -60, -128, 96, -18, 127, 127, 127, 127, 127, 127, 127, 127, 127, -65, -128, -128, -128, 127, 0, 127, 127, 127, -128, 127, -87, 127, 64, -113, -110, -128, 127, 127, 83, 127, 109, -128, -128, -128, -128, -128, -128, -75, 127, 127, 55, 127, -128, -48, -128, 10, 127, 127, 127, 89, 106, 30, -128, -32, -70, -128, -128, -128, -2, -128, -6, -128, 56, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 56, 127, 127, -128, 127, 119, 127, 127, 127, -85, -128, -128, -77, -128, 127, -42, -72, 127, -128, -128, -128, -128, -128, -93, -96, -128, 98, -128, -27, 127, 64, -44, -98, -12, -128, 127, -128, -26, 127, -128, -128, -128, -128, -7, 127, -128, 127, -128, 127, 51, 122, 127, 127, 127, -88, 116, -88, 47, 95, 127, 127, 127, -116, 122, 114, -128, -128, 24, -128, -128, 127, -128, 127, -128, -26, 127, -68, -25, 62, 127, -128, 127, -128, 127, -128, 66, 66, 127, 127, 127, 109, -128, 55, -128, -128, -128, -12, 127, -128, 127, -70, 99, -128, -128, -39, -128, 127, 75, 127, 108, 127, -128, -128, -128, -128, 126, -64, 127, 127, 127, 127, 36, 32, 87, 126, 127, 127, 127, 127, -128, -128, -128, -128, -106, -76, 127, -41, -68, 127, 127, 127, 127, 127, 127, -95, -5, 97, 59, 127, 127, -36, 95, 73, 127, 127, 127, -30, -85, -128, 127, -128, 127, -128, 30, -57, -128, 115, -128, -128, -90, -128, 127, 127, -65, -109, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -80, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 104, 127, -128, 127, 83, 127, 127, 127, 127, 74, 127, 127, -114, 127, -128, -128, -99, -128, -27, -128, -4, -128, -128, 46, -53, -22, 31, 127, 127, 127, 127, 127, 127, 119, 127, -128, 127, -111, -128, -128, -128, 127, -128, 127, 127, 127, 77, -22, -128, 127, -128, 123, 127, -128, 127, -80, 127, 53, -128, -107, -128, -40, -128, 127, 65, -128, -128, -128, 127, -128, 22, 127, 51, -83, -44, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 9, 127, 127, 127, 127, 17, 127, 127, -128, -91, 127, -128, 127, -9, 127, 23, -128, 107, -128, 127, -24, 127, 28, -128, -128, -128, -60, -128, -128, -53, -128, 126, 47, 90, -66, -128, 127, -128, 127, -26, 36, 127, -128, -128, -28, -128, -1, -128, -128, -128, -43, -109, 127, -23, -128, 127, -128, -60, -128, 127, 66, 127, 127, 127, 127, -41, 127, -128, -128, -128, -30, 58, 59, 127, 127, -82, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 99, 127, 127, 127, 99, 127, 127, 7, 127, 127, 127, 127, 127, 109, -12, -128, -128, -128, 104, -128, 127, -128, 127, -105, -128, -128, -128, -109, 127, 127, 127, 127, -54, 127, -128, 6, -128, -128, -128, -128, -116, -23, 127, -128, 127, -128, 105, -128, -103, 76, -128, 95, -128, -128, -12, -128, 127, 127, 127, 127, 69, 127, -128, 127, 0, -9, 127, 64, 127, 18, 127, -128, 127, -116, 80, 127, -128, -89, 127, -128, -31, 127, 3, 127, -89, 127, -19, 127, 95, -128, 4, -128, -128, -128, -128, 88, 24, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, 90, 127, 127, 127, -80, 127, 75, -70, -128, -128, -128, -9, -3, 104, 119, -128, 72, -128, 71, 127, -128, 127, -128, 43, -128, -128, -106, -128, 38, -128, 127, -4, 127, -65, -37, -73, -128, -29, -76, -128, -128, -19, -128, 127, -128, 64, 98, -128, -128, -128, -128, -128, -128, -128, -74, 117, 30, -128, 124, -128, 87, -128, -128, -32, -128, -128, 127, -128, 127, -128, -128, 127, -128, 0, -128, -109, -128, -128, -128, -128, -128, -128, -127, -128, -128, -128, -128, 127, 127, 127, -3, 127, -128, 127, 127, 127, 127, 127, 112, 127, -128, -128, -128, -128, 127, 25, 127, 127, 127, -11, 13, -128, -128, -128, -128, 120, -48, -52, 6, -128, 78, -128, 127, -128, -128, -128, -128, -7, 127, 127, 127, -114, 51, 36, -128, 127, 127, 127, 127, 127, 40, -128, -120, -128, 123, 127, 127, 79, 27, -128, -128, -128, -128, 127, -19, 82, 127, -128, 127, -44, 127, 127, 127, 127, 127, -1, 127, -110, 127, 127, 127, 35, 127, -128, -28, -128, 100, 127, -81, 127, -102, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -75, 56, 127, 127, 127, 20, -128, -107, 127, 127, 127, 127, 127, 21, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -55, 127, -128, -128, -128, -128, 109, -21, 127, 127, 127, -128, -128, -128, -128, -128, -11, 3, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 64, 127, 96, 60, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 66, -128, -128, -75, -128, -24, -128, -128, -27, 70, -128, 60, -128, 127, 127, 127, 127, -36, -128, -126, -128, 127, -128, 127, -128, -128, -96, -128, 127, 113, 127, 127, -128, 127, 127, -37, 127, -128, -128, -128, -128, -111, -128, -128, -40, -128, -87, -128, 1, 76, 127, 48, 127, 127, 127, -128, 127, -128, 38, 79, 127, 127, 127, 127, -80, 60, -119, 127, -4, 127, 127, -128, -66, -128, -24, -128, 36, -128, 127, -128, -58, -30, -128, 108, -63, 107, 94, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 119, 127, 1, 127, -128, 127, -128, 127, -128, -128, -128, -105, -21, 127, 127, 127, 58, 127, -128, 111, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -42, -128, -128, 2, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 105, 127, -104, -22, -114, -128, -83, -128, -128, 127, -128, -128, 127, -128, -40, 36, -128, 68, -79, -128, 127, -128, -128, 46, -128, -128, -128, -61, -128, 127, 116, -69, 127, -128, 127, -94, -107, -128, 51, -128, -128, -128, -128, -128, -128, -128, -128, 3, -128, -29, 79, -128, 127, -62, 127, 127, 127, 127, 127, -19, -128, -128, -128, -128, -116, 127, 127, 127, 127, -94, -128, 127, 127, 43, 127, 127, 127, -128, -109, 127, -86, 127, 127, -82, -99, -128, -32, -128, 127, -63, -128, 0, 55, -128, 127, -128, 127, 127, 22, 127, 127, -128, 104, -128, 127, 127, -128, -112, -128, -128, 127, 127, 127, 127, -128, 127, -69, 30, -87, -128, 23, 10, -96, 127, 127, 127, 127, 124, 127, 93, -128, -128, -128, -128, 127, -128, 71, -128, 37, -45, -128, 72, -128, 64, -83, 41, 127, -128, 29, -128, 107, 127, 11, 127, 44, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -22, 127, 127, 127, 52, 127, -128, -128, -128, -128, -128, -128, -27, -128, 6, -128, -128, -128, -128, -87, -106, -27, 99, -71, 20, 127, -95, -128, 37, -111, 17, -108, 127, 127, 127, 127, -8, -65, -128, -128, -128, -6, -65, 127, -17, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -75, 127, -47, 31, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 89, 46, 60, -128, -61, -90, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 5, -128, -128, 127, 127, 127, -128, 127, 127, -56, 127, 30, -128, 48, -128, 113, -128, 12, 127, 120, 127, 127, 80, 27, -128, -128, -128, 3, 127, 127, 127, 127, 127, 127, 127, 46, 92, -128, -51, 127, -2, 127, 127, 127, -128, -128, -128, -128, -128, 127, -2, 127, 127, -128, -5, -128, -128, 111, -128, -43, -128, -128, -128, -128, -47, 7, 22, 127, 43, 127, 64, 64, 127, -128, 127, 127, -8, 127, 127, 92, 127, -128, -128, -24, -122, 127, 127, 127, -76, 127, -128, 127, -128, 127, -128, 127, -128, -27, -128, -114, -128, -128, -128, 1, 82, -14, 108, -128, -128, -128, 109, -128, -124, -65, -128, -128, -104, -128, -57, -128, -128, 127, -128, 127, 40, 127, -128, 72, -128, 126, -128, 127, -123, -86, -128, -128, -128, -93, -128, 23, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 63, -128, 127, -128, -128, -128, -17, -128, 23, -128, 127, -128, 127, 62, 127, -128, -128, -128, -128, -128, 127, 127, -32, -128, -128, -128, 47, 9, 127, 71, 127, -128, -53, -10, -40, -128, 100, 69, -128, -80, -128, -128, -128, -128, -91, 73, 127, 127, 127, 127, -128, 127, -68, 96, -92, 127, -128, 127, -128, -36, 127, 3, 111, -128, -128, -128, -128, -128, -128, 117, -128, 17, -128, 44, -128, 112, 52, -128, 127, -18, -128, 127, -128, 102, 12, -62, 127, -128, 127, -128, 127, -128, -81, -128, -128, 26, -128, 127, -77, 37, -128, -128, -128, 127, -128, 93, -128, 127, -13, -18, 127, -128, 127, -128, 29, -20, -85, -128, 127, -128, 127, -128, 127, -128, 127, -128, 70, 104, -61, 99, 127, 127, 73, 119, -39, 127, -104, 127, 127, 127, 127, -128, -128, -74, 18, 39, 127, 112, 17, 90, -128, 127, -128, 14, -128, -82, 127, 65, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 39, 62, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 76, -128, -128, -128, 58, -128, 94, 127, -128, 127, -128, -107, -128, -128, -9, -128, -128, -128, -128, -25, -128, -128, 127, -128, 127, -62, 127, -24, 127, -128, -128, -128, -128, -128, -128, 12, -128, -128, -128, -128, -128, -128, -128, 44, -128, 127, -43, 127, 127, 127, 127, -20, -46, -128, -128, -128, -128, -128, -128, -128, -71, -107, 127, 117, 127, 127, -128, -107, -128, 1, -128, 57, 123, 127, 127, 127, 127, 127, 97, -128, -120, -128, -128, 4, -58, 127, 87, 127, 127, 127, 127, 127, -1, -128, -26, -128, -128, 65, -128, 127, 127, 127, -32, 80, -128, 63, -128, -128, -128, -128, -128, 29, -128, -128, 32, -25, -128, 31, 30, -128, -128, -128, 110, 127, 127, 127, -128, -55, 18, -54, 87, -128, -128, -128, -128, -128, 127, -56, 127, 127, 127, 112, 127, -128, -128, -128, -128, 100, -128, 127, -128, 7, 0, -128, 20, -128, 112, -25, 95, -15, 127, -128, -69, -128, -38, -79, 127, 114, 127, 127, 127, 96, 127, -14, 127, -128, 127, -14, -62, 21, 127, -128, -128, 127, -49, 127, 127, 110, 127, 127, 127, 127, 127, 127, 127, 25, -57, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 37, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 89, -128, 127, -128, -80, 127, -128, -59, -43, 119, -128, 127, -20, 127, -54, -128, 10, -128, -128, -128, -128, 127, -128, 127, -89, 37, -128, -128, -128, 23, -128, -106, 51, -41, 127, -7, 127, -128, -43, -128, -128, 127, 127, 127, 127, 62, -128, -128, -128, 81, -128, -69, 127, 81, 127, 127, 127, 127, -12, 127, 10, 59, 127, 127, 127, 20, -128, -128, -128, 12, -128, 79, -128, -128, -128, -90, -128, 127, 15, 127, 54, -128, 119, -103, -128, 69, -128, -22, -128, 89, -128, 1, -128, 52, -128, -111, 127, -128, 127, -128, -104, -76, -128, 127, -128, 34, 127, -19, 127, 127, -128, -91, 27, -128, 127, -11, 127, 127, 127, -128, 127, -23, 12, 127, -91, 49, -128, 74, 127, 127, 127, -89, -42, -128, -128, 80, -128, 127, -128, -73, -128, -128, 41, 127, -128, 127, -128, 127, -128, -128, 127, 7, 127, 127, 127, -128, 127, -128, -128, 92, -128, -128, 1, -128, -37, -128, 127, 56, 127, -6, 127, -63, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 83, 127, -128, 127, -128, -128, -128, -128, 127, -111, 127, 127, 127, 127, 60, -128, -8, -128, -88, -128, 14, 127, -128, 127, 127, 127, 80, 127, -128, 0, -128, 127, 127, 127, 127, 127, 87, -128, 127, -128, 103, 127, 127, 127, -128, 127, -3, -49, -27, 39, -128, -128, -128, 91, -128, 127, -57, 127, -128, -128, 127, -128, 57, -128, -128, -128, -103, 127, 127, 127, 127, -128, 72, -128, 127, -85, 127, 127, 79, 127, 127, 127, 0, -110, -128, -128, -128, -128, -128, -43, -128, 25, -99, -128, 7, -128, 127, 127, 117, 127, 127, 39, 127, -128, 127, -112, -128, -17, -128, -128, -128, -128, 127, 127, 127, 127, -9, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -32, -128, -83, 75, -78, 127, 127, 127, 127, 127, 127, -2, 40, -128, 127, -58, 127, 127, 127, 127, 127, 124, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -108, -128, 127, -68, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -80, 17, -18, -128, 127, 127, 127, 127, -128, -30, -36, -128, 127, 127, 107, 124, -128, 127, -120, 127, 106, 127, 57, 103, 127, 127, 127, 65, -128, -113, -128, 127, -128, 15, -34, 127, -25, 127, 82, 127, 127, -128, 127, 127, -80, 127, 127, -128, 79, -128, -128, 98, -128, 127, 127, 127, 127, 127, 88, 57, -128, 127, -57, -128, -37, -128, -128, -128, -128, -100, -128, -62, -128, -27, -128, -128, 75, -51, -88, -18, 58, -46, 44, 60, 122, 127, 127, 15, 127, 127, 127, 127, 127, 127, 60, 127, -59, 25, -128, 28, -128, 13, -128, -128, 127, -128, 127, 126, 127, -2, 71, -122, -128, -128, -93, 127, 127, 127, 127, 127, 127, 127, 20, -113, -128, -128, -128, 36, 54, 127, 127, 127, 105, 127, -2, 127, -128, -128, -128, -128, -119, -83, -128, 114, 2, 127, 127, 127, -128, -128, -128, -128, -28, 127, 32, 127, 96, -128, 127, -128, 127, -45, 127, 127, 15, -115, 127, 49, 127, -69, 127, 23, -10, 82, -11, 127, -128, 127, -128, 82, -128, -128, -128, -128, -47, 4, 53, 127, -128, 44, 94, -128, 89, 37, 127, -128, 127, -128, 127, -14, 127, 127, 127, 88, 88, -8, 5, -31, -128, -128, 18, -128, 43, 127, 127, 127, -63, 49, 25, -128, 2, -128, -128, -128, -2, -128, -128, 127, 20, 117, 41, 127, 59, 29, 61, -73, 127, -23, -128, 127, -128, 59, 58, 126, 127, 127, 127, 127, -68, 127, -128, 68, -128, -116, 127, 27, 127, 127, -128, 127, -128, 6, -128, 127, -83, 123, -128, 127, -128, 127, 127, 127, 127, 127, 87, 127, 9, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 70, 127, 127, 127, 127, -93, -128, -128, -65, -8, 127, 127, 127, -128, 127, -128, 127, 98, 127, 127, -13, 127, 46, 127, 127, 127, 112, 127, -128, 11, -128, 127, -128, 127, -128, 43, -58, -128, 127, 55, 127, -128, -125, -128, -128, -128, -128, 127, 52, -128, 47, -128, -128, -77, 11, 127, 127, 127, 127, 127, 29, -56, -128, -128, -128, -128, -71, 127, -15, 127, 127, 127, 0, -128, 127, -38, -49, 127, 127, 127, 127, -128, 127, -128, 127, 127, -26, 127, -92, 127, 80, 127, 127, 127, 127, 127, -119, -128, 121, -128, 127, -128, 127, -128, -55, 96, 127, 127, -96, 127, -58, 127, 127, 44, 117, -44, -128, -128, -128, 72, -128, 127, -128, 127, -128, 127, -128, -128, -116, -128, -128, 127, 127, 127, 127, 127, 92, -128, 29, -128, 127, -128, -40, 127, 37, 127, -11, 54, -128, -128, -128, -128, -126, -21, -23, -83, -128, -128, -128, 127, -128, -128, -106, -128, 127, -128, 127, 127, 127, 52, -128, -117, -128, 127, 62, 127, 127, 127, 127, 127, -126, -128, -128, -128, -128, 46, 127, -128, 127, -128, 58, -128, -128, -48, -128, -128, 43, -128, -74, -128, 127, -128, 127, -128, 127, 54, -94, 127, -128, 127, -128, 127, -128, 127, 10, 127, 127, 127, 121, -48, -128, -128, -128, 127, 122, -2, 127, 12, 127, -48, -128, -128, -128, -128, 127, 102, 127, 127, -128, 62, -108, -56, -71, 127, 127, -128, 127, -128, 127, -128, 127, 112, -128, -105, -128, -128, -128, -128, -128, -72, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -109, -128, -9, -128, 127, 127, -100, 127, -128, -41, -128, 127, 127, 127, 127, -62, -128, 127, 125, 127, 127, 121, -125, 72, -70, -73, 127, -128, -128, -128, -128, -128, -6, 127, 127, 127, 71, 127, 35, 127, 127, 95, 127, -45, -128, -128, -128, -128, 71, 31, 127, 127, 127, 127, -128, -128, -128, -128, 100, -128, 127, -128, 127, -77, 127, 127, 127, 127, 127, -19, 127, -14, 127, -20, 127, 127, 127, -26, 127, 66, 127, 13, -28, -128, -29, -128, 66, -128, -107, -128, -128, -123, -128, 127, 77, 127, 127, 25, 127, -128, -10, -128, -115, -128, -85, -128, 127, -58, 127, 127, 127, 127, 127, 127, -128, -24, -128, -128, 127, -128, 127, 26, 127, 127, -128, 127, -128, -128, -128, -128, -20, -128, -128, -128, 127, -41, 127, -128, 2, -128, -128, 83, 127, 127, 127, -55, -128, 127, -128, 127, -128, 127, 77, -128, 85, -128, -128, -128, -128, 78, 71, -55, 127, -128, -114, -128, -128, 0, -128, 127, 47, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, 122, -128, -128, -128, -128, 127, 7, -31, 127, 127, -6, 127, -128, 127, -128, 120, -128, -120, -128, 14, -55, 91, 127, 31, 127, 37, 13, 127, -23, 127, 127, -128, 127, -128, 87, 127, -128, 127, -128, -64, 127, -78, 127, -51, 19, -128, -128, -128, -128, -87, 1, 127, 75, 127, 127, 127, 127, 127, 127, 22, 127, -128, -128, -108, -128, 19, 127, -128, -35, -128, -128, -46, -18, 127, -128, 106, -128, -128, 68, 6, 127, 127, 127, -70, -45, 112, -128, -128, 94, -100, 127, -128, -95, 127, -128, 127, 41, 100, 127, -128, 40, 6, -128, 19, 65, 40, 127, 85, -4, 127, -128, -128, -128, -128, -128, -128, 123, 58, 127, -128, 127, -128, -127, 116, -88, 127, -128, -72, -128, 127, 78, 127, 127, 127, 64, -128, -128, 46, -128, 127, -128, 127, 127, 127, 127, -128, -28, -128, 127, -69, 127, -68, 127, -128, 127, -128, 95, -128, 127, 127, 74, 81, -128, -128, -128, -128, 32, -128, 36, -128, 1, 127, 63, 127, -39, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -58, 127, 127, 127, 127, 80, -128, -15, -128, 25, -128, 127, 127, 55, 127, 127, -128, 127, -128, -128, -128, -128, -82, 30, -128, -128, -13, -47, 11, -87, -128, -128, -128, -82, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -55, 127, 127, 127, 127, 127, 127, 127, -40, 127, -128, 127, 109, 127, 127, 117, 127, 127, -65, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -19, -128, -80, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -108, -128, -128, -128, 127, 29, 127, 127, 127, -128, -128, -128, -85, 127, -128, -21, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -55, 127, 127, 127, 127, 127, 127, 90, -12, -128, -109, 127, 127, 127, 127, -128, -128, -48, -128, 127, 48, 127, -27, 42, -12, 68, -128, 127, -128, -128, 127, -76, -128, -15, -47, 127, -62, 127, 127, 127, 127, 127, 127, 40, 90, -128, -128, -128, 127, 21, -26, -75, -128, -128, -128, 127, 127, 127, 127, -128, 127, -122, 127, 127, 127, 127, 66, 127, -128, 127, 5, 127, 127, 127, -54, 127, -128, 127, -124, -128, 69, -128, -128, -128, -128, 4, -128, 127, 97, 73, 126, -128, -41, 127, -128, 127, -128, 127, -73, -128, 127, -128, 127, -74, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, 107, 127, 127, 127, 127, 127, 127, 127, 127, -128, -127, 12, -128, -2, -128, -128, 127, -128, 127, 127, -94, 81, -128, 127, 127, 127, 127, -128, -128, -128, -63, 37, 7, -114, -78, -128, -31, -99, -89, -128, -128, -128, -128, -43, -128, -10, -128, 127, -128, 127, -128, 77, -128, -128, -88, -58, 127, 127, 127, 127, 127, 127, -26, 127, -98, 127, 87, -122, -34, -128, -126, -128, 127, -128, 127, 127, -80, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -27, 0, 127, 127, 127, 127, 127, 127, 127, 127, 127, 23, -48, -123, -128, -128, -128, -128, -57, -128, 127, -128, 44, -128, -128, -128, -58, -128, 127, -99, 127, 2, -128, 122, -128, 45, -128, 127, -128, -21, -128, -128, -128, -9, 127, 127, 83, -90, -128, -128, 58, 81, -128, -128, -128, -128, -128, -128, 71, -128, 127, -128, 77, -128, 127, -128, 127, -128, -128, 127, -128, 121, -128, -128, 86, -20, -128, -9, -53, -128, -128, -128, 127, 127, -3, 109, -58, -128, 127, -96, -22, 127, 120, 127, 127, 127, 127, 71, 127, -128, 127, -128, 127, 93, -128, 127, -128, 20, -128, 127, -94, -91, 127, -7, 94, 127, -117, 127, -128, -128, -128, -128, 105, -128, 24, -128, -82, -17, 56, -69, 127, -128, 127, -128, 127, -117, -128, -111, -128, -128, -128, -128, -128, 64, -12, -74, 127, -59, -53, 55, 127, -89, 127, 93, 127, 78, -128, -128, -126, -128, -39, -128, -128, 127, -128, 127, 127, 127, 110, -128, 111, -128, -128, -128, -128, -12, -128, -57, 127, 127, 127, -128, 127, -128, -128, 89, -128, 9, -43, -128, -128, 127, 127, 127, 75, 127, 9, 127, 127, 91, 127, 127, 96, 127, 127, 3, 70, -128, -128, -128, -128, -128, -127, -128, -128, -94, -13, -128, 30, -128, 72, -128, -128, -83, -128, -128, -23, 32, 127, 18, -128, -45, -128, -128, -128, -128, 85, 127, 115, 127, 127, 127, -115, 127, 10, 127, -128, 46, -128, -128, -128, -128, -128, -128, -128, 127, -58, 127, -128, 127, -21, 127, 119, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -34, -128, 127, -128, 127, -128, 127, -6, -9, 127, -128, 127, -39, -38, -128, 127, -128, 127, -128, -3, 127, 11, -128, 54, -79, 126, 21, -66, 127, -128, 24, -104, 127, 127, 24, 127, 108, 127, 103, -128, 127, -128, 127, -128, -113, -128, -128, -128, -128, -128, 95, -20, 29, 127, -128, 127, -96, 127, 8, 127, 127, -29, -31, -51, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 23, -57, -31, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 19, 127, -1, -128, -28, -128, -128, 108, 66, -2, 127, -128, 127, 127, -128, 127, 7, 127, 127, 127, 127, 127, 68, 127, 127, 127, 127, -128, -116, -128, -128, -128, 127, 41, -123, 9, -128, -41, -128, -26, -128, -106, -128, -128, -128, -128, -128, -96, -128, 76, 127, 127, 70, 85, 127, -128, 127, -128, 127, -128, -128, -55, 58, 127, 127, 127, 127, 127, 25, 58, -110, -128, 127, -128, 127, -128, -10, -57, -128, -128, -13, -128, 49, -21, -74, -128, -128, -83, -128, 127, -128, -52, -128, -128, -128, -128, -128, -128, -62, 114, 6, 127, 127, 127, 28, 60, 117, 91, 127, 127, 127, 87, -108, 127, -128, 127, -51, 127, -128, -61, -128, -128, -128, 91, 127, 98, 93, -128, 24, -128, -128, -128, -128, -9, 127, 127, 127, 127, 127, 127, 127, -48, -128, -128, -128, 114, 127, 127, 127, -128, 89, -90, -128, 127, -128, 127, -128, -128, 127, -128, 127, -85, 127, -128, 43, -128, 127, 1, 127, -128, -105, -128, 125, -89, 127, 127, -128, 127, -91, 127, -128, 127, -128, 86, -128, 127, -128, 127, -128, 126, -65, -128, -128, -128, -128, 127, -76, 127, 18, 127, -108, -128, -128, 127, -128, -2, -37, -128, 72, -128, 71, -128, -108, -128, -128, 9, 127, 127, 127, -27, -128, -128, -128, -128, -128, -128, -128, -15, 127, -1, 127, -128, 127, -95, -128, -31, -128, 127, -9, 127, -48, -128, -128, -128, 38, -128, 68, -128, 127, -128, 127, 127, 127, 127, 127, 42, -128, -128, -128, -128, 127, 127, 127, -41, 127, 108, 127, -48, 127, 127, -128, 127, -128, 127, -89, 30, -128, 127, -128, 127, -128, -13, -128, -59, -128, 96, -64, 127, 35, -112, 127, -36, 127, 127, 127, 127, -60, 127, -106, -128, -128, -128, 7, 127, 127, 127, 127, 120, 127, -128, 127, -128, -128, 105, -128, 127, -128, 97, -49, -128, 127, -128, -128, 127, -128, -6, -104, -128, -128, -128, 127, 127, 127, 127, 117, 127, 127, 127, -128, -128, -128, -128, 127, 85, 127, 122, -128, 114, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 121, -128, 127, 69, 127, 127, -128, 11, -128, 127, -128, 127, 127, 127, 127, -128, -58, -128, 127, 115, -128, 127, -128, 127, -128, 127, 127, 127, 52, 127, 55, 127, 127, -128, -62, -128, -128, -128, -128, -54, -57, 127, 0, 127, 127, 127, 127, 127, 127, 127, 58, -128, -128, 76, -34, 127, -128, 26, -128, -96, -128, -56, 127, -58, -13, -65, -128, 127, -65, -128, -7, -128, -128, -128, -22, -128, 127, -128, 127, -128, 127, 125, 21, 127, -128, 127, -128, 127, -128, -128, -38, -128 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
