-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            -36, -78, 119, -95, -93, -11, -10, -101, 56, 56, 86, 83, -91, -54     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( 81, 12, 0, 48, 11, -41, 64, 39, 1, -76, -40, -124, 124, 45, -109, -121, 28, 94, -78, -50, 13, 43, -117, 14, -26, 67, -103, 32, 124, -30, -110, -97, -28, 109, -67, 35, -52, -24, 5, -13, 61, 105, -19, -125, -47, -72, 14, 50, 127, -1, -104, -37, -70, -109, -16, -19, -56, -98, -127, 92, -23, 42, 45, 25, 9, 2, 59, -104, -80, -100, 106, -7, -47, 109, 119, 19, 41, 125, 118, -104, -68, 48, -98, 10, -24, -13, -69, -4, 97, 76, -1, -23, -29, 22, -3, 5, 89, 37, 127, 86, -51, 89, -11, 91, -84, 87, 57, -81, 106, -35, 82, -63, 56, -83, -74, -50, 121, -32, -112, -105, 118, 111, -93, -14, 41, -50, -114, 115, 95, -10, -46, 95, -125, -94, -28, 16, -93, 124, -17, 11, -21, 83, 105, 71, -11, 13, -65, 28, -20, 47, -34, -75, -56, -75, 127, 116, 55, 38, 127, -33, 3, 126, 50, 81, -87, 113, 106, 78, -48, -77, 51, 33, 90, -104, -49, 88, -109, 24, 11, 40, -108, 40, 112, 68, -81, -111, -87, 43, 59, 108, -80, -13, 82, -94, -22, 11, -78, 67, 125, -40, -118, 28, -52, 106, -84, -60, -86, -107, -95, 69, -93, -22, -96, 24, -36, -57, 46, 32, 113, -60, 63, -52, 18, -94, 3, -2, 12, 122, -41, -35, 8, -59, 126, -68, -4, 63, -11, -50, -17, 118, 68, 33, -3, -92, 72, 61, -27, 34, 125, -14, -79, 32, -78, 10, 75, -3, 38, -70, 79, 56, 109, 25, -64, 18, -2, 16, -68, 112, 86, -115, 60, -80, -103, -92, -28, -95, -87, -39, -115, 81, -35, -107, 110, -40, -114, 105, -52, 93, -80, 112, -4, 43, 87, -121, -119, 86, 1, 6, 25, -4, -65, 3, 114, 63, -12, -54, -124, 32, -111, -98, 17, -47, -112, -1, 100, -8, -101, 15, 24, -116, 122, -2, -122, 35, -69, -63, -33, -95, 4, 84, 81, 126, 5, 67, -23, 66, 1, -92, 31, -126, 48, -116, -127, 3, 121, 76, -103, 0, -87, -35, -105, -86, -38, -22, 78, 30, 8, 92, 42, 46, -103, 34, -30, -2, 76, 110, -68, -43, -126, 33, -67, -33, 68, 47, -126, -41, -20, 100, -51, -120, -5, 58, 66, 42, 115, 86, 58, -89, -112, 42, -36, 72, 94, 109, -106, -28, -70, 115, 38, -29, -8, 37, -11, 52, -36, -59, -16, -5, -25, 3, 13, -35, -57, -73, -65, -66, -32, -47, -82, -80, -61, 16, -121, 50, 124, -91, -50, -106, -43, 57, 96, 30, -20, -82, 53, 22, 93, 125, -25, -8, 124, -123, 29, -24, -10, 81, -70, -101, -40, 35, 70, -119, -98, 31, -51, -6, -48, 75, 31, 91, -121, 19, -51, 75, -59, -67, -15, -57, -88, 125, 20, 29, 11, 105, 126, -111, -20, -81, 41, -128, 19, 97, 71, -37, 41, -47, -2, -120, -116, -38, 108, -70, 24, -113, -55, 60, 42, -93, -62, -44, -8, 48, -7, -9, 75, 30, 95, -121, 41, -125, 2, -51, 61, 114, -4, 55, -35, 16, -30, -63, 37, 105, -126, 32, -63, 91, 112, 69, 105, 77, -15, -40, -39, 15, -127, 117, 64, 111, 14, 77, 95, 81, -50, -101, -128, -86, -63, 77, -79, -55, -4, -82, 100, 51, -47, -119, 64, 8, 57, -32, 22, -57, -100, 26, 103, 43, 44, -28, 51, 39, -54, -73, 1, 63, -117, -66, -45, -63, 127, -75, -70, -43, 71, 102, -57, -62, 124, 39, -57, 18, -19, -14, -83, 68, 112, -117, -80, -122, 37, 98, 32, -7, 69, -16, 28, 20, 79, 88, -94, -27, 19, 97, -4, -38, 11, 0, 61, -8, -48, -48, 78, 68, -69, 92, -106, 3, 122, 74, 117, 62, -63, -20, -3, -85, 57, 0, 46, -109, 36, 13, 109, 8, -20, 60, -50, 24, -26, -72, -72, 105, 83, -69, -109, -90, 114, 25, -11, 34, 76, -20, 91, -47, 98, 61, 53, 76, 72, -43, 126, 38, -60, -47, 3, 123, 45, -22, 33, -99, 86, -77, 86, 40, -50, -45, -65, 19, 96, -87, -107, -10, -127, 97, 41, -118, 72, 45, -60, 27, 124, -91, -58, -79, 42, -106, -120, 56, -105, 126, 105, 87, 52, -9, -71, -9, 108, -19, 12, -70, 26, 96, 44, -28, 100, 61, 24, 72, -78, 65, 125, -117, -57, 102, 74, 45, -67, 9, 71, -76, -64, 27, 64, 118, 80, 88, -75, 12, 107, 40, -36, -128, 18, 23, -94, 71, -107, 94, -122, 6, -96, -79, -74, -113, -1, -106, -125, -103, -24, -16, 122, 63, 123, -13, 44, -67, 36, -58, 97, 61, 41, 20, 36, -36, -73, 31, 125, -5, 38, 93, 61, -92, -122, 65, -70, 37, 95, -48, -51, 107, 111, -35, -21, 127, 110, 97, -126, -42, -54, -92, 43, -121, 117, -97, 113, 44, 32, 20, -72, -75, -116, 127, -46, -73, 16, -56, 4, 45, -65, 44, -118, -102, 70, -28, 35, -62, -116, 125, -86, 99, -36, -15, 120, 23, -56, -72, -45, 24, -119, 50, 47, 88, -62, 91, 114, -70, -19, 17, 57, -125, 6, -115, 84, -45, -125, -63, 32, -99, -13, 60, -3, 25, -19, -107, -109, -113, 45, 3, 20, -26, 33, 44, 47, -57, 114, -57, -49, -8, 47, 35, 112, -29, 85, -10, -21, 18, -93, -33, 58, 81, -111, -74, 85, 118, 4, -18, 13, 36, 45, -7, 54, -99, 92, 27, -92, -66, -91, -56, -56, -85, 29, 75, 56, 113, 89, -77, 92, -16, -97, 26, -27, 41, 70, -38, 90, 47, -51, 41, 5, 39, -126, 114, 11, 65, 11, -117, -4, 116, 83, 16, -67, -48, -43, 125, 52, -24, 94, -4, -77, -110, -17, 37, 49, 86, -104, 86, 82, -74, -86, 56, 119, 34, -89, -16, -8, -70, -25, -27, 99, -103, 62, -9, -36, 116, -54, 70, -90, 90, 103, -66, -126, 127, -28, -93, 6, -113, -15, -3, 17, 127, -2, 90, 102, 36, -123, -94, 100, -105, 4, -40, 16, 81, -98, 33, 0, -98, 22, 97, -106, 48, 124, -105, 94, 39, -75, 74, 101, -80, -128, 11, -92, 37, 54, -26, 25, -56, -101, 41, 35, -73, -22, 14, 36, 23, 20, 99, 36, 107, -23, 122, 66, 29, -43, 74, -67, -61, 103, 61, 79, -118, -101, 3, 62, 37, -30, 43, 87, 29, -67, -105, -7, 44, 76, 33, -46, -96, 112, 75, 14, 97, 34, 126, 98, -117, 43, -106, -106, -45, 29, 76, -120, -27, 33, 24, -23, 28, 82, -47, -9, -35, 120, -24, 58, -3, -109, 40, 112, -115, -23, -8, 40, -87, -110, 23, 101, 11, 126, 115, 126, -112, 32, 43, 40, 111, 41, -85, -27, -122, -54, -33, 12, -22, 73, -77, 118, -83, 115, 42, -116, -83, 67, 57, 52, 78, -28, -12, 42, -22, -70, 11, -79, -24, -61, -74, 44, 49, 127, 91, -18, -69, 100, -62, 11, -61, -125, -63, -74, 87, -44, 71, 3, 106, 95, -105, 58, -12, -30, 120, 0, 48, -79, 111, -116, -8, -121, -62, 52, 68, 58, -48, -67, -82, 24, 49, 1, 84, 20, 74, 120, -79, -104, 33, -107, 46, -93, 95, 17, -20, -92, 70, -30, 8, 20, 98, -26, 78, 80, -119, 100, -41, 57, -75, 58, 110, -92, -102, -71, 69, -13, -9, 24, 94, -118, 97, 56, -12, -122, -11, -15, -114, -106, -93, 80, -42, -14, -110, 89, -57, -81, -87, 120, 116, 86, 98, 121, -33, 34, -13, -53, -34, -60, 68, 95, -37, -71, -61, -35, 16, -61, -21, -98, -28, 107, -46, -113, -102, 23, -49, 84, 93, -91, 58, -32, 98, 126, -68, 23, 86, 84, -103, 22, 62, 16, -23, 12, -52, -45, -42, 24, 61, -90, -49, -21, -8, 23, 14, 53, 92, -58, -30, -23, -2, 83, -3, 121, 45, 14, 89, -92, -126, -6, -116, 18, 37, -2, -50, -63, 13, -127, 87, 2, -62, 11, 49, 69, -19, -1, 93, -117, 113, -118, 44, 91, -48, -68, 81, -31, 46, -107, 110, -5, -62, 113, 17, 1, -85, 90, -116, -48, 98, -86, -43, -2, -2, -55, 118, -13, 87, -119, 46, 107, 82, -31, -51, -89, -123, -30, -67, -121, -47, -50, -93, 93, -60, 74, -59, 3, 27, -100, -2, 70, 4, -120, 115, -17, 117, -122, -116, 23, 66, 36, 127, -127, 13, 45, -99, -37, 55, 86, -120, -110, 6, 54, 47, -93, 72, 120, -94, 121, -97, 7, -5, 85, -10, 79, 15, 35, 83, -67, 46, 23, 96, 98, 63, 49, 22, 33, -36, 45, -12, 70, 60, 98, 20, -101, -16, -29, -22, 112, 63, 84, -122, -88, 61, 72, 6, -36, 125, -57, 79, -98, 57, -90, -37, -18, 75, -46, -60, 76, 35, 76, 27, -21, 95, -108, 1, -23, -47, -121, -108, 33, -63, -77, -76, 103, 67, 17, -44, -21, 60, 10, 94, -104, -54, -45, 57, 107, -9, 22, 90, -35, 117, 45, 1, 115, -41, 55, 34, 7, 78, 98, 120, -43, 90, -23, 56, -12, 17, -39, -43, -73, -56, -101, -73, 1, 84, 110, -104, -93, -31, 73, 59, -98, -40, -16, 37, 18, 71, 30, 105, -82, 7, -33, 33, 29, 0, 13, -92, -80, 94, -87, -28, 37, -81, 13, 66, -70, -92, 78, -53, -124, 62, 106, -112, -17, 96, -58, -24, 32, 38, 87, -116, -28, 42, -119, 107, -50, 21, 13, 13, -44, -56, -86, -69, 74, -65, 6, -71, 112, -110, 14, -114, -58, -28, 37, 23, 107, 9, -51, 42, -115, 10, 126, -3, -46, 108, -20, -112, 11, -97, 44, -59, 112, 76, 20, -31, 68, -109, -119, 31, 67, 28, 11, -99, -57, 103, -26, -60, -81, -40, 62, -32, -12, 125, -1, 31, 6, -76, 124, 91, 35, 22, -44, -73, -87, -123, 75, -4, 36, 93, 59, -118, 80, -101, 104, 55, -71, -65, 100, 125, 38, -9, -42, -82, 114, -124, 48, -32, -112, -115, 107, -26, 80, -44, -71, -99, -12, -65, -25, 45, -4, 89, -121, 100, -25, -29, 57, -55, -88, 74, 27, 31, 100, 9, -98, -87, -111, 25, 48, 104, -13, 125, -96, 55, 106, 123, 115, -79, 121, -73, -21, -14, -34, -93, -12, 89, -50, -15, -87, 17, 105, 104, -55, 51, 121, -112, 72, -4, -8, -90, 9, 99, -120, -21, 31, 74, -84, 96, 49, 22, -102, 60, -59, 79, -48, -104, -81, 5, 65, 36, -19, -91, -112, -18, -96, -33, 96, -95, 4, -105, 49, 10, 12, -17, 93, 84, 104, 95, -82, -18, 4, 95, 109, 108, 20, 4, 3, -27, 108, 88, -51, -108, 97, -46, -106, -19, -68, -57, 5, -122, -56, 38, -118, 48, 5, -92, 4, 115, 127, -115, 98, -11, 70, 4, 111, -8, 12, -87, -46, -9, -61, -3, -93, 52, -124, -88, 9, 5, -40, -65, 115, 3, -28, 17, 9, 124, -53, -29, 113, -49, 41, -61, 14, 106, -20, 80, -85, -31, 9, 78, -119, -42, 7, -49, 122, 65, 47, -9, -11, -97, 79, -72, -82, 45, -14, -114, 53, -81, 113, -66, -124, -94, -122, 38, 49, 98, -74, 121, -74, -30, -113, 75, 114, 90, 19, -17, -6, -20, -127, 67, 24, 68, -78, 106, -120, -57, 64, 95, -117, 57, 104, 33, -58, -118, -28, -37, 14, 55, -103, -85, -123, 113, 4, 12, -128, -34, -128, 4, 102, 23, 114, 37, 64, -37, 62, 82, 94, 88, 124, -107, -5, -82, 27, -52, 0, -42, -111, -113, 126, -63, 34, 53, -11, 75, 123, 67, -36, 114, -85, 111, 89, 111, -36, 53, -36, -8, -36, -70, -46, -79, -83, 54, -62, -40, -14, -46, -63, 17, 107, 122, 109, -30, -41, 111, 50, -70, 18, 127, -102, 25, 36, -1, -67, 33, 97, -122, -8, 87, 5, 9, -14, -108, -66, 25, 27, 105, 122, -25, 86, -100, 58, -114, -93, -127, 91, -24, -37, -9, -23, 119, -20, 62, 105, 33, -114, 51, 9, -27, -79, 80, -45, 68, 48, -120, -67, -15, -65, 62, 7, -48, 71, 28, 14, 124, 93, 102, -34, 51, -43, -54, 57, -73, 55, 48, 27, 115, 65, 48, 53, 60, 34, -73, -21, -6, 45, -125, 94, 120, -27, 6, 7, -30, -91, -78, -56, -6, -112, 111, -110, 34, -53, 108, 107, -54, -93, -45, -111, -122, 75, 73, -86, -106, 17, -51, 73, 31, -66, 38, 41, -33, -67, -111, 81, -28, 92, 53, -12, -125, -15, 56, 110, -86, -81, 112, -47, 78, 36, -106, 115, 108, 94, 99, -61, 111, 99, -92, -65, 47, 27, 15, -114, 49, -99, -30, 28, 108, -125, 86, 68, 52, -27, -43, 3, 85, 68, -26, -44, -47, -88, -43, 103, -17, -118, 2, -123, 7, 32, 91, -90, 3, 40, -72, -111, -119, -99, -125, -83, 33, 43, -121, 41, -49, -64, -69, -109, -77, 19, 48, 23, -4, -125, -125, -50, -88, -85, 66, -112, -90, 117, -82, 17, -90, -16, -96, 40, 53, 82, 18, 33, -22, 75, -64, -124, -93, 74, -119, 80, -40, 8, 44, -36, -8, -87, -125, 73, 12, -9, -32, -25, 117, -17, 91, -71, -125, 107, -121, 77, 121, -56, -51, -88, 22, 43, 87, -1, 52, -111, -40, -73, 120, -19, -70, -72, -78, -55, -83, 7, -11, 111, 16, -114, -89, 63, 34, -56, 64, -4, 66, -43, -53, -110, -34, 75, -73, 104, -72, 111, -80, 111, -111, 105, -7, 4, -38, 42, -39, -5, -44, -19, -7, 114, 36, 10, 87, -99, -117, -61, 20, -50, -46, -51, -35, 117, -119, -53, 113, -22, -43, -89, -42, 47, -7, 113, 34, 5, -30, -6, -9, 18, -85, 50, 103, 1, -42, 19, -117, -58, 105, 63, 30, -117, -90, -21, -72, 44, 10, -68, 9, 63, 9, -6, 110, -8, -6, -51, -112, 86, -94, -92, 23, -29, 33, 125, -55, 43, -69, 87, 122, 18, -113, 114, 119, -18, -73, 107, -109, 83, 57, 25, 63, 98, -111, 52, 77, -122, -55, -19, 111, 15, 69, 92, 85, -123, 5, -65, -63, 108, -45, 22, 109, 97, 93, 66, -32, -73, 114, 97, 54, 15, 51, 15, -39, 38, -102, 5, -106, 72, -78, -74, 34, -33, 120, 101, 51, -58, -40, -23, 53, 110, -86, 101, 21, -23, -51, -101, 85, 41, -77, -71, 89, -59, 83, 90, -45, -66, 119, 121, -64, 32, -52, -32, -114, -111, 73, -1, -14, 106, -115, 100, -83, -111, 113, -30, -69, 4, -76, 106, 102, -76, -82, 112, -34, -20, 113, 31, 50, 41, 102, 100, -48, -86, 125, 46, -53, -51, 92, 21, -120, -29, -128, 55, -79, 48, 42, -81, 37, 2, 80, -106, -59, -24, -119, 28, -78, -12, -78, 126, -11, -45, 87, 8, -88, -8, -15, -70, 117, -109, 23, -80, 69, 19, 35, 50, -54, 105, -79, -93, 71, -16, -102, 93, -112, 59, -83, -37, 71, 77, 1, -41, -36, 111, 75, -105, -111, -97, 127, 102, -54, 62, -87, 10, 30, 29, -57, -29, 55, 21, -70, -104, 0, -90, 8, 80, 123, -5, 20, -128, -84, -46, -47, 124, 78, -7, -83, -11, -15, -15, -10, -4, 47, -118, -36, 7, 1, -30, 47, 35, -120, 107, 61, -63, -25, -29, -47, 103, -6, 102, 26, 93, 59, 60, 64, -18, 103, 0, 14, -68, -72, -12, -22, -124, -34, -45, 84, -96, 115, -54, 17, -123, -128, -13, 99, -39, 40, -60, -97, -44, 81, 109, -48, -117, -21, -14, -46, 60, -51, 96, 104, -11, -49, -90, 46, 64, -120, 10, -34, -73, -100, -54, 55, -19, -17, -102, -75, -58, -21, -63, 114, -18, 79, -65, 116, -49, -13, -94, 56, 23, 99, -109, -92, 95, 16, 49, 96, 38, 52, 49, -17, -31, -41, 65, -26, -49, -28, 21, 54, -45, 120, 72, 98, 44, -97, 108, 19, 33, 13, 82, -95, 109, 126, -83, -122, 117, -8, -63, 33, 31, -98, 11, -122, 93, 76, -49, -11, -61, 105, -44, -99, -38, 122, 81, -1, -90, 111, -43, -14, -121, -85, -62, 24, -55, -80, -46, -73, -1, -89, -75, -29, -81, 47, -128, 81, 76, -88, -64, -52, -92, -16, -128, 15, 49, -113, 83, 24, 102, 24, 39, -12, 43, 94, 74, -38, 116, -32, -42, -66, -10, 94, -86, -66, -102, -6, 118, 59, -106, -85, -102, -14, 53, -18, 75, 118, -21, -103, 46, -116, -19, 22, -52, -53, 56, 104, -62, 67, -32, 88, -30, 111, -15, 10, 0, -62, 122, 112, -96, -92, -84, 20, -30, 124, -7, -41, 103, 110, 116, 12, -5, 76, 34, -19, -125, -112, -86, -42, -90, -25, -35, 32, -44, -34, 91, 9, 106, 84, 124, -55, -126, 96, -76, -110, 101, 10, 124, -107, -54, -74, -35, 110, 98, -25, 75, 73, 86, 120, -102, -10, 123, -48, 102, 93, 35, 110, -63, -77, -61, 83, -96, 82, -13, 37, -107, 29, -79, -26, -77, 68, 28, 25, -87, 127, 62, -119, -40, 67, -15, 80, 1, 75, -2, -29, 62, -69, 85, -97, -16, -67, 93, -53, 83, 38, -111, -73, 72, 99, 114, -75, -10, 106, 74, 108, 66, -11, -2, -42, 26, -95, -1, -36, -45, 28, 48, -77, 103, 78, -103, -82, 89, 82, 38, 5, -96, 44, 117, 43, 117, 79, -105, -80, -2, -44, 106, 126, 60, -4, -84, 1, 45, -44, -85, 55, -108, -28, -11, 59, -5, 49, 20, -31, -120, 64, -4, -15, -58, -77, -23, -79, 83, 21, -63, 17, -41, -87, 87, -62, -6, 17, 62, 121, -48, 77, -112, 61, -17, 71, -83, -3, 109, -65, 53, 57, 59, -62, -113, -28, 21, -26, -69, -118, 114, -52, 33, -128, 26, -89, 87, 66, 31, 30, 32, -99, -85, -57, 81, -126, 30, -13, 99, 83, -120, 20, 105, -25, -109, -108, 64, -58, -86, -107, 67, -72, -17, -31, -79, -24, 4, -11, -50, 25, 65, 17, -46, 87, 62, 17, 68, 87, -19, -58, -35, 32, 25, -115, 15, -116, 41, -60, 9, -97, -18, -81, 58, -104, -24, 90, 68, -26, 9, -17, -29, 84, -109, -85, -15, -40, 33, -29, -44, 94, -72, -103, 23, -99, 70, -58, -8, -10, 50, 119, 93, 119, -6, -115, -50, 104, 33, -25, -27, -37, -48, 85, -96, 67, 37, -96, -81, 105, 12, 65, -11, 9, 122, -23, 37, 0, 94, -10, -112, 88, 40, 94, -11, 117, -6, -19, 103, -91, -103, 38, -17, -42, 90, 55, 82, 3, 54, -56, -126, 39, 64, 73, -31, -41, 44, -99, 83, 113, 10, -51, -85, -25, -82, -39, 77, -100, -51, 18, 123, -72, -17, -61, -22, -56, 30, 110, 60, 12, -89, 84, -53, 111, 47, -100, 22, -34, -51, -56, 36, 45, 31, 98, 40, -91, 25, 27, 117, -113, 120, -105, 62, 14, -44, 76, 14, -25, 49, -120, 102, 110, -37, 75, -22, -10, 5, -116, -15, 33, -124, 80, -92, -62, -76, 121, 106, 87, -25, -26, 76, -56, -45, -107, 36, 5, 35, -17, 26, 3, 126, -101, -87, 81, -89, -15, -118, -13, -63, 111, -46, 113, -83, -103, -88, -113, 73, -41, 1, 117, 47, 87, 36, 41, -98, 117, 13, -4, 94, 49, -101, 97, -56, 119, -32, -5, 113, -14, -92, 27, -21, 118, 5, 117, 55, 123, 77, 59, 46, 29, -128, -75, -86, -30, -51, -49, -118, 80, 2, -114, 73, 59, -118, 33, -19, 1, -30, 31, -58, 89, 38, -77, 85, -3, 107, -92, -93, 118, 27, -94, -44, -57, 105, -32, -24, 65, 39, -49, -45, 118, 115, -115, -37, 74, -121, -88, -26, 25, -111, -20, -94, 89, -79, -96, 89, -100, 116, 27, -83, -105, -68, 124, 115, -91, 34, -71, 26, 81, 66, 25, -72, 68, 80, 94, -114, -113, 14, -98, 59, -69, -76, 56, -38, -128, -128, 20, 71, -18, 36, -95, 29, 41, 118, -32, -68, -92, 14, 76, 5, -101, 124, -5, -41, -99, -6, 60, 77, -90, 9, 11, -62, 75, 56, -83, -20, 127, -128, -118, -106, -11, 101, 117, -121, 62, -89, 100, 58, 24, -74, 81, 43, -80, -60, -95, -82, -58, -59, -122, 72, -104, 69, 109, -104, -11, -36, -118, -33, 96, -68, -82, -92, -59, 57, -119, 26, -61, 34, -88, -15, 36, -13, -103, -76, -76, -23, -8, 85, -78, -16, 32, 81, -55, 59, -5, 52, 114, 11, -95, -107, -59, -91, -81, -120, -107, 25, -121, 21, 91, 59, 15, 50, 111, 47, 34, 25, -114, -70, 72, 103, -39, -118, -53, 78, 119, -10, 91, -52, 47, 21, 98, 48, -108, 22, -5, -122, -5, -27, -43, -93, -106, -82, 78, -56, 31, 101, -30, 125, 33, -16, 87, -116, -21, 94, 79, -10, 73, -66, -10, 12, -107, 7, -50, 110, 21, -21, -21, -119, -112, -53, 71, -52, -84, -57, 103, 106, -83, 14, -85, -39, 120, 25, 23, 95, 77, 68, -15, -100, 22, -71, -18, 22, -82, -84, 94, -95, -13, -122, 67, -64, 52, -59, 112, -65, 20, -21, 103, 14, 64, 95, 35, -29, -61, 25, 22, -114, 88, 57, 93, -32, 68, 57, 17, -62, 12, -90, -122, -27, -53, 79, 78, -77, 27, 96, -61, -111, -12, 106, -84, -41, 95, -16, 11, -35, -83, 64, -78, 1, -100, -38, 1, 21, 82, -30, -43, -79, -68, 73, -13, -28, -77, 39, -100, -86, -86, 106, -99, -32, -50, -121, -75, -5, -11, 65, -69, 76, -54, 112, 35, 0, 108, 59, -36, 72, -88, 113, 83, -70, -61, -70, 64, -78, 59, 1, -26, 11, -19, 67, 112, -84, -95, 110, 70, -7, 91, 82, 62, 14, 8, -6, 57, 85, 60, 126, -28, 121, 1, -120, -120, 107, -25, -33, 15, 107, 17, 61, 52, -39, 113, 62, 67, 104, -89, -25, -11, -24, 106, -38, -8, 26, -119, 92, -30, -12, -47, -45, 110, 66, 22, 93, 33, 108, 115, 38, -27, -8, 43, 101, 68, -102, 20, 78, -39, 113, -118, -76, 27, 115, -4, 29, -25, -29, 67, 30, -54, 8, -21, 43, 1, -26, 38, 98, 8, -32, 20, -98, 125, -40, -123, -24, -48, -56, 23, 93, -27, -108, -11, 109, 50, 67, -51, -66, -6, -69, -81, -88, -121, 42, -58, 87, -96, -78, -112, -62, 2, -50, -68, 21, -87, 74, 99, 121, -106, -64, -15, -43, -83, 111, -115, 118, 27, 33, 108, 33, -38, 52, 86, -121, 53, 40, -23, -127, -121, -5, -37, 111, -22, 127, -124, -29, -17, -85, -122, 29, 29, -1, 96, -36, 45, -68, -81, -97, -65, -58, 102, 5, 26, 55, 57, 58, -18, 44, -83, 96, 73, 106, -73, 45, -79, 92, 8, -50, -69, -22, 94, 10, -69, -89, 87, -44, 1, -86, -86, 58, 8, -107, -56, -20, -99, -61, -121, -104, 103, 1, -103, -3, 109, -55, 125, -43, 27, 38, 88, -59, 117, 4, 10, 55, -105, 94, -20, 13, -56, -106, 109, -24, -117, 53, -92, 51, -105, -111, -79, 18, 39, -45, 83, 76, 125, 94, 86, -109, 12, 108, 10, -10, 69, 33, 81, -8, -121, 24, -5, 121, -20, 98, -80, -113, 11, 57, 35, -86, 126, 3, -47, -114, 82, -14, -73, 10, 14, 95, -108, 87, -79, 82, -29, 83, 98, 115, -7, 34, 125, -15, -63, 107, 24, 120, -106, 108, -80, -4, 111, 20, 118, 115, 44, 16, -58, 70, -93, 60, -119, -57, 7, -126, 12, 114, -86, -32, 103, 82, 122, -120, -97, -116, -35, -112, -25, -103, -88, 107, -21, 76, 83, -124, -80, 31, 67, 70, 97, -93, -80, -16, 124, -117, -11, -121, -119, -21, -107, -13, 40, -89, 75, 57, 90, -37, -101, 41, 81, 36, 9, -76, -13, 86, -46, -45, 74, -107, 100, 40, -128, -96, 51, -81, 119, -5, -84, -49, 63, 120, -122, -90, -21, -41, 113, -67, -92, 121, 88, 125, 102, -26, 89, 104, -11, 101, 14, -15, -120, 36, -116, -106, 34, -74, -5, 88, 35, 87, -127, 66, 5, 97, 104, -56, -16, -118, -111, 14, -61, -64, -113, -107, 115, -69, 51, -70, 98, -93, -121, 32, 97, -52, -36, 2, 22, -90, 113, 6, 120, -29, 16, -36, -14, 100, 118, 21, 103, -86, -28, -102, 62, 90, 12, -80, 34, -90, 53, 40, -63, 113, -26, -103, -116, 58, 27, 88, -95, -94, 58, -97, 58, -42, 113, -52, 86, -105, -51, -76, 59, 57, 113, 61, 4, 5, 102, 106, 124, -1, 125, -97, -105, 46, 66, -43, 109, -83, -2, 125, 39, -67, -117, 18, 88, -1, 60, -105, -19, 119, -15, -76, 44, 52, 28, -83, -49, 18, 45, 80, 56, -3, 69, 49, 108, 72, 125, -80, -121, -64, 91, -54, 44, -121, -89, -95, 20, -64, 14, 96, 56, -17, -120, 88, -24, 101, 96, 8, -97, -18, -63, 56, 67, 88, -64, -108, -83, 109, 115, -18, -112, -37, 31, -2, -106, 86, -121, 26, 23, -34, 18, -122, -21, -95, -101, 107, -6, 36, -94, -120, -5, 14, 30, 110, 34, -46, -58, -63, -48, 50, -7, 15, 3, 17, 89, 112, 125, -7, 122, -34, -101, -86, -7, -117, -12, -83, 102, -125, -40, 122, 38, -117, -55, 82, -87, -125, -3, -127, 91, 44, 26, 24, -87, 108, 76, 102, -96, 15, -84, 88, -12, 16, -122, -54, 60, 0, -68, -12, -53, -26, 89, -75, 56, 67, -107, 11, -128, 62, -49, 99, -61, 40, 0, -41, 74, -96, -47, -35, -128, 108, 33, 13, -38, 45, 119, 29, 70, -87, -25, -18, 38, 99, -14, -34, -78, 119, -85, -4, -26, 79, -115, -80, 63, -87, -66, -81, 41, 113, -114, 79, -10, -17, 34, 0, 5, -44, 18, -60, -49, -93, -75, -41, -73, -38, -110, -39, 104, 7, -92, -6, -11, -45, 112, -34, -64, -96, -110, -69, 77, -76, -71, -22, -116, -88, 125, 100, -41, 49, -120, 10, -17, 63, -96, 59, -43, 81, 103, -115, 120, 123, 97, -52, -5, 120, -61, 25, -31, -109, 123, 98, 113, 26, -55, 102, 5, -37, 93, -117, -113, 127, -65, -34, -59, 120, -30, 39, -101, 85, 66, 70, -58, 15, -106, 73, -4, 100, -76, 72, -30, -17, 50, 73, -48, 18, 17, -41, 127, -103, 40, -77, -2, -23, 60, -113, -25, 61, -119, -38, -58, -46, 106, 4, 63, -65, -128, -23, 79, 80, -70, -11, 87, -89, 115, 111, -48, -102, -40, -64, -75, 124, 113, 71, -75, 44, -100, 114, -59, 8, 35, 45, -40, -115, -6, 37, 108, -51, 18, 58, -26, -127, -127, 65, 31, 12, 78, -54, 56, 25, -94, 19, 55, 50, -81, -36, 104, -109, 10, -110, 2, -21, 78, 113, -6, 81, -85, 44, -119, -6, -36, 47, 105, 48, -40, 64, -80, 120, -14, 63, 112, 94, 11, -23, -97, 8, -43, 81, 1, 104, -110, 124, 46, -107, -95, 91, -27, -95, 73, -13, -128, 1, -99, 18, 107, -35, 11, -119, -108, 16, -66, -44, -44, -41, 76, -65, -2, -1, -5, 102, -121, 87, -59, -88, 3, 5, -41, 89, -124, 76, -62, -35, -94, 85, 32, -80, -30, 20, -108, -109, -128, 12, 96, 49, 16, 37, -60, -127, -68, 37, -41, -106, 45, -67, 38, -117, -46, -67, -91, -26, 24, -96, -29, 39, 121, -83, 99, -90, 99, -24, -62, 34, -48, 126, 77, 8, -17, 50, -54, -25, -18, -73, -91, 47, -76, 113, 18, 12, -39, 33, -71, 40, 63, 36, -105, -40, 110, -28, -109, 43, -65, 52, 119, 92, 29, 48, 18, -9, 125, 96, 101, -126, -64, 16, 113, 77, 65, -49, -5, -15, -111, -117, 7, -83, -1, -119, 84, 15, -91, 70, -106, -33, 117, 125, -29, 47, 108, -43, -127, -45, 13, -35, -73, -104, 67, 101, -13, 74, 32, 9, -82, 15, -61, 88, 111, 34, -47, 88, 27, -2, -31, 122, 83, 60, -24, -104, 103, 59, 83, 62, 112, -33, -118, -79, -41, 6, 20, -37, -102, -23, 67, -102, -58, 56, -42, -116, 7, 40, 28, 7, -123, -1, -85, 12, -9, 9, -26, 120, 41, -17, -16, 120, 118, -110, -37, -87, 77, 9, 104, -120, -13, 56, 87, 75, 27, 122, -10, 120, -56, 123, 45, -120, -108, 42, 104, 32, 10, 29, 1, -8, -103, 46, 0, -86, -82, 67, -81, -104, 53, -37, 39, 36, -34, -127, -32, 11, -69, -83, -108, -39, -99, -100, 51, 91, -19, 1, 45, 86, -43, -120, 92, -124, -5, -123, -13, -87, -61, 56, -90, 38, 38, 24, -37, -123, -105, 41, -21, 105, 102, -26, -27, -115, 16, -50, 79, -14, -63, 64, -108, 35, 43, -102, -13, 122, -56, 19, -119, 23, 40, 21, 113, 124, -41, 64, 29, 13, 91, -96, 15, -53, 14, -69, -100, -48, -87, 48, -43, -41, 32, -49, -17, 12, 38, 45, -3, 99, 57, -72, -89, -34, -49, -113, 108, 84, -90, -77, 101, 7, -28, 84, -41, -58, 11, -61, 111, -80, -63, 116, -6, -2, -2, 18, -110, -28, 99, -57, 9, -68, 88, 5, -73, 33, 28, -72, 56, 108, -115, -81, -64, 107, 67, 45, -12, 87, -16, 18, -36, -89, -24, -80, -45, -78, 84, 65, 95, 27, -29, 92, 105, 93, -19, -17, -109, 73, 85, -74, 108, -78, 57, 38, 24, -86, 45, 13, 125, -99, 92, -82, 93, -52, 31, -83, -110, 32, 70, -88, -36, 125, 8, 4, 110, -100, -66, -48, 8, 76, -76, 42, 5, -34, -60, 73, 55, 28, 96, -54, 106, 117, 36, 101, 99, -90, 116, 73, -57, -2, 113, -66, -15, 4, -87, -36, 35, 126, 106, -53, -61, -11, 36, -37, 42, 19, -50, 80, -19, 14, -12, -94, -14, 8, -66, -13, 64, 33, -12, -108, 67, 71, 110, -111, -53, 67, -27, 58, -73, -87, -78, 42, -111, -58, 56, 68, -67, -119, 126, -62, -58, -123, 52, -18, 13, 122, 67, 38, -61, 10, 71, -102, 37, -124, 21, -103, -58, 5, 55, 45, 99, 94, -36, -124, -15, -121, 65, 116, 19, 87, -118, -11, 117, 83, 91, -55, -113, 52, -23, 25, 123, 97, 106, -7, -116, -99, 116, -6, -75, 65, 3, 109, -117, 30, 68, -28, 102, 10, 43, -36, 113, 79, 19, 114, -71, -122, 68, -94, 122, -14, -109, -100, 127, 19, -91, 40, -24, 121, 111, 82, -97, -91, -69, 1, 119, 56, -67, 76, 110, 2, -92, 99, -80, -102, 9, 29, 9, -62, -34, 115, -83, 28, 31, 102, 23, 65, -23, 22, 75, 65, 24, 33, -102, 110, 43, -37, -127, 42, 15, 4, 31, -59, -35, -92, 115, -40, 53, -39, -39, 8, 115, -36, -74, 60, 58, -26, -54, -121, 7, 76, -24, -40, 44, 32, 66, 77, 40, -27, -107, 47, 77, -25, 41, -77, 59, -76, -57, -68, -102, -39, 63, 64, 83, -54, 122, -65, -126, 44, -106, -7, 122, -23, 13, -15, 32, -106, -46, 81, 112, -118, -15, 33, 9, -45, -104, -97, -69, -15, 111, 75, 58, -89, 28, -74, -125, 61, 105, -51, 113, 117, -53, -75, -96, 47, 24, -68, -35, 90, 87, 26, 8, 22, 20, -17, 52, 105, 89, 122, 101, 91, 29, -35, 15, -48, -27, 44, -53, -93, 10, 107, -39, 27, -33, -32, -21, 51, -80, 67, 66, 68, -22, 6, 102, -31, 95, -28, 44, 63, -77, 15, -55, 94, -14, -128, 81, -64, -115, -106, 48, -98, -121, 75, 70, 120, 5, -14, 125, -33, 47, -36, -60, -5, 55, -128, -111, -105, 76, -40, -57, 63, -71, -5, -45, -62, 24, 35, -61, 74, -50, -123, 124, 71, -70, -115, 31, 47, -67, 89, 28, 15, -17, 59, 67, 55, -75, 126, -71, -49, 104, 83, 105, 84, 126, -66, 64, 58, -88, -87, 28, 100, -16, -23, -3, 11, -91, 83, 7, 25, -54, 28, 22, -66, 77, 31, -78, -108, 59, -28, -97, 120, 94, -61, -60, 55, 107, -27, 76, -47, 28, 113, 117, -75, -16, -37, 23, 57, -58, -46, -63, -40, 35, 33, 16, -70, 105, 53, -24, 12, 56, -117, -65, -97, 66, 30, 115, 11, -37, 13, 122, -92, 0, -102, -46, -86, 70, 101, 92, 22, -31, 77, -83, -73, 29, -81, -21, 56, -34, -31, -46, 55, 18, 111, 102, -63, 82, -13, -15, 95, 86, -37, -53, 115, -46, -98, 66, -112, -65, -95, 10, -113, -51, 87, -24, 113, -119, -109, 78, -57, 48, -77, 18, -34, 28, 98, 5, -126, -23, -35, -47, -75, 29, 75, -4, 62, 24, 55, -58, -103, -119, 6, 20, 7, 93, -108, 39, -46, -31, -56, 92, 82, -53, 39, 104, 85, -79, 22, 39, 10, 116, -110, -14, 53, 28, -124, 36, 116, -64, 89, 49, -99, -97, 122, 88, 123, -113, 109, 25, -98, 47, 73, -35, 82, -77, -34, -24, -97, 90, -7, -20, -123, -85, 104, -69, 0, 25, 29, -88, -103, 76, 89, 64, 60, -5, 127, -26, -54, 59, -34, -35, 3, 102, 53, 93, -104, -66, 65, -48, 45, 88, 43, 25, -35, 109, -42, 4, -73, -51, 17, -88, -80, 116, -66, -89, -1, -76, -128, -125, -21, -90, 96, -56, -108, 94, -34, -110, -105, -31, 70, -3, -78, 32, -85, 126, 11, -103, -57, 108, 17, -19, 75, 64, -34, -42, -114, -103, 87, -85, -49, 27, 4, -97, 91, -61, 90, -111, -70, -31, 18, 7, -50, 116, 115, -48, -4, 11, 48, -6, 88, -21, 60, -49, 3, -67, -45, 29, 85, -32, 91, 90, 120, -109, 73, 105, -23, 115, 103, -56, -116, 75, -94, 26, -118, 87, 115, 101, -1, 123, -13, 117, 87, 92, -119, 117, 80, 30, -39, -82, 60, -94, 126, 10, 127, -93, -122, -54, 79, -66, -10, 52, -37, -69, -77, 72, 121, -121, 66, 14, -56, -59, 67, 87, -117, -81, 3, -66, 77, 53, 17, 117, 76, -41, 48, 89, -81, -86, -41, 89, -83, -33, -22, -83, 126, 10, 72, -95, 0, 126, -109, 22, 13, -121, -77, 1, 88, -83, -64, 29, -75, 47, 58, 92, 62, -112, -104, -5, 118, 106, 0, -115, 69, 23, -76, 44, 84, 126, -99, -70, -59, 72, 71, 21, 64, 58, 75, -95, 109, -95, -21, -84, -50, 89, 61, 101, -58, 43, -91, -23, -89, 35, 36, 124, -84, 64, 118, 92, 55, 82, 89, -77, 54, 9, -34, -71, -96, -14, -51, -99, -105, -80, 50, 111, 93, 37, 45, 75, 11, -17, 87, 28, 110, 109, -99, 112, -46, 13, -92, 16, 78, -42, 125, 95, 41, -77, 78, 24, 48, 20, -107, 120, 115, -8, 101, -107, -15, 108, -106, -28, -127, -122, 126, -95, 77, -60, 31, -66, 79, 1, -83, 101, 55, -87, 127, 89, -101, 32, -26, -41, 52, 116, 45, -53, -110, -20, 1, -68, 56, -5, -48, 12, 107, 102, -1, -40, -53, 80, -46, 72, 47, -50, -91, 24, 30, -79, 105, -88, -54, -9, -73, 25, -115, 15, -46, -89, 8, -84, 59, -11, -108, 108, 108, -52, -59, 50, -54, 68, 8, 60, -40, -41, 95, 14, 29, 36, -6, -9, -44, 84, 5, 1, -30, -10, -78, -34, -109, -18, -47, 82, 18, -9, -114, 70, -86, 97, -118, -29, -34, -25, -102, -6, 125, 50, -89, -93, 125, -108, 98, -87, 50, -113, -35, -4, -105, 16, -11, 75, -24, -118, -112, 28, 75, 69, -100, 117, 27, 101, 6, 52, 53, -22, -53, -109, -1, 5, 39, -68, 103, 17, 122, 15, 98, -91, 58, 119, -80, 113, -60, -86, -23, -108, -59, 26, 77, 124, -15, 88, -78, -103, 126, 124, 29, 115, -105, -31, 12, -1, -121, -76, 7, -112, 47, -77, 41, 34, 8, 67, 68, -23, -109, -122, 39, -13, 76, -18, 2, -25, 87, 38, 122, -65, 105, -58, -33, 63, 97, -2, 90, -101, 99, 27, 114, 65, 72, -111, -105, -72, 71, 40, -49, 93, -76, 94, 61, -70, 127, -87, -50, 110, -2, -56, 52, -127, 8, -114, -101, 110, 119, 69, -113, -10, -119, -97, -54, 86, 32, 107, -3, -2, 85, 55, 57, 127, -43, -55, 69, -108, 105, 81, 100, 61, 120, 89, -98, -87, -21, -47, 121, -122, 79, 54, 123, -125, -16, 17, 33, -74, -95, 64, 71, -14, -4, 122, -99, -25, 103, 63, 71, 52, 117, 4, -56, -31, -126, -80, -114, -68, 33, -122, 57, -92, 3, 123, -32, -108, 33, -125, -55, -44, 17, -22, 10, -52, -42, -8, -69, -36, -108, 60, -49, -125, -51, -103, 41, 104, 22, -16, 46, 45, 58, 83, -43, 69, 31, 58, 114, -13, -103, 63, -71, -112, -124, -60, -96, 42, -40, -69, 41, 3, 98, 119, -78, -47, -16, -103, 104, -23, 88, -126, 111, 103, -57, 19, 63, -70, 113, 86, -62, 54, -110, 61, -5, -66, -58, -37, -58, 43, 95, 78, -12, -28, 18, -73, -78, -78, -63, -66, 44, -43, -21, -39, -29, -1, 43, 111, -13, 83, 105, -107, -23, -62, -35, 65, -78, 52, 67, 56, -22, 36, 46, 101, -97, 62, 60, 107, 106, -78, 85, 61, 82, 11, -46, -106, -41, -4, -1, 26, 45, -8, 12, -127, -82, -85, 122, 69, -120, 49, -36, 103, 66, -21, -11, -28, -1, 17, -76, -74, 37, 25, -94, 23, 93, 87, -67, 108, 78, 12, 60, -19, -110, 123, -44, 62, -81, 116, 121, 111, -112, -17, 105, -74, 87, -91, -121, -100, -75, 32, 41, 93, 81, -64, 71, -37, 55, 120, -104, -62, 19, 124, -44, -43, 17, 86, 123, 74, -115, 41, 66, -85, 27, 23, 10, 72, 99, 99, -2, -107, 95, 62, 42, -47, 15, -94, -68, -53, 122, 44, 105, -68, -2, 72, -63, -13, -31, 62, -10, -127, 11, -32, 63, -14, -19, 55, 2, 37, -27, -72, 114, 48, 44, 90, 123, -97, -105, 15, -75, 127, -40, -54, -79, -59, -34, 110, -120, 9, 21, 69, -77, -109, -21, 75, 109, 3, 7, 1, 25, -66, 12, 64, -36, -113, 78, 82, -73, 113, -39, 77, -110, -117, 81, 1, 90, 96, 61, -54, -80, -39, -40, -54, 93, -113, -92, -59, 120, -34, 1, 60, 44, -36, 34, 110, -20, 112, 16, -39, 80, -38, 71, 109, 43, 53, -90, 85, -67, -96, -84, -11, -110, -33, -5, -40, 95, 91, 102, 88, 55, -92, -128, 120, 41, 24, -12, -104, -89, 64, -45, 127, -42, 89, 94, 26, -112, 99, 70, -9, -39, 13, -41, 104, -89, 49, -72, 88, -68, -4, 29, -8, 59, 22, 77, 43, 19, -112, 39, -124, -117, -99, 67, 12, -82, 95, -109, 83, -66, 98, 19, 105, -125, -18, 80, -70, 18, 101, 126, 90, -52, -14, -45, 48, -42, -110, 52, 18, -115, 63, 18, 10, 73, 24, 98, -124, 121, 112, -93, 126, 119, 118, -45, -80, 39, -42, 100, 55, 66, 51, 91, -65, -42, 109, 100, 80, -59, 51, 86, 19, -43, 89, 112, -17, 12, 5, -40, -116, 20, -15, -67, 43, -28, 99, 16, -44, -94, 111, 80, -124, -109, 57, 93, -111, 26, 112, 41, -82, 70, -92, -2, 105, -29, -102, -38, 90, -123, 8, -53, -4, 107, -7, 86, -70, -102, -24, -1, 69, 86, 2, -17, -122, 106, -35, -36, 123, -117, 98, 48, -25, 102, -90, 15, 54, -104, -69, 122, 9, -2, 48, -67, 107, -6, 110, 125, 15, -104, 22, 70, -66, 39, -119, -111, 4, -52, 4, 67, -112, -60, 41, -80, -118, 14, 8, 40, -58, 14, -41, 30, 30, -60, -110, -97, 15, 79, 77, 109, -50, 37, 82, 97, 40, -82, -104, 5, 113, 29, 116, -118, 38, 108, -48, -89, -9, 77, -113, -10, -57, -76, 121, -72, -118, 2, 105, 65, 121, -20, 89, 38, 120, 112, 124, 29, 4, -40, -45, -78, 52, 31, -91, -26, 57, 1, -118, 119, 72, 31, -21, 45, 87, 56, -126, 37, -46, -127, -81, -44, -104, 20, 104, -15, 88, 19, -98, -53, 53, 4, -16, -13, 68, -103, -67, 94, 117, 35, -120, -61, 8, 110, 64, -38, 110, 8, 123, -50, -46, -98, -104, -17, -121, -13, 110, -1, 114, -48, -7, -90, 85, 77, -31, -14, -112, 45, 111, 70, -44, -60, 85, 19, -60, -38, 22, 66, -125, 91, -99, -75, -59, 77, 111, -30, 7, 68, -100, 94, -7, -6, -100, 17, -47, 1, 82, -22, -110, 31, -9, 124, -78, 88, -57, 76, -83, 81, 108, 28, 57, -8, -103, -89, -56, -125, 29, -82, -88, 56, -3, 100, 22, -47, -20, 47, 114, 52, 83, 79, 80, 111, -14, 72, -41, 67, 77, 79, 31, -84, -74, -72, 42, 62, -17, 15, 109, -80, 120, 77, 80, 9, 109, -90, 23, 13, -44, 47, -42, -85, -106, 92, 15, -128, -97, -110, -122, -87, -65, 111, -25, -90, 24, 50, 19, -54, -33, 116, 127, -43, 116, 107, 86, -20, -118, -76, 114, -82, -78, -39, -88, 75, 86, -95, 22, -15, -14, -106, 127, 89, 35, -37, 101, 119, 25, 9, 102, -95, -125, -97, -115, 60, -30, -51, -11, 16, 66, 111, -11, 121, 62, -34, 63, -52, 70, 97, -68, 121, -99, -108, -51, -43, -102, -27, -12, -31, -22, 79, -106, 15, -92, -93, 93, 112, 24, -64, 40, -86, 20, 3, -61, -114, 102, 15, 4, 101, -16, 10, -127, -42, -61, 17, 80, -90, 44, 22, 57, 59, -48, -20, -11, 43, 122, 99, -2, 107, 24, 97, 49, -106, -56, 88, -27, -78, 66, -40, -106, 53, 115, -14, -30, -18, -59, -17, -60, 38, -119, -8, 89, 42, 27, 19, 10, -102, -2, -57, -40, 80, -108, -103, 49, -123, -122, 52, -15, -19, -79, 29, 124, 27, 10, 39, -1, 124, 100, -61, 30, -87, -49, -41, -4, 66, -104, 68, -49, 89, -27, -101, -51, 117, -82, -108, 14, 83, 68, 120, 87, -47, -22, -123, 76, 42, -20, -2, 104, -77, -78, -113, -89, -21, 110, 97, -97, 87, -119, -85, 120, 36, -23, -54, 106, 121, -61, -33, 108, 10, -9, 69, -66, -56, -6, -71, 107, 9, 85, -19, 80, 22, 48, 116, 91, 81, -7, 127, -29, -122, -8, 95, -18, -93, -47, 64, -62, 90, -81, 35, -11, -97, 69, -32, 77, -102, 59, -4, -98, -60, -16, -58, 57, 82, 110, 88, -32, -25, 106, -26, 21, -24, -101, 35, 107, 0, 30, 41, 125, 12, 65, -93, -108, -72, 109, -22, 46, 78, -7, -111, 7, 18, 121, 65, -76, 88, 40, -51, 105, -40, 18, 75, -21, 93, -59, 34, 42, 66, 43, -99, -103, -74, -60, 110, -61, 47, 126, 82, 78, -3, -7, -32, -4, -5, -118, 61, -20, -14, 33, -67, 104, 56, -51, 60, 74, 107, -2, 110, -36, -48, -110, 2, 48, 123, 72, -68, -89, -119, 91, -27, 64, 66, -120, -77, 29, 39, -51, -45, 46, 104, 98, 17, 22, 100, 55, 49, 49, 49, -96, -83, -49, 125, -78, -63, 107, -86, 107, 55, 73, -54, -20, -95, 34, -119, -32, 56, 48, -62, 66, -98, -125, -61, 6, -77, 15, 32, -124, 119, -30, -29, 9, -20, 25, -86, -9, -79, 92, -12, -101, 60, 82, 73, -118, 26, -83, 37, -102, -26, -37, -69, 0, 36, 120, -4, 104, -123, -56, 60, -45, 125, 14, -51, -121, -99, 122, 58, 111, 16, 107, 88, 3, -120, 76, -88, -47, 84, 0, -58, 77, 86, -121, -52, 106, 58, -64, -41, 2, -128, 37, 49, -46, 24, -19, -29, 56, 23, 99, -18, 32, 43, -87, 61, 47, -27, 51, -24, 111, 5, -113, -34, 53, -77, 3, -61, 40, -111, -121, -33, -103, 126, 84, 31, 107, 24, 20, -32, -61, 112, 74, -7, -14, -120, 42, 42, -55, 75, 59, -35, -120, -33, 77, -106, -44, -53, 54, -87, 22, -34, 64, 42, -102, 0, -34, 7, 126, 64, 99, 45, 53, 123, 102, 122, -119, -108, 9, -96, 113, -12, 90, -25, -87, 96, -52, -22, -123, -63, 35, 28, 10, -114, 53, 59, 126, -32, 1, 43, -18, 42, -49, 118, 117, -88, 12, 29, 9, -50, 21, 7, -71, -83, -13, 120, 87, 86, -98, -73, 108, 28, -48, -62, -72, 117, 73, -12, -28, -49, -115, -116, -103, 102, -115, 6, -93, -109, 58, -49, 30, -59, 36, 112, 73, -86, -4, 38, 108, 88, -14, 96, 58, -117, -10, -80, 24, 108, 21, -32, -14, -100, 74, 72, -27, 34, -68, -3, 118, -59, 122, -95, -83, -80, 121, -52, -115, -90, 64, -12, 90, -35, 71, -103, 32, 22, 25, -70, -82, -79, -101, 71, 108, 82, 97, -44, -118, 65, -57, 69, -9, 52, 64, -62, -1, 94, -62, 121, 36, 20, -72, 123, -35, 50, -21, 98, 92, -119, 26, -56, 2, 63, -26, 4, -73, -88, 69, -126, 44, 115, 80, 17, 116, 103, -4, 109, 19, -5, 64, -36, 77, -99, 5, 11, -38, 76, -99, 12, 124, -55, 107, 35, 64, -7, 92, 77, -21, -10, -54, 25, -125, -75, -53, 7, -27, 80, 63, -47, -44, 62, -76, -94, -28, -34, -112, 123, -85, -110, -65, -59, 27, -67, 57, 76, -92, 9, 1, -13, -109, 18, -88, -116, 12, 117, 4, -74, 33, -109, 71, 64, -22, 113, 1, 91, -72, 102, 124, -65, -22, 66, 94, 32, 119, 9, -102, 119, -117, -60, 118, 100, -63, -39, -81, 42, 5, 36, -35, 104, 85, 120, -44, 93, 117, 44, 17, 16, -34, -75, -110, 69, 78, 73, -127, 5, 16, 121, -121, -57, -46, -115, -13, -101, 103, 118, 126, 30, -58, -122, -7, -47, -20, -54, 109, 89, 126, -127, 72, -78, 43, 8, 39, -49, -75, -77, 114, 89, -74, 124, -32, 10, -10, -54, 121, -22, 18, -61, 33, 100, -67, 48, 104, 98, -89, 82, -27, 33, -32, -63, -43, 58, 52, -83, 34, -18, -41, -70, 75, -15, 81, -57, -66, 122, 127, 52, -42, -103, -80, 10, -32, -85, 86, -96, 74, -28, -36, 89, -81, -67, -120, 117, 68, -119, 109, -110, 10, -128, 64, 93, 52, 91, -63, -71, -105, 87, 123, 1, -104, 64, -107, -40, -31, 98, 117, 3, -68, 48, 88, 11, -27, 113, -68, 4, 32, -64, -123, 83, -115, -80, -59, -67, -83, -120, -91, 115, -119, 21, -123, 105, 1, 71, -104, -39, -14, 68, -56, 119, 48, 77, 10, -15, 58, -17, -74, -37, -18, -33, 81, 109, -123, -61, -127, -57, 43, -37, -29, 72, -75, 110, 91, 105, 12, -115, -90, 81, -16, 33, -84, -42, -111, 17, -104, -79, 28, 6, -86, -86, -34, -116, 11, -74, 39, -32, -73, -55, 92, 6, 31, 29, 78, 27, -55, 80, -56, -22, 49, 43, -39, 97, 32, -86, 59, 57, 18, 126, -117, -64, 121, 119, 67, -110, -1, -51, 122, 1, -11, -126, 71, 20, -58, -92, 97, 17, 46, -38, -58, -70, 42, 16, -19, -86, 28, -54, 118, -122, -107, 74, 71, 12, 50, 77, 29, -124, -106, 125, -47, 50, 97, 18, 114, 41, -121, -84, -127, 45, 40, -60, 58, -119, -22, 68, -57, -1, 16, 68, 75, 126, -31, -67, 29, 16, -21, 15, -87, 116, -43, 71, 30, -95, -52, -57, -87, -20, -120, -15, -85, 117, -37, 41, -93, -19, 13, -74, -71, -86, 8, -65, -47, 127, 97, -6, -11, -125, 119, 124, -20, -61, -90, -82, -125, -128, 111, -84, -45, -23, 124, 85, 109, -66, -46, 74, 16, 44, -6, -31, -19, 35, 78, 94, 48, -72, -88, 67, 118, 17, -43, -42, 15, -61, 124, 15, 73, 13, 95, 64, 27, 28, 73, -31, -109, -84, -2, 118, 70, -111, -95, -91, 1, 49, -80, 54, 35, -56, -109, 126, -73, 102, -34, 32, 104, 42, 46, 33, 3, -91, -110, 20, 2, -55, 63, -58, 55, -82, 76, 88, -120, 84, -73, -36, -8, 104, -80, 20, -117, 98, 57, -64, -24, 66, 86, 64, -39, -23, -33, -43, 114, 3, -70, 73, 86, -108, -76, 116, -93, -48, -41, -42, 22, 13, -89, 61, 28, 91, 31, 43, -89, -71, 24, -87, 108, 77, 22, -46, 16, -76, -75, -122, -38, 14, -82, 127, -6, 60, 64, -67, 54, 117, -116, 69, -46, 55, 16, 11, -2, 5, -88, -60, -84, 106, 84, 53, -85, 46, 83, 122, -3, 33, -16, 71, -100, -124, 82, 89, 67, -13, -78, 106, 123, -94, 108, -24, 73, -89, 74, -20, 77, -103, -126, 92, -55, 49, -117, -41, 110, 47, -124, -103, 91, -46, -121, -41, 25, -95, 30, -87, -67, 100, 60, -101, -28, 51, -95, 117, -86, -47, -30, -1, 105, -77, 39, 78, -97, 58, -59, -22, -115, 32, -89, 118, -32, -78, 28, -58, -16, 26, 65, 78, 44, 16, 78, 72, 34, 52, 108, -40, -81, 100, -71, -8, 64, -1, -15, 113, -41, -85, -6, -71, 32, 77, 105, -55, 38, 32, 91, -3, -42, 87, -121, -61, -6, -30, -33, -65, 127, 57, 57, -83, 41, -114, 75, -116, 64, 20, 18, -4, 22, 24, 51, 59, 31, -55, -72, 44, -13, 17, 40, -28, -93, -88, 1, -6, -60, 105, 59, -85, -117, 102, -69, -79, -43, -116, 106, 60, -98, -6, 101, -12, -95, -120, 0, -99, 99, 102, 9, 17, 82, 56, 102, -44, -66, -26, 126, -30, -99, -31, 39, -106, -6, -27, -32, -30, 21, 81, -62, 48, -121, 125, -78, 105, -4, 57, 28, 21, -1, 121, -26, -117, 18, 54, -122, -21, -10, -6, 70, -122, 114, -43, -69, 12, 57, 60, -114, 83, -106, -110, -52, 124, -40, -117, -118, 48, -68, 115, 8, -122, -89, -30, -58, -44, -105, -99, -104, -58, -66, -99, -81, -119, -24, 57, 98, -90, 8, -47, 32, -8, -87, -111, -35, 0, 66, -105, -73, -45, -121, -98, 111, 58, 44, -48, -75, -96, 76, 71, -36, -123, 71, 103, 94, 102, -29, 26, 12, -82, 8, -4, 45, -85, -52, 78, -31, 125, -42, 5, -9, -105, 124, 110, 95, -65, 105, -128, -116, -7, 25, -117, 35, 5, 35, 61, 101, 5, 12, -73, -54, 10, -18, 74, -29, 9, -89, 43, -102, -33, 30, -119, -16, -83, 43, -40, -61, -39, 19, -2, 115, -102, -51, -47, 66, 31, -85, -23, 33, -30, 36, 104, -1, 32, -11, 42, 98, 79, 77, 102, -59, -16, -78, 104, -123, 110, 81, -113, 80, 100, -90, -49, -32, -41, -51, -97, -120, 35, 4, -56, 71, -97, -21, 78, 109, -122, 68, -20, -85, 32, 67, 91, -92, -84, -59, 68, 23, 64, -124, -33, -34, 20, -121, -31, 106, 112, -62, 69, 47, 122, 51, -76, 73, -9, -101, 9, 95, -92, -18, 5, -67, -77, -21, -107, -101, -127, -89, -13, -110, 6, 94, 106, -107, 40, -64, -58, 27, -8, -66, 46, -89, -43, -103, -96, 93, -3, -109, -37, -16, 89, 106, -48, 85, -74, -60, -51, 11, -117, 25, -125, -104, -57, -88, 50, 55, 2, -127, -38, -90, 123, 31, 42, -39, 96, 9, 5, -28, -46, -49, -7, -98, 10, -84, 114, -109, 115, -5, -18, 106, 48, -88, -74, 41, -114, -105, -32, 98, -19, -82, 107, 103, 30, -110, -35, -17, -87, -56, -123, 80, 62, -97, -24, 116, -97, 66, -4, -70, 87, 44, -42, -43, 43, 90, -18, -64, -16, -43, -3, -64, -49, 28, -61, -124, -102, 92, -44, 8, 98, -62, 36, -22, -82, 119, -29, 6, 33, 36, -66, -58, -2, 19, 21, -47, -94, -68, -111, -75, 115, -69, 125, 22, 7, 68, 105, -90, 94, 46, 0, 88, -103, 11, 38, -60, 85, -127, 16, 13, 79, -122, -73, -77, 121, -127, 94, -105, -5, -11, 45, -109, 25, 43, -8, 81, -10, 94, 34, 51, -53, -46, -81, -125, 87, -100, -100, -23, -13, 122, 108, 13, -32, 10, 35, 96, 49, -100, 108, 40, -5, -5, 5, -1, -39, -53, -43, -15, 55, 98, -70, -51, 56, 28, 93, -108, 63, -7, 54, -63, 37, -92, 60, 17, 120, -128, -101, 97, 121, -52, 50, -72, 125, -106, 54, -79, 64, 127, 13, 11, -89, -120, 115, -37, -16, -2, 8, -15, 112, -57, -1, 122, -23, 61, -40, 81, 91, -6, -125, -30, 59, -106, -57, 4, 82, 125, 51, 119, 89, -45, -120, -93, -106, -46, -93, -112, 27, -64, 96, 101, 38, 81, 47, 101, -20, -41, 116, -124, -51, 22, -113, 69, -83, -69, -105, 35, -48, 72, -119, -63, 101, 35, 71, -57, 99, -20, 120, 46, 98, 120, 41, -62, -125, 60, -8, -55, 110, 3, -28, -31, -80, 42, 92, 35, 69, 41, 123, 105, -26, 34, 100, -13, 68, 41, -91, 67, 36, 7, -58, -69, -124, -69, 76, 29, 59, -77, -116, -31, -128, 31, -99, 56, 26, 100, -18, 9, -95, -78, -26, 6, 35, 110, 103, 6, -59, 112, 61, -96, 51, 116, 99, -127, 12, 73, 73, 1, -56, -105, 79, -82, -123, -76, 92, -128, -51, 64, 46, 111, -16, -72, 100, 54, -86, 15, -123, -113, -113, 5, -99, 7, -106, -37, 55, -34, 120, 93, -15, 15, -29, -125, 12, 111, 15, -10, -51, 97, -83, -105, 9, 87, 5, 62, -34, 118, 74, 8, -53, -112, -104, 0, -84, 102, 99, 84, 122, -64, -125, 117, -109, 12, -3, 100, 84, 15, -15, -33, 80, -3, 94, -97, 110, 62, -102, -1, 112, 28, -82, -113, 69, 78, -82, -45, 34, 0, 127, -110, -102, 77, -81, 85, 7, 3, -75, 5, -25, -37, -54, -77, -39, 51, -78, -18, -14, 100, 91, -60, -18, 37, 14, 13, 16, 4, 20, 99, 118, -51, -44, 18, -114, 36, 17, -5, 56, -10, 5, -118, -43, 98, 68, 3, 13, -22, -92, -120, -22, 19, -89, -114, 18, 65, -92, 16, 70, 86, -96, -128, 63, -6, 102, -100, 57, 94, -39, -24, 6, 103, 102, 27, 94, -27, 85, -65, -125, 86, -124, -99, 10, 1, -43, 43, -89, 97, -28, 107, -95, -53, -1, -63, -91, 91, -33, -39, -47, 67, -49, 69, -9, -61, -87, 116, 29, -47, 117, 118, 115, 28, 43, 111, -79, -88, -119, -97, 113, -96, 67, -94, 34, -51, -5, -29, 88, -61, 99, 97, -55, 9, -4, -34, -73, -76, -16, 25, 70, -80, -113, -35, -62, 90, 57, 29, 85, -58, 80, 108, -33, -83, -127, -13, -13, -125, -52, -50, 19, 121, -45, 50, 43, -51, -71, -18, 74, 10, 50, 95, -74, 110, -90, -46, 123, 19, 18, 58, -22, 91, -73, 108, 13, -116, 43, 87, 29, 60, 126, -97, 111, 39, -29, -70, -111, -13, -72, -39, -80, 92, -74, -67, -21, 49, -96, -120, 106, 41, -79, -62, 116, -99, -95, 36, 106, 57, 73, -24, -34, -64, 59, 86, -23, -37, -56, -42, 91, -121, 101, -87, 97, 61, 72, 27, -110, 112, 127, 95, -113, 57, -106, 122, -28, -29, -57, 56, 34, -60, 69, -13, -62, 11, -7, 98, -109, 93, 105, -23, 78, -14, -27, 126, 112, 34, -85, -3, -10, 35, -122, -109, 59, -74, -120, -104, 15, 122, 37, -123, 101, -20, -42, -36, 112, -112, 91, -70, 90, 52, 17, -61, 53, -58, 115, 28, 107, 28, -68, 118, -106, -71, 33, -103, 84, -63, -60, -34, -19, 65, -24, 24, 84, 111, 92, -34, 123, -125, -86, -27, -65, -23, -89, -33, -66, -119, -101, 1, 54, -71, -47, -6, -8, 116, 97, -65, -125, 104, -65, 86, 94, -72, 46, 29, -36, 70, -66, 92, 89, -59, -14, -114, -85, -22, -121, 22, -126, 103, -35, -40, 12, 115, 122, -125, -127, 122, 48, 18, -113, -22, 18, -108, 90, 24, -55, -30, 30, 111, -83, -40, -120, -26, 78, 95, 64, -68, -64, 96, 101, -21, 90, 44, 29, 126, -101, -43, -28, 16, -127, 86, -27, -25, -120, -56, -101, 3, -121, 25, 51, 86, 55, -122, 35, -7, -8, 89, -83, -123, -120, 61, -42, -27, -32, 96, -107, -51, -1, -72, 77, 91, -19, 16, -41, 23, 50, -29, 55, 51, -74, 80, 31, -35, 36, -103, -9, -67, -66, -1, -1, -32, -103, -63, 105, -101, 100, -108, 26, 93, -76, -55, -1, -49, 12, -66, 59, 10, -45, -74, 74, -83, 18, -53, -66, -61, -79, -44, 123, 67, 48, -52, 30, -34, 79, 82, 45, -16, -45, -23, 83, 120, -103, -37, -7, 31, 19, 12, 88, -84, -20, 40, 123, 56, -22, 24, -80, -118, -122, -121, -96, -81, 85, -80, -79, 114, 71, -106, -93, 65, -34, 78, 120, 68, 82, -46, 61, -85, -5, -17, -12, 52, -66, -51, -56, 106, 92, 97, -22, -111, 98, 73, -49, -22, 114, 27, -116, -28, -107, 86, -9, 100, -115, 83, -111, 39, -5, 27, 52, 57, -101, -62, 124, 27, 40, -23, 10, 32, 125, -12, -70, 23, -104, 72, 50, 81, -100, -128, -103, -75, -50, -8, 16, -85, 98, 75, 119, 37, 83, 38, -8, -116, 114, -54, -76, 7, -27, 20, -106, -64, 85, -121, -92, 58, -13, 26, -117, 100, -6, 45, -39, 116, 25, -1, 11, -7, -100, 3, -125, 69, 64, -128, 22, 36, 112, -99, -107, -115, -86, -51, 55, -128, 61, -108, 51, -94, -11, 1, -74, 122, 127, -37, 69, -70, 121, -42, -56, -45, 15, 88, 75, -98, 16, -90, -53, -19, 34, -105, -47, -1, 26, -10, -118, -23, 24, 70, -14, 10, 63, -44, 59, -118, 101, -74, -28, 82, -107, 104, -80, -94, 47, -3, -72, 15, 35, -41, 33, -86, -109, -39, 10, 22, 1, 67, 95, -67, 70, 46, 72, 55, -12, -9, 80, 110, -90, 69, 33, -53, -89, 52, 40, -25, 12, -24, 26, 34, 103, -14, 47, 85, -86, 64, -15, 45, -58, 73, -32, -80, 116, 59, 57, 15, 73, -62, -97, 3, 39, -23, 49, -3, 90, 100, 116, 101, 126, 6, 71, -114, -9, -111, -93, 121, 74, -128, -89, -9, 94, 59, 25, 108, 97, 97, 13, 7, -35, -61, -64, 11, 4, 36, -119, 1, 26, 69, -61, -38, 62, -119, 17, 49, -41, 77, 16, 0, -18, -65, 70, -29, 20, 59, -43, -5, -46, -47, -6, -90, 34, 39, 97, -95, -28, -11, -98, 30, -44, -87, -86, 115, 10, -20, 86, -6, 17, 5, 79, -112, 98, 106, 78, 66, -36, 14, 91, 120, 103, -11, -47, 49, 90, 115, -57, 103, 33, -94, -124, -51, 47, 32, 10, 37, -107, -107, -82, 87, -83, -61, -40, -69, -58, -103, -7, -7, 75, -71, -22, -62, 59, -41, 95, 55, -38, -33, 75, -107, 19, -68, -79, 10, -18, -94, -7, -52, -91, 97, -98, -62, 16, -120, 63, -28, -72, 76, -93, 105, -110, 0, 22, -124, 75, 4, -57, 6, -10, -90, -37, 26, -4, -18, 111, 15, 125, 88, -124, 82, 98, 101, -53, -64, -12, -108, 64, -75, -12, 16, -14, -40, 60, 124, 26, 41, -47, -69, 107, 88, 85, 0, 66, 15, -50, 90, -15, 102, 6, 120, 81, -60, -85, -3, -46, -109, -43, -38, 81, -88, 50, 5, -58, -76, 67, 11, -69, -40, -5, 103, 60, 13, -120, -61, 104, 42, -104, 89, 46, 76, 119, 98, 37, 40, 118, 87, -96, -40, 26, -73, -86, -57, 33, 63, -25, -104, -17, -70, 60, 4, 16, 33, 68, -47, -30, 33, 70, 12, 122, 109, -108, 22, 47, 22, 69, -24, -98, 58, 112, 119, 32, 46, -86, -111, -127, 107, 25, 116, -114, 7, 79, -128, -63, 87, -124, 77, -52, 112, 92, -74, 72, 57, -27, -44, -73, -94, 65, 13, 32, 97, -113, -107, -34, -74, -6, -81, -32, -110, -53, 7, -19, -91, -84, -8, 40, -40, 86, 88, -7, 52, 88, -115, 66, 100, 115, -37, 12, 119, 21, -41, -119, 0, 48, 12, -1, -86, -113, -54, -18, 43, -98, 68, -65, 64, -64, -84, -104, -108, -75, 53, -52, 92, -107, 62, 55, 57, 38, 72, -89, 21, -118, 110, 76, -71, -113, -126, -86, 126, 114, 31, 110, -123, 89, -55, -20, -125, -90, -3, -92, 108, 117, 75, -97, -39, -47, -120, -7, -11, -95, -34, -53, -34, 123, 77, 14, 24, 37, 80, -60, -102, -80, -22, -22, -63, 112, 14, -87, -45, 59, -37, -2, 18, 21, -51, -53, -58, 30, 108, -57, -121, -53, -7, 46, -6, 64, 124, 97, -43, 61, 28, 70, 56, 90, -55, 114, -48, 73, 52, 39, -105, -123, -25, 63, 99, -58, 40, -12, -113, 45, 58, 22, 110, -84, 92, 20, 51, 38, 18, -107, 73, 92, 17, 58, 124, -117, 42, -45, 46, 54, -8, 5, 28, 74, -70, -99, -29, 27, -117, 40, 26, -31, -51, -15, -82, -53, -107, 95, -115, -30, 9, 48, -32, -20, -68, 26, -80, -51, -85, 73, -70, 0, -85, -34, -73, -61, 89, -101, 86, -8, 8, 65, 22, 37, -67, 6, -85, -60, 0, 99, 95, 32, 114, 18, 65, -107, -4, -26, -55, -3, 76, -111, -1, -90, 103, 0, -84, -14, 85, -38, -88, -58, -70, 111, -15, -59, -82, 97, 67, 7, 115, 57, 107, -51, 46, 66, -49, 69, -13, -18, -7, -56, 29, 69, -11, -127, 57, -115, -4, -83, 8, -78, 103, 10, -121, -6, -91, 70, 39, 106, 20, -111, 102, -43, 43, -89, 9, 63, -109, 86, 86, -125, -125, -15, -16, -31, 84, -27, 101, -13, 10, -26, -61, 20, 113, 109, -70, -36, -69, 61, 14, -103, -123, 55, -73, 71, 75, -17, 48, -55, -10, 117, -125, 3, -66, 5, 93, -56, -111, 21, 9, -61, 14, 37, -42, -103, 30, 23, -65, -59, 40, -57, -119, -120, -60, -69, -14, 126, -87, -50, -1, -32, -57, -17, 86, -46, -104, -108, -26, 100, 59, -63, 94, 119, 101, 3, 41, 112, -62, -91, -18, -31, 3, -99, 59, -121, -91, -59, 27, 30, -100, -57, 81, 73, -9, 99, -34, -11, -8, -64, -35, 23, -31, -25, 25, 11, -111, -106, 104, 9, 99, 111, -86, -47, 95, 77, 112, -125, 119, 54, 87, -51, -50, -48, -57, 15, 7, -18, -110, -20, 127, 63, -46, -53, 72, -111, 52, 110, -81, 78, -71, -61, 26, 120, 46, 84, -27, -72, -63, -17, -72, 4, 42, 95, -68, -5, 63, -123, 107, -24, -14, -27, 88, -106, 27, 43, -114, -84, -39, -23, -11, 14, 16, -35, 21, 15, 81, -7, 27, 17, -58, 44, 56, -45, -6, 98, 67, 48, 123, -22, 100, 9, -34, -49, 95, 123, -26, 116, 57, -11, 77, -47, 22, -16, -5, 92, 99, 36, -2, -22, 39, 58, -46, -25, 79, 63, -30, -6, -56, -43, 80, -7, 120, 42, 37, 110, -54, -98, -9, -84, -121, -59, 18, 34, -60, 98, 16, 104, -128, 3, -65, 37, 89, 7, 25, -34, 107, 123, -99, 46, 50, -99, 105, 73, 82, 70, -53, 103, -120, 42, -50, -26, 6, -4, -40, -105, 53, 24, -39, 69, -128, -29, -58, 5, 26, 32, 58, -80, 7, 22, 18, 66, -119, 4, -12, -28, -46, 111, 20, 16, -73, 19, -23, -93, -54, 11, 46, 82, -63, 9, -48, -37, 21, 118, -25, 8, -119, -14, -52, -86, -102, 101, -82, -27, 9, -106, 31, -73, 1, 88, -111, 38, 53, 41, 26, 37, -123, -122, 80, 78, -119, -37, 93, -57, 97, -65, 87, -48, -121, -122, 56, 120, 36, 116, -69, -55, -58, 103, -99, 119, 52, 46, -77, -91, -38, 26, 39, 118, -72, 90, -117, -25, 72, -103, 47, 18, 37, 114, 66, -2, -120, -60, -22, -10, -21, 96, -33, 76, -102, -56, 41, 4, -57, -27, -24, 3, 112, -95, -22, -54, -29, 12, -127, -6, -49, -108, -124, -53, -91, 96, -45, -28, -21, 54, 9, 42, -82, -42, 107, -29, -60, -59, -77, -51, -16, 115, 123, -13, 126, 88, -31, 39, -68, 108, -59, -91, 62, -21, 56, 108, -113, -18, -93, 101, 78, -42, -11, -41, 11, 17, -40, 120, -86, -45, 29, -22, -54, -127, -121, 76, 11, -86, -74, -99, -53, 91, -4, -50, 95, 127, 79, -5, -35, 91, 107, -94, 75, -21, -67, 96, 4, 62, -61, 87, 14, -14, -68, -29, 94, -106, 126, -127, 109, 78, -40, 71, -73, -98, -117, 17, 18, 7, -34, 39, -81, 19, 22, -67, -81, -26, 10, -101, -104, -39, -7, -32, 0, 1, -5, 113, 115, -104, 82, -35, -58, 62, 3, 36, 21, 45, -119, -3, 38, 52, 39, 66, 88, 102, 62, 111, 69, -10, 67, 40, 51, -106, -14, -19, 24, 29, -12, -54, 74, 48, 27, 101, 122, 56, -111, -127, -76, -33, -34, 16, -28, -83, 48, 118, -80, 38, 122, 36, 62, 51, 64, 40, 26, 46, -3, -90, 119, 80, 28, 91, 5, -83, -16, 47, 115, 19, -101, -52, -103, -42, 48, -57, -45, -128, 116, -100, 91, 23, 30, 1, -85, -112, -23, 90, -81, -2, 90, 42, 71, -73, -8, 23, -122, 78, 78, 102, 12, -87, -58, 95, -52, -90, -121, 102, -61, 84, -16, -48, -77, -25, 77, 37, 88, 7, 43, 96, -116, -53, -3, -52, -76, -45, 70, 25, 119, -53, 87, 98, -95, 77, 78, 57, 49, -49, 91, 41, -120, 102, 81, -39, 52, 127, 125, 18, -83, -5, -58, 26, -17, 31, -52, 52, 68, -8, 17, -113, 26, 84, -120, 106, 42, 19, 46, 24, 107, 32, 127, -66, 54, -2, 68, -67, 103, -100, -79, 51, -104, -35, -103, -77, 94, 89, -100, -42, 52, -74, -6, 78, 101, 38, -67, 84, -4, 60, 101, 78, -19, 102, 33, -92, 113, 85, -72, 78, -40, 44, -104, -16, 101, 42, -97, 8, -14, -26, -43, 20, 60, 61, -123, -72, 7, 19, 113, -98, -18, -42, 16, 111, -55, -104, -36, 105, 95, -99, 122, 34, 72, 6, -92, -88, -14, -92, 64, 74, -72, 5, 24, -19, -77, -49, 45, -64, 76, -79, 57, -82, -97, 112, 16, -55, -31, -17, 117, -17, 42, 113, -50, -1, -110, -62, 3, -87, 3, 91, -41, 67, -111, 79, -23, 77, 55, 15, -56, -1, -85, -50, 24, -12, -16, -105, 37, -3, -28, 17, 112, -88, 22, 82, -33, -11, -70, -110, -45, -122, -10, -94, -19, 29, -119, -48, 7, 90, -116, 41, 0, 93, -100, -41, -18, -33, 16, 103, -128, 98, -116, -111, 88, -93, -125, 4, -82, -90, 35, -24, 38, 27, 17, 77, -36, 29, -90, -70, 65, 100, 35, -84, -122, 62, 121, 109, -42, -73, -64, 64, 62, -40, -120, 116, 113, 35, 105, 31, 94, -24, -67, 22, -5, 41, 44, -49, -90, -22, -42, -126, 5, 42, 23, 22, -112, 46, 48, 73, -84, -3, -71, 31, -126, 30, 35, 52, 83, -72, 79, 104, -73, 37, 74, -52, -4, 2, 87, -93, -22, 17, 61, 39, -30, 2, 93, 10, 86, -45, 45, -117, 78, 105, -79, -84, 86, 36, 116, 0, -76, -31, -97, -100, -109, -62, -110, 38, 122, -7, 90, -17, -105, -112, 97, -124, -62, -17, 14, -86, 119, -20, 90, 19, -86, -115, 82, -41, -55, 87, -25, 76, 61, -9, 5, -68, 102, -100, -12, -49, -12, -110, -83, -86, 80, 11, -27, 86, -31, 96, 84, -36, 69, 82, 11, 75, 59, 98, -95, 127, 84, 100, -83, -115, 61, 61, -29, -42, -85, -9, -39, -90, -73, 96, 44, 103, -55, 52, -60, -9, 107, -43, 58, 14, -58, -5, 7, -95, -82, 70, 15, -22, 1, -51, -69, 12, 37, 71, 86, 86, 112, -55, 125, -63, 0, -5, 40, 72, -36, -31, -22, 115, -100, -6, -119, -34, 91, -72, 69, 110, -8, -17, 13, 38, 28, 65, -74, 113, -9, -56, 107, 102, 44, -41, 102, -74, -101, -68, -97, 59, -77, -56, -29, -79, -119, 11, -113, 83, 18, 79, -81, 92, 63, 20, 0, -53, 48, 71, 97, -15, 41, -25, -125, -54, 23, -15, -112, -110, -21, -83, 106, 37, -44, -41, 43, 86, 113, 120, -51, 42, 87, -83, 82, -110, 21, 18, 70, 115, 16, 57, 0, -56, 86, -34, -66, -41, 88, 89, -45, 72, 85, -38, -106, 17, 103, 104, 12, -74, -93, -99, -127, -27, -66, -34, -91, 24, -88, -35, -86, -117, -109, 72, 36, -79, 6, 57, -87, 82, 68, 70, -122, 22, -52, 37, 47, -29, -110, -64, -109, -60, 72, -73, -53, 67, 27, -78, -122, -22, -86, 30, 32, -113, 121, 32, 105, 8, -100, -38, -20, -75, -17, 122, -111, -114, -3, -113, -98, -16, -1, -52, 67, -104, -123, 79, 73, 115, -33, -123, -96, -79, -75, 123, 41, -20, -115, -66, 19, -94, -5, 85, 52, -91, -116, 84, 2, -12, -112, -110, -78, 93, 68, 100, 44, 106, -40, -124, -38, -115, 112, 75, -24, -105, -92, 50, -2, 103, -55, -24, 61, -43, 2, 114, -26, -102, -111, 25, 112, -3, 76, -90, -50, 66, -120, -87, 104, 66, -8, 95, -53, 6, -41, -48, -11, -92, 121, 25, -41, 66, -80, -77, -35, -89, 70, 35, 69, 13, 18, 125, -53, -50, 24, -100, -10, -62, -46, 94, 64, 40, 57, -122, -85, -32, -52, -32, -89, 125, -85, 110, -6, 42, -34, -81, -87, -121, 76, -86, 77, -114, -73, -88, 106, 38, 98, -41, -55, -102, 37, -76, -3, 125, 66, -26, 46, 42, -120, 83, 107, -49, 105, 80, -92, 4, 1, -107, -51, 22, -120, 74, -23, 25, -93, 83, 114, 63, 84, -5, 99, -123, 47, -107, 121, -43, 8, 90, 108, -77, -41, 34, -17, -81, -85, 41, 77, 79, 40, -127, -8, -42, -5, 124, -102, 35, -17, -29, -20, 98, -75, -63, 45, 21, 43, 26, -89, 48, -37, -9, 10, 1, -127, -13, 80, 69, 68, -25, 95, 77, -21, -49, 78, -112, 83, -72, -116, -75, -23, 89, 79, 115, -43, -115, 121, 49, 58, 20, -88, -72, -63, -93, 9, 59, -81, -6, 84, 91, -6, -98, -105, -100, 80, 5, -44, 59, 46, -54, -70, -70, -115, 0, 127, -126, -98, 95, 123, -83, 78, 73, 64, -55, 21, -91, 90, 81, 111, 64, -73, -120, 86, -44, -97, -128, 46, -99, 55, -21, -23, 47, -29, 29, 67, -63, -54, -33, 16, -126, -49, 80, 57, -128, -98, -60, 57, 83, 84, 70, 122, -6, 105, -36, -102, 82, -109, 38, -46, -66, -3, 20, 65, 70, -49, 56, -44, 48, 46, 27, -25, 51, 28, -80, 68, 24, -39, 35, 99, 117, 76, -3, -88, -2, -11, 123, 50, 27, 126, 13, 112, -108, 57, 127, 94, 117, 126, -104, 113, 107, 90, 76, -99, -62, 97, 12, 18, -39, 26, 9, -3, -62, 116, 11, 110, 16, -39, 77, -65, -119, 24, 75, -86, 38, -30, -98, 28, 10, 113, 34, -83, -62, -100, 41, -21, 37, -19, 73, -127, -127, 5, -114, 58, -41, -98, -79, -124, 28, -128, 79, 14, 67, 63, -77, 77, 8, -86, 36, -98, -82, -41, -128, -32, 126, -115, -96, -121, 66, 12, -28, -126, 3, -74, -22, 105, -12, 8, 127, -2, 98, 8, -54, -31, -80, 63, 93, 117, -41, -75, -120, -92, -113, 47, -8, -76, 20, -114, 107, 94, 95, -48, 20, -62, 15, 68, 80, 111, -128, 87, 115, 18, 15, -31, -36, 73, 21, 0, -18, -50, -108, 109, 25, 123, 89, -38, 67, -35, -109, -23, 2, -69, 43, -27, 36, -5, -78, -91, -57, -87, -60, 108, 89, -81, 50, 125, 68, -69, 18, 40, -29, -20, -23, -46, -122, -1, 44, 34, -64, 6, -57, 86, -79, 11, -83, 67, 115, 73, 68, 122, 99, -60, 65, 57, -85, -102, -49, -41, 32, 105, -70, 54, -25, -58, -85, -51, 124, -53, -9, 40, 58, 38, -90, -8, 49, -25, -60, 106, 117, -122, 120, -6, 109, 12, -80, -110, 80, 79, -25, -107, -9, -104, -53, 66, 51, -1, -10, 76, 36, 112, -19, -27, 111, -4, 54, -103, -128, 73, -99, -82, 72, -51, 122, 57, -88, -48, 94, 15, 62, 37, -51, -46, 46, 54, -25, -66, 85, 38, -123, 119, 8, -68, -8, -22, -51, 76, -94, -102, 30, -13, -94, -36, 126, 89, -56, -54, -93, -29, -27, -74, 99, -16, -90, -40, -60, -86, 18, 64, 58, 123, 110, -104, 119, -122, 57, -64, -17, 40, -61, 111, 63, -80, 68, -124, 91, 93, 116, -99, -112, -126, 97, 75, -43, 22, 104, 82, -59, -115, -37, 44, -125, 18, 98, 59, -5, 92, -74, 81, -35, -14, 0, -25, -102, -113, 24, -65, -47, 116, -112, 108, -95, -51, 95, 29, 117, 106, 92, 110, 18, 84, 19, -127, 73, -93, 63, -60, -75, -42, 71, 105, -6, 14, 69, -82, 37, -117, -67, -44, 98, -22, -4, -86, -99, 79, 92, -36, -14, -121, 40, 95, -5, 103, 73, -51, 96, -108, 111, -69, -91, 28, 49, 35, 29, -125, -40, -15, 42, 8, 70, -110, 3, 62, 58, 19, 96, -50, -86, 64, 95, 33, 60, 106, -55, -106, -113, -79, 63, -30, -27, 35, 126, 47, -24, 48, -43, 120, -33, 88, 121, 42, 46, 45, -124, 112, 93, -88, -95, -14, -54, -127, -24, -50, -83, -77, -78, 35, -86, -127, 122, -66, -113, 70, 54, 39, -39, -102, -17, -66, -96, 1, -1, -43, 15, -9, -105, -101, 54, 37, 30, 95, 44, 119, -37, -69, 85, 23, 46, 7, 45, -102, 69, -120, -25, 106, 96, 57, -93, 41, -21, -51, -2, -112, 51, -18, 84, -33, -51, -125, 34, -4, -56, 118, 23, -64, -65, -105, -84, 36, 23, 67, 121, 3, -42, 61, 47, 85, 86, 19, 113, -44, -40, 8, 67, -122, 115, -68, 6, -108, -12, 92, -121, 90, -58, 109, -14, 42, -91, -125, 108, -105, 66, -82, -3, 10, -82, -29, -41, 42, -66, 0, -48, 45, -1, -7, -76, 4, -52, -117, -36, -50, 93, 79, 25, 12, 112, 13, 49, 74, 37, 118, -91, 96, 48, -81, 111, 85, 21, -41, -43, -27, -96, -126, -58, -44, -91, -56, 98, -97, -93, 69, 35, -4, -81, 93, 12, 52, -94, -54, 108, -56, -56, -69, 122, -118, -31, -58, 117, 102, 71, 90, -78, 6, -97, -73, -123, -73, -126, 127, -71, -23, -49, -14, -56, -50, -93, -108, -121, -38, 70, -105, 123, 97, 117, 4, 115, -18, 56, 48, 107, -79, 0, -45, -59, 20, 86, -33, -32, -105, -52, 66, 125, -110, -100, 52, -116, -45, 22, 106, 55, 105, -21, 70, -86, 109, 91, -73, 77, 53, -85, 78, 32, -29, 50, 107, 10, 91, 91, 61, -3, 66, 112, 6, 79, 125, -13, -83, -119, 66, 27, -94, 2, -23, 93, 31, 4, -105, 29, -41, 53, -1, 0, 40, 16, 57, -72, 86, -21, -31, -123, 37, -23, 41, -111, -111, 107, -97, 85, 99, 16, 119, -117, -49, 83, -96, -105, 74, -117, 15, -93, 126, 99, -11, -57, 36, 102, 87, -110, -109, 70, -71, -60, -33, 8, -18, 80, -95, 32, 0, -21, 77, -61, 110, 80, -79, -97, -2, 16, -77, -43, -52, -4, -90, -101, -99, -113, 34, 19, -80, -76, 120, 20, -55, -114, 57, -34, -80, -113, 22, 11, 36, 117, 76, -26, -91, 74, 37, 17, 18, -83, 51, -45, -52, 54, 3, 36, -5, 84, 23, -74, -47, 108, -122, 123, -69, -43, 109, -6, 21, 112, -128, -62, 91, 6, -64, 31, 120, 45, -80, -86, -23, -127, -43, -127, 28, 124, 43, 43, 69, 17, -122, 50, 124, 10, 82, 15, 76, 83, 16, -15, 53, -124, 11, -18, -74, 43, -20, 12, 9, -9, -71, 47, 52, 28, 122, -53, 56, -70, 82, -54, 61, -108, 103, -84, 107, 124, 123, 1, 117, -80, 109, 18, -65, -34, 81, -17, -101, 20, -78, 49, -15, 61, 66, -125, 74, 62, 22, 34, 114, 93, 44, -57, 38, 104, -18, 5, -22, -18, 123, -86, 79, -108, -49, -118, -64, 69, -87, -28, 35, 80, -24, 126, 78, -32, -68, -72, 111, 66, -71, -56, -4, -56, 1, -127, -30, -110, 107, -95, -93, -89, -31, -107, 86, -72, -59, -62, 32, 66, -99, -95, -44, -36, 114, 31, -14, -85, 47, -65, 25, -3, -85, 8, -14, 109, -107, -121, 21, 72, 99, -85, -121, -113, -107, 80, -87, 28, 108, 3, -102, 70, -57, 40, 47, 78, -32, -82, -89, 123, 20, 37, -6, -85, 45, 106, 101, -114, -121, 108, 116, 110, 15, 2, 126, 49, 16, 65, 34, 61, 28, -3, -56, -74, 115, 50, 29, -112, -64, -85, -32, 86, -71, -54, 51, -58, 52, 22, -126, 28, 42, -48, 88, -47, 50, -21, -42, -93, 7, 37, -68, 124, -23, -35, 92, -55, -47, -71, 66, -43, -37, 42, 103, 71, 109, -6, -54, 76, -104, 28, -84, -46, -19, 102, -84, 78, -85, 102, 79, -88, -126, 124, 14, 121, 13, 75, -102, 78, -17, 32, -96, -125, 122, -39, -86, 95, -118, 72, -20, 29, -40, 124, -48, 124, -18, 52, 98, -6, -55, -64, -11, 121, 118, -70, 9, 50, -61, -119, -24, -62, -54, -54, -88, -89, 51, 52, -91, 37, 26, -16, -120, -109, 106, -68, 114, -59, 104, -22, -102, 115, -25, 75, 67, -96, 13, 88, 10, 45, 89, -41, 78, -27, 76, -71, -1, -74, 117, -121, 127, -122, -43, -24, 120, 81, -105, -26, -66, 53, 121, 34, 46, -47, -4, 80, 39, -103, -119, -96, -17, -54, -84, 68, -112, 64, -3, -96, -41, 115, -77, 24, 23, 35, 113, -32, -10, 34, 88, -121, -58, 103, -43, 5, -24, -33, -52, 91, 9, -105, 58, -102, 106, -84, -91, -23, 105, -45, -73, -47, -9, 119, 111, 78, 54, -77, -62, 71, -4, -45, -60, 78, 65, -13, -19, 124, 7, 12, 46, -30, -119, -40, -103, 54, -44, -106, 61, -48, -95, 48, -111, -14, -68, 79, -30, -43, 103, -57, 81, 7, 105, -12, -28, 119, -81, -59, 72, -88, 75, 48, 34, 16, 100, -65, -110, 103, -17, -13, 39, -62, -6, -90, 113, 2, -112, 71, -41, 4, 25, -37, -75, 9, -123, 63, 10, -15, 82, -51, -92, -54, 12, -27, -126, 2, -92, -86, 25, -79, -79, 17, -61, -59, -116, -68, 31, -126, -120, -103, 5, -41, 52, -111, -15, -68, 47, -29, 32, -110, -66, -1, -13, -23, 56, 6, 64, -33, -17, 88, -72, 73, -77, 13, -6, -84, 86, 111, 122, -77, -116, -39, -107, -33, 28, 95, -54, 75, -58, 87, -61, 116, 50, 19, 27, 60, -28, 88, -114, 93, -78, -71, -1, 11, -80, 15, -115, 51, 116, -61, -117, -98, 32, 4, 31, -12, -105, 22, 104, -62, -82, -75, -72, -46, -67, -85, 4, 44, 58, 48, 35, -51, 114, 1, 92, 127, 122, -78, 122, -110, 127, -83, -127, -50, -102, -5, -7, 53, -103, 22, -81, 63, 31, 60, 31, -12, -83, -108, -123, -41, -116, -66, 54, -88, 88, 94, -25, 71, -121, 37, 93, -81, 13, -46, 11, 119, -37, -58, -38, 54, -3, 50, -125, 102, 86, -21, -39, 118, -47, 7, 108, -59, 49, 36, 63, 14, 35, 122, 94, -10, -85, 98, -116, -44, -123, -4, 30, 122, 55, -86, -70, 8, -69, -11, 22, -33, -46, -107, -12, 50, 33, -34, 7, -65, -46, -71, -107, -8, 56, 35, 23, 80, 53, 59, 108, -87, -98, 49, 48, 16, -96, -96, 18, -25, -112, -77, -22, -41, -94, -119, -59, 30, 118, -91, 109, 47, -113, -83, 126, 3, 78, -10, -128, 67, 34, 52, -23, -84, -112, 56, -123, 103, -100, -55, -18, 33, 34, -60, -60, 70, -14, -23, 112, 2, 20, 105, -55, 27, -70, 78, 87, -126, -105, 10, 103, -118, -60, 33, -91, -15, 49, -112, -117, -126, -12, 2, -113, -94, 11, -38, 20, -81, 11, -36, 91, -14, -100, 114, 88, 56, -64, -17, -98, 96, 37, -95, 127, -1, -16, -12, 83, 7, 106, 23, -127, 104, 106, 27, 7, -112, 85, 91, -111, 57, -7, -8, -51, 103, -36, 31, -80, 56, -46, -26, 67, -61, 63, 83, -76, 96, -16, 115, 49, 116, 77, 14, 98, -81, -14, 96, 73, -38, 21, -38, 8, 82, -122, 2, -21, 113, -43, 47, -81, -11, 39, 87, 63, -111, -52, 64, 65, 4, -91, 16, 121, -111, -126, -47, 101, -29, 101, 6, -68, 45, -113, -117, -2, -127, -55, -1, 100, -14, -83, 122, -51, -105, -31, -10, 118, 113, -47, -85, -120, -82, -35, 15, -34, -81, -22, 89, 75, 64, 40, -24, 28, 114, -126, -9, -114, -86, -58, -116, 36, -126, -68, 44, -78, -18, -36, -33, -78, 127, -55, -50, -127, 30, -72, 81, 12, -16, 114, -78, -20, 117, 30, 73, 10, -120, -107, -1, -70, 1, -122, -108, 40, -87, 95, -37, -76, -106, -40, -38, 101, -102, 43, -65, -62, -12, 7, -124, -118, 79, -128, -2, 40, -72, -99, -8, -85, 123, -90, -24, 123, -121, -127, -85, 36, -8, -120, -44, 59, 7, 91, -97, -68, -126, -114, 73, -84, 92, 43, -94, -125, -11, 35, 71, 44, 101, 74, -56, -91, 15, 73, 4, 37, -85, 60, -52, 116, 38, 57, 56, 59, 96, -90, -60, -120, 79, -87, -7, -9, -104, 64, -71, -31, 69, 116, -118, 47, 115, -100, -76, -52, 17, 13, -109, -128, -104, 34, -18, -106, 61, 5, -97, 35, 91, 74, -69, 6, 108, 61, 40, -24, -119, -47, -127, 101, 12, -76, -51, 117, -49, -29, -70, 89, -105, 90, -80, -106, -6, -77, 85, 1, 18, -85, -70, 81, 67, 52, -57, 78, -97, -93, 29, -106, 26, -121, -66, -123, 86, -69, 94, 43, 8, 110, -126, -13, -84, -90, 89, -48, 70, 25, -4, -86, 5, 68, 92, -85, 124, 64, -21, -22, 57, 87, 61, 40, -110, 14, 25, -69, 104, -55, -116, -98, 44, 114, -45, 61, 38, -126, 106, 67, -123, -39, -65, 121, -62, -118, 65, 44, 23, 58, -18, 37, -44, -52, 54, 4, -53, 105, 91, 94, -126, 66, 4, 56, -58, -82, -71, -117, -23, 19, 28, -111, 33, 44, -37, -45, -105, 106, 74, -89, -107, -84, 32, 99, -66, 120, 118, -51, 101, -27, 22, -62, -28, -56, -71, 74, -116, 64, -31, 14, -5, 6, -99, 75, -80, 38, 9, 24, 13, 103, 107, -128, 16, -97, -8, -94, 67, -103, -86, -103, -76, 39, 24, -65, -119, -22, 97, -22, -119, 67, -123, -43, 119, 126, -80, -49, -118, -95, 21, -114, -90, -72, 97, -11, 49, 81, 38, -126, -124, 71, 39, -92, 81, 4, 109, 34, -94, -67, -12, 4, 79, 120, 36, -30, 113, 71, -114, 22, -30, -109, -118, -60, -70, 106, -34, 42, 19, 123, 7, 7, 7, 71, -26, -55, -47, -62, 26, -62, -74, 126, -26, -92, -18, -48, -90, 3, -93, -84, 12, -42, 123, -42, 75, 103, -3, 20, 127, 108, 32, -28, 119, -6, -15, 25, -27, -18, 99, -28, 68, -45, 61, 48, 19, -39, 103, 49, 4, -124, 89, 106, 68, -30, -126, -34, -113, -72, -47, 7, -3, 108, 32, -55, 63, 68, -106, 33, 57, -126, -107, 68, -84, -26, -28, -51, 39, 53, 81, 51, -14, 109, -89, -91, -12, 65, -38, 124, -43, 126, 119, 0, 32, -26, -16, 122, 127, -81, 126, -110, 11, -11, -80, 69, -60, 65, -40, 43, -50, -65, 72, 22, -43, -12, 39, -121, 70, -22, 114, 102, -87, 44, -1, -108, -50, 64, -48, -107, -92, 3, -105, 84, 27, -87, -54, 66, 66, 3, 0, 123, 17, 124, -90, -18, -66, 102, 60, 65, 93, -31, 84, -43, 5, -113, -44, 2, -119, -119, -29, 81, -11, -44, 107, 38, 24, 91, -30, 123, 31, 90, 36, -128, -94, -58, 42, -13, 79, 33, 61, 6, 81, 56, -105, -31, -24, -4, -110, 118, -31, -105, 9, 41, 34, -73, 78, 104, 45, 107, -7, 60, -12, 12, -67, -28, -123, -56, 42, 107, -86, 51, 109, -56, 12, -82, 110, 35, 45, -128, -37, 103, -90, 86, 27, -3, -93, -103, 105, -30, -81, 101, -64, 82, 66, 65, -14, -33, 3, 8, -64, 60, -82, 70, 75, -51, -109, -117, -14, 34, 90, -100, -14, 124, -64, -113, 39, -13, -1, 45, 94, -72, 22, 3, 10, 10, 97, -60, -124, 49, -59, 123, 92, 100, 106, 19, -10, -30, -99, 87, 121, 105, 62, -60, 106, -2, 110, -113, -51, 86, 9, -75, 102, -103, 67, 71, -56, 41, -84, -30, 94, 107, -28, 14, -75, -41, -3, -9, 63, -54, -111, -67, -73, 44, -64, -67, 124, 16, -66, -59, -89, 32, 99, 66, 127, 107, -1, -113, 95, -88, -88, -4, 38, 97, 62, 114, -115, 80, 26, -38, 29, -42, -17, -71, 88, 50, -86, -1, -31, -99, -28, 88, -76, -54, -118, -76, 20, -40, 92, -107, 1, -14, 39, -120, -104, -120, 76, -68, 62, -117, -120, 103, 122, 30, 106, 43, -96, -55, 57, -101, 87, -39, 57, -111, -115, 46, -17, 101, -127, -62, -100, -64, -9, 10, -103, -86, -60, -38, -17, -100, 85, -126, 52, -75, 46, -101, -31, 77, -79, 13, 85, 15, -51, 16, -89, -1, 26, 29, 91, -107, 22, 110, 7, -53, 56, 28, -56, 113, 97, 0, 58, -91, -104, 24, -72, -23, -81, -45, -93, -13, 119, 47, -65, -36, 53, 96, 50, 11, 35, -17, -17, -70, 124, 103, -78, 84, 126, 5, 123, 4, -93, 119, -67, 47, -19, -33, 97, -82, -81, 96, -15, 93, -127, -6, -1, 33, -79, 114, 23, 102, 8, 30, -11, 127, -59, 1, -4, -18, -85, 55, 99, 123, -18, -36, -119, -74, 4, 80, -16, -109, -30, 116, -114, -121, -91, -34, -90, -43, -62, -114, 116, 5, 8, -83, 124, 2, 73, 80, 60, -27, -58, -20, 31, 35, -46, 15, 59, -84, 59, 5, -1, -37, 58, -47, -108, -81, -99, 62, -95, -57, -2, 59, 17, 58, -21, -72, -119, -88, 0, -33, 31, -87, -80, -39, 43, -21, -69, 108, 89, -121, 118, -96, -96, -46, -34, -52, -123, -104, -24, -1, -93, -29, 2, 16, -47, -113, 106, -33, 15, 104, 26, 18, -124, -31, -95, 122, 111, 10, -54, 42, 35, -63, 75, -5, -77, 19, -63, -17, -113, -124, 52, 12, -81, -57, 30, -117, -84, 115, -40, -33, 76, -1, -46, -72, -104, -114, -90, 2, 26, 18, -90, -9, -123, 94, -6, 70, 16, 37, -65, -47, 126, 66, 113, -54, 83, -80, -23, 87, 64, -27, 115, -56, 72, -123, 107, 36, 121, 18, 116, -57, -16, 25, -38, 104, 6, 45, 10, -25, 97, 82, -114, -109, -37, -46, -49, 115, -103, -2, -29, 112, -96, -112, 20, 0, -98, 18, 74, 4, -40, -33, -4, -30, -115, 11, 70, -4, 29, -7, 127, 75, -38, -80, -101, -121, -53, 96, 61, -24, 84, -68, 94, 100, 72, 112, -66, -5, 76, 87, 1, 100, 30, -89, 98, 70, -114, 11, -66, -70, 101, 40, 10, -57, 89, 77, -113, -91, -119, -8, -106, 91, 66, 104, -35, -75, -100, -101, -22, -65, -120, 26, 24, 29, -47, -104, -102, -54, 17, 6, -122, 65, 107, -1, -52, -17, 86, -78, -101, 125, 1, -106, -90, -94, 23, 45, 33, -55, -21, 84, -107, -46, -114, 66, 92, 49, -14, 23, 108, 114, 90, -90, 32, -48, 14, -101, 56, -30, 53, -3, 36, 99, 76, -76, -73, -27, 103, 57, 36, 116, 73, -43, 68, 97, -30, -125, 125, 81, 28, -21, 124, -3, -27, -126, -90, -125, -58, -10, 111, -59, 77, 117, -52, 8, -25, -23, 123, 29, 62, 10, -52, 43, 0, 65, -75, 116, -101, 117, 112, -59, 1, 53, 17, -84, 72, -31, 22, -70, 124, -19, 5, -82, 69, -28, -33, 127, 8, 89, 108, -15, 19, -57, 57, -77, 12, -102, 70, 99, -86, -85, -78, -96, 68, -124, 38, 85, 71, 55, -47, -7, -48, 84, 104, -103, -78, 55, -97, 52, 68, -28, 73, -59, -122, -113, -90, 47, -107, -46, 5, 44, 47, 45, -45, 40, -6, 58, 27, 90, -101, -79, 117, -6, -107, -42, 47, 35, -69, -20, 30, -38, 59, 30, 19, 35, -21, -19, 42, -97, -33, 107, 112, 111, -97, 61, -104, 40, 13, 43, -128, 20, 89, 108, -126, 71, 71, 90, -76, 40, 26, 82, -95, -25, -11, 45, 79, 109, 66, 10, -13, -96, 25, 13, -48, 80, -9, 12, -5, 35, -18, 110, 35, -6, -42, 42, 27, -11, -105, -37, 69, -63, 58, 30, -113, -47, 118, 46, -2, 15, -127, -54, 23, 3, -12, -90, -76, 121, 38, -17, -29, -13, -128, 70, -100, 10, 105, -64, -48, 28, 78, -5, 4, -73, -85, -54, -40, 64, -126, 109, 122, 121, 55, 7, 99, -16, -71, -5, -34, 74, -74, -20, -111, 22, 95, 60, -65, 111, 24, 51, -8, -111, -75, 13, 42, 74, -63, -87, -95, 39, 106, -63, 1, 56, -55, 5, 39, 52, -116, -14, -59, 123, 75, -85, 19, -76, -20, -45, 19, -6, -92, 91, -20, -11, -9, -19, 54, 26, 20, 118, 81, -44, -17, 116, 24, -57, 125, 11, 108, -75, 54, -105, -122, 118, 56, 94, -6, -24, 54, -16, -77, -79, 87, 21, 33, -110, -30, -124, -113, 115, 2, -45, 122, -97, 71, -67, 40, 74, 2, 121, 12, -46, -24, 54, 7, 57, -3, -3, -125, -128, -77, -52, -111, -108, -34, -127, 112, -107, -26, 78, -75, 13, 4, -121, -10, -119, 43, 11, -64, -6, -31, 106, -126, -89, -88, -117, 69, -45, -53, 29, 53, 46, -81, -3, -12, 31, -60, -98, 27, -23, -21, 30, -85, -11, -81, -13, 37, 27, -6, -121, -42, -63, -65, 125, -64, 18, 66, 69, 3, -108, 28, 49, -108, 83, -98, -22, -103, -55, 79, -8, 124, -125, -110, -52, 23, 85, -69, 30, 69, -78, 109, -34, -83, 1, 72, -51, 34, 94, -58, -41, 32, 14, -101, 10, -97, -75, 81, -56, -93, 65, -2, 76, -33, -122, -55, 45, 90, -95, 11, -31, -20, -104, 94, -55, 46, -36, -18, 76, 30, -112, -69, -55, -112, -40, -95, -62, 71, -89, 97, -68, 61, -124, -57, -11, 123, 101, -94, 88, 32, 25, 127, -107, -42, -41, -107, 27, -85, -107, 124, 43, 82, -34, -112, 58, 78, -59, -40, -108, 126, -107, 84, -89, -19, -23, 54, 98, 82, 117, 91, 94, -106, -87, -125, -35, -44, -24, 105, 116, 40, -24, -38, 21, -83, 60, 85, -44, -91, -127, -116, 72, -22, 88, -23, 54, -93, -2, -120, -101, -126, -2, 16, -43, -92, 97, -22, 64, -69, 12, 21, 62, 14, 68, -1, -100, -2, 77, -15, 85, 38, 119, 83, 6, 117, -54, -1, 126, 47, -100, 32, -40, 67, -70, -101, 103, -2, -12, -16, 70, 120, -52, -22, -21, -10, 10, 99, -19, -15, -112, -53, 64, -30, 43, -67, 59, 16, -20, 122, -90, -21, -42, -86, -62, -37, -37, -51, -63, -4, -96, -99, -27, 32, -24, -107, -24, -70, 107, -41, 72, 35, -33, 84, -94, 58, -21, 113, 78, 37, -9, 63, 115, -37, 39, -100, 33, 25, -31, -87, -2, -89, 119, -8, -30, -50, -4, 37, -13, -10, -53, -107, 33, 51, -91, 29, -124, 76, -91, 17, 101, -9, 67, 110, 103, -120, 5, -57, -46, 89, -22, 65, 108, 37, 19, -21, 10, 120, 84, -34, -11, 118, -59, -23, -97, -81, -91, -18, 93, -19, -33, -3, -20, -68, -18, 0, -53, 127, 46, 9, -88, -70, 110, 26, -19, -62, -44, 116, -24, 113, -18, 108, 42, -79, 126, 109, 95, 127, -3, 16, -63, 104, 19, 9, -77, 93, 83, -116, 8, 10, -38, 6, 54, -12, 93, -28, -37, -38, 50, -69, -9, -91, 53, -37, -98, -101, -44, -77, -86, 48, 41, -114, 42, -14, 10, -59, 121, 52, -26, 74, 102, -86, -24, 30, -59, -49, 31, -119, 110, -19, -115, 91, 68, 94, 59, 106, -115, -53, -45, 116, 127, 85, -118, -128, -120, 54, 115, -44, 47, -34, 30, -20, 15, 40, 17, -60, 99, 71, 118, -21, 35, 98, -85, 31, 88, 5, -26, 44, -32, 67, -96, 85, -124, 54, 1, -101, 29, 56, -66, -51, -88, -106, 34, 24, -123, -18, 54, 57, -94, 73, 71, 82, -80, -49, 92, 51, -8, 79, -17, 12, 95, -35, 6, -56, -36, -81, -87, -29, 49, -40, 70, 114, 73, 62, -101, -73, -28, 104, 89, 125, -11, 52, -19, 13, 41, 74, -21, -53, -126, 22, 91, -81, 63, -29, 65, 124, -105, 4, 95, -79, 69, -22, -97, 22, 20, 83, -26, -104, -100, -48, -20, -59, -110, -89, 123, -67, 62, -64, -16, -46, 36, 18, -117, 36, -60, -96, 3, 41, -50, 109, -18, -74, 18, -71, 16, -127, -108, -84, -57, -87, 127, 111, 32, -101, 39, -89, -64, -89, 63, 4, -47, -99, -21, -127, 23, -111, 38, 22, -2, 5, 32, -30, 81, -99, -113, -75, -117, 111, 69, -21, -25, 18, 98, 5, 110, 24, -39, -70, -24, 123, 51, 53, 28, -21, -50, -101, 65, 105, -71, 14, 56, -113, 81, 17, 10, -62, -8, -69, -82, 104, -124, -5, -87, -112, -22, 58, -86, -124, 125, 9, -13, 96, -103, 83, 6, -54, 68, 16, 89, -30, -64, -123, -4, -64, -78, -7, 31, 77, -80, 53, -70, -4, -123, 87, 110, -50, 30, 30, 86, -44, 2, 31, -21, -45, -82, -38, -35, -94, -10, 71, -51, -112, -36, 67, 77, 58, 87, 27, 79, 49, -90, 124, 125, -66, 53, 35, -101, 34, -83, -3, -102, -111, -38, 94, 121, 54, -18, -120, -10, 39, -59, -7, -114, -81, 28, 62, 60, 46, -24, 0, -115, 20, -23, 49, -101, -38, -6, -78, -29, -26, -15, -14, 39, 104, 108, 92, -43, 82, 78, 91, 83, 17, -122, -90, 64, -58, -114, 94, 63, 59, 21, -117, 59, 125, 101, 115, 48, -68, 67, 101, 103, 58, -35, 124, -31, -49, 56, 79, -87, 72, 104, 105, -96, -56, -4, -4, 93, -70, 103, 125, 0, 30, -113, 15, 70, 23, 97, 5, -83, -69, 61, -13, 81, 63, 39, 51, 14, -72, 76, 70, -86, 117, 49, 121, -69, -77, -79, 96, -119, 16, 49, -39, -18, 105, -68, -5, -43, 91, 83, 65, -123, -114, -107, -9, -69, 76, -105, 65, 109, 102, -20, 29, 61, -7, 21, -30, -90, 44, 82, -12, 88, 85, -73, -97, 34, 98, 15, 97, -29, -116, -107, -82, 115, -9, 21, -80, -5, 37, -21, 54, 31, -52, -10, -80, 19, 64, -20, 75, 98, 99, -97, 73, 3, -35, -114, 5, -50, -17, -120, -28, -102, 83, -13, -22, 12, -54, 94, -55, -7, -91, 42, -72, -61, 11, -18, -21, -79, -7, 1, 66, -79, 114, 122, -75, -85, -71, 48, 15, -30, 23, -45, 12, -80, -6, -120, -100, -63, -28, 24, 7, 63, -79, 89, 26, -25, 92, -109, -7, -109, -70, 53, -20, 89, 23, 96, 2, -96, 92, 21, 60, 95, 72, 113, 12, -63, 109, -67, -113, -81, 85, -74, 65, 59, -50, -112, 103, -110, -93, -92, 119, -69, -78, -54, 81, 67, -122, 87, -21, -81, -17, -105, 76, -96, 126, -16, -80, -47, -9, -53, -81, 72, -61, -55, 36, -51, 74, -27, -105, 86, -54, 23, 83, -44, -66, 16, 20, -118, -48, 120, 82, 113, 124, 23, 9, 97, -120, 60, -14, -122, -23, -40, -114, -22, 40, -114, -1, -110, 76, -41, -123, 109, -63, -46, -51, -7, 88, 84, 39, -1, -68, -16, 14, 121, -18, 68, 76, -10, -17, -115, 86, -98, -75, 52, 82, 49, 29, 22, -119, -3, -77, 28, 72, -101, -95, -1, -98, -121, -106, -17, -65, 45, 106, 41, 44, -52, 0, 34, 6, 91, -123, -47, -16, -37, -57, 71, 53, -57, -85, -123, 127, 97, -67, -24, -20, 121, -1, 44, -90, -105, -32, 73, -117, 88, 76, -30, 32, -88, 42, -23, -111, 23, -15, -60, 117, 45, 23, -28, 40, 106, 107, 125, -69, 25, -116, -108, 79, 89, 39, 103, 84, 103, -27, 79, 27, 106, 101, -99, -23, -85, 25, 108, -8, -5, -55, 0, -98, 71, 89, -6, 71, -5, 111, -54, -107, 0, -110, 113, -34, 65, 12, -95, 112, -47, -119, -52, 22, 30, -75, 122, 9, -121, -26, -48, 109, -73, -88, 44, -100, -103, -79, 117, 14, -104, 127, 88, 9, -72, 18, -110, 104, -92, -25, 8, 47, -36, 118, 28, -124, 61, 59, -33, 49, -47, -25, -26, -26, 27, -19, 122, -65, -49, -108, -90, -54, -34, 88, 1, -78, -123, -74, -95, -36, 7, -40, -99, 110, -63, 81, 20, 51, 37, 13, 100, -11, 119, -67, 118, -45, -57, 108, -89, -7, -52, -44, -65, 110, -48, -108, 111, -39, -78, -77, 11, -1, 36, 16, -127, 88, -87, 84, -43, -23, 23, -100, -29, -6, -22, 120, 71, 97, -126, -7, -123, 75, -108, -121, 107, 90, 46, -84, 7, 127, 105, 55, -9, -15, -43, -106, -75, 98, -107, 123, -47, 93, 72, 47, -109, 104, -96, 37, -9, 103, -76, 41, -115, -22, -50, 117, 21, 43, -87, 18, 127, 5, -126, -50, 1, 6, -43, -113, -69, -118, 69, -96, -98, 77, 25, -43, 38, -87, 23, 48, -126, -33, -112, 91, -64, 33, 98, -128, -128, -98, -7, 70, -107, -37, 44, -49, -127, 37, -106, 19, -47, -58, -120, 103, 125, -30, 92, 37, 14, 88, 37, -11, 103, -30, 53, -26, 113, -50, -56, -3, -125, 81, 79, -94, 85, 10, 13, 82, -110, -19, 116, -67, 61, -62, -118, -107, 63, -127, -85, 33, -71, 4, -58, 88, -102, 60, -7, 85, 104, 44, -50, 42, -94, -51, -94, -40, -97, 42, 69, 5, 45, 32, -59, 63, -128, 36, 1, 89, 30, -85, -81, -57, -93, -123, -48, -28, -6, -2, -94, 4, 84, 0, 26, -60, 118, -121, 76, -113, 8, -4, 123, -81, -55, 22, 41, 34, 1, 75, -2, 27, 56, -36, -11, 62, -9, -41, 34, 127, -74, 91, 86, 32, 82, 118, 48, 125, -30, 18, 91, 93, -96, -103, -11, -101, 1, 97, 23, 73, -118, -99, 122, -8, -28, -63, -26, -62, -9, 121, -25, -117, 46, -114, 8, 112, -95, 38, 35, 36, 6, 100, 77, -16, 107, -54, -44, -16, 28, -14, -10, 81, 86, 71, 116, 125, 105, -83, 76, 50, -10, 51, -50, 48, -91, -40, -12, 4, 113, 114, 78, 111, 19, 37, 57, 50, -43, 105, 88, 95, 118, -94, 107, 126, -7, -29, 35, -86, -9, 51, 126, 113, -69, 94, 62, 34, -74, 117, -70, -66, 57, -3, -120, 67, -42, -31, -48, 40, -22, 20, 21, -34, -124, 23, -16, 124, 69, 117, 62, 35, -94, 89, 29, 78, 67, -1, 78, -13, -124, -103, 98, 119, 61, 41, -103, 38, 11, 2, -37, 24, 118, -38, 12, -66, -92, -41, 73, -109, -25, 58, 38, -26, 77, -12, 66, -87, 109, -39, -16, 18, -41, -62, -107, 84, -66, 87, 4, 19, 106, 82, 58, -34, -3, -2, -49, -87, -125, 19, -12, 109, 28, -39, 29, -56, -50, 46, 84, -5, -31, 125, -24, -102, 109, -117, 40, -84, -19, 110, 64, 120, 55, -41, -17, -62, 101, -56, -103, -128, 6, -43, -104, 36, -26, 4, 5, -41, 64, 11, 108, -14, -93, -65, 17, -95, 11, 108, 55, 76, 34, -64, 28, 110, -11, -44, 126, -97, -27, 78, 75, 106, -41, 57, 16, 56, 17, -20, -3, 107, -115, 113, 69, -56, 30, 123, 101, -24, 127, -97, 28, -73, 117, -27, -41, -106, 35, -24, -20, -63, -128, -30, 99, -95, -26, 120, -113, -3, -23, -94, 69, -128, -29, 126, 33, -110, -19, -122, -79, -55, -57, -66, -84, -81, 54, -33, -52, 117, -86, -99, -113, 55, -71, -73, -77, -35, -128, 88, 69, 111, -121, 11, -36, -49, -75, 16, 92, -95, 73, -90, 39, 86, 2, 38, 106, -19, 122, 13, 73, 48, -1, 117, -111, 77, -42, -78, 116, -55, 11, 66, -62, -61, 44, 63, 106, -12, 70, 32, -64, 65, -121, -65, -113, -127, -115, 26, -15, -46, 46, 66, -22, -4, 45, 1, 74, 26, 13, -106, 83, -64, -104, 104, -57, 84, -72, 27, 38, 114, 117, 35, 41, 104, -68, -74, -107, -76, 50, 107, -53, 69, 25, -12, 78, -8, 112, -126, 24, -75, 33, 76, 90, -124, 72, 99, -119, 44, -76, 77, -13, 107, 42, 122, -122, 39, 16, -29, 82, 39, -8, 76, 15, -76, -35, 77, -85, -37, 119, -47, 20, -19, 2, 68, 125, -23, 78, -121, 104, 64, 62, 70, 124, -29, 43, -49, 125, 34, 4, 96, -18, -70, -64, -33, -28, 69, -70, -77, -5, 35, 123, 79, -90, -42, 119, 32, 104, -46, 101, 85, -61, -115, -126, -64, -7, 123, -47, -74, 50, -109, -96, 25, -95, 42, 77, -86, -13, -50, 23, -82, 60, 101, 54, -8, 28, 45, -97, 110, 32, 105, 125, 62, 26, -108, -57, -76, -122, -107, 114, -6, 59, -28, 11, 19, -70, -117, 86, 104, -19, 19, 23, 90, -108, -41, -4, 109, 116, -45, 35, 89, -45, -54, -21, -51, -89, -121, -10, 13, -76, 32, 124, -109, 25, 70, 73, 32, 47, 62, -122, 16, -40, -98, 105, -97, -118, 110, 103, -9, 110, -71, 117, -101, -37, 96, 50, -67, -49, 55, -111, 109, -8, -79, 72, -30, 117, 116, 77, -100, 79, -122, 16, -68, 28, 74, 33, 52, -94, 117, 10, 30, -76, -73, 106, 125, 46, 119, -37, -103, -45, -89, 97, 112, 112, 0, 28, 9, 55, 101, -74, -40, -55, 51, -86, 13, -15, 106, -122, -37, 12, -90, -57, 80, -10, 112, -9, 5, -107, 121, 72, -47, 11, -97, 69, 75, -41, -27, 122, 60, 15, -96, 58, -23, 127, 103, 111, -19, -46, -36, 99, -67, -75, 60, 94, 85, 27, -117, 119, -60, -14, 64, -101, 78, 116, 11, -6, -38, 58, -20, 56, -17, 59, -16, 20, 65, -39, 22, 11, -47, 10, 41, -124, -43, -15, 50, -127, 31, 101, -95, 64, -117, -108, -90, 7, 117, 114, -77, -33, -29, 7, 99, 60, -26, -121, 71, -119, 54, -28, -82, -26, 77, -120, -24, -19, 125, 49, -120, -1, -82, 61, 101, -47, 24, -94, -20, -27, 109, 64, -11, -33, 32, -60, -50, 90, -93, -125, -104, -123, -3, 101, 40, 87, 42, -41, 53, 45, 57, -15, 86, -97, 47, 121, 96, 8, 0, 91, 11, -67, -23, -100, 87, -110, -1, -128, 58, -65, -120, 23, 35, -43, -82, -20, 7, -40, 14, 30, -118, 72, 119, -128, 64, 92, 45, 105, -38, -120, 118, 31, -9, 106, -85, -81, 22, 46, -18, -98, 52, 74, 43, -112, -28, 103, -86, -40, 10, -9, 2, 74, 124, 48, 81, 101, -84, -100, -37, 120, -34, 87, -13, -47, 54, -50, 52, -5, -58, 90, -74, -61, 72, 112, 74, -121, 75, 6, -119, 81, -74, -120, -43, 95, -20, -83, 22, 29, 101, 26, -106, -19, 97, 51, -11, -38, -33, 69, -5, -36, -91, 122, -29, 29, 36, 4, 87, -97, -46, -16, -8, 17, 9, 125, 11, -57, 47, -126, 32, -91, -71, -1, -61, 101, 15, 106, -88, 51, 66, -15, -87, -74, -110, -81, 95, 26, -34, 9, 53, 1, -35, -110, 30, 92, -38, -46, -11, 85, -29, -128, 74, 15, 105, -32, 60, 50, 21, -8, -128, -1, 74, -101, -36, 0, -4, 51, 84, 75, 4, 9, 45, 23, -51, 99, 6, 68, 77, -23, -24, 80, -102, -125, -26, 10, -127, 56, 102, -111, 5, 70, 35, -55, -82, 47, -1, -124, -44, -127, 53, -128, -73, -22, -67, 76, 126, 27, -72, 115, 41, 47, 101, 84, 98, -21, -2, 4, 64, 5, -22, -2, 37, 89, 33, -37, 120, -97, 64, 116, -30, -128, -53, -120, 104, 73, -94, 80, 30, 45, 29, -38, -54, 15, 84, 22, -20, 116, 43, -57, -68, -22, -48, -76, 107, -21, 112, 98, -71, 111, -28, -104, 61, -75, -87, 94, -105, -103, -26, -34, 80, -118, 127, -18, -16, -24, 108, 21, -9, -122, -82, 46, -98, 109, 47, -39, -124, 46, 97, -65, -68, -8, -74, 32, 91, 54, 23, -18, -50, -112, -20, -63, 69, -84, -35, -65, 19, -51, -104, 113, 115, -98, -21, -122, 37, -46, 57, 42, 51, -81, 38, -8, 46, -33, -96, 31, -8, -92, -107, 31, 51, 26, -54, -59, -49, -17, 101, -30, -62, -120, 118, -17, 34, 127, -31, 9, -35, -23, -118, -48, 54, 59, -43, -59, 43, 56, 70, 28, -79, -43, 78, -98, 108, -19, -108, 75, 117, -120, -100, -101, -102, 64, -18, 122, -43, 66, -66, 81, -110, -37, 88, 83, 19, 2, 57, 87, 34, 12, 56, 47, 28, 12, 2, 21, -23, -66, 42, -89, 64, 91, -126, 99, -106, 77, -85, 28, -74, -42, -28, -87, -35, -9, 60, -28, -45, 84, 95, -28, 35, 40, -97, 114, -2, 50, 33, 86, 96, 123, -43, 123, 100, 69, -78, 23, 39, 6, -100, -53, -62, -34, -23, 81, -48, -82, 49, 82, 40, -69, -74, 94, 42, 107, 24, -60, -49, 105, -51, 21, -8, -21, -70, 82, 121, 53, 29, 0, 12, 122, -10, -68, -8, 67, 119, 26, 119, 87, -119, 110, -83, -128, 85, 40, -10, -26, -105, -1, -82, -74, 42, 80, 81, 35, -83, -8, 15, 60, -13, 61, 28, 51, -23, 16, 38, 22, 6, 99, -12, -66, 102, -13, -124, 126, -94, 75, -63, 127, 86, -120, -120, -55, -95, 27, -44, -66, 96, 17, -29, -43, 40, -73, 70, -105, -57, 111, 123, -57, -48, 117, 87, -27, -52, 69, 18, 114, 54, -116, 36, 96, 74, -97, -99, -128, 28, -79, 5, -40, -35, -6, -40, 103, 67, 16, -104, -45, -5, -40, 16, -32, -90, 124, 7, -117, -120, -83, -29, 69, -2, 19, 39, 40, -70, -31, 17, -15, -38, -75, 117, -103, 80, 84, 93, 22, 62, -81, -24, 40, 16, 100, 64, 84, -74, 36, -72, -65, 18, 29, 68, -66, 13, 117, 78, 18, 90, 25, 23, -77, -31, 55, 83, -71, 21, 121, 2, -65, -16, -127, -100, -49, -70, -108, 50, -16, -82, -8, 89, -65, 94, -30, 47, 117, -120, 78, 94, 110, -66, 73, 90, 63, 58, 100, 119, -46, 101, 94, 9, 100, 37, -100, -121, -58, 33, -47, 59, 89, 110, -113, 24, -97, -11, -30, 90, -3, -61, 96, -36, -65, 34, -72, 9, -66, -75, 25, -87, 121, 27, -13, 4, -28, 58, 89, 20, -77, 4, -16, -62, -27, 105, -66, -90, 114, 48, 10, 108, 17, -77, -86, -55, -114, 54, -120, -70, -39, -46, -95, 69, 103, 11, 41, -91, 97, -120, -109, -103, 70, 103, -6, 1, 63, -26, -123, -42, 48, -20, -30, -97, 98, 99, 53, 71, 98, -48, -59, 22, 111, -26, 15, 41, -22, -44, -25, 75, -109, 42, 8, 57, -78, 115, 59, -47, -120, -87, 16, 58, -85, 6, 82, -81, -20, 2, -104, 123, -3, 89, 56, -65, 90, -8, -44, -50, 59, 31, 74, -96, -10, 109, -43, -66, 96, 99, -101, 46, 43, 46, -56, -117, 0, 89, 42, 101, 35, -83, -52, -13, -73, 75, -116, -9, 84, 108, 66, 121, 127, 5, 90, -34, 125, 124, -111, 38, 105, -59, -95, -81, -121, 42, -98, 59, 102, -102, 66, 72, 116, -94, -57, 21, -53, 78, -29, 114, 76, 55, 33, 7, -4, -127, 95, 126, -52, -32, -1, 45, -51, -36, -126, -118, -27, 112, 107, -77, 71, 64, 43, 40, -74, 8, -20, -5, 98, 5, 13, -110, -38, 13, -41, -96, -63, 18, -61, -64, -27, -88, 3, 45, 80, 107, 22, -76, -2, 102, -76, 86, -58, -63, 111, -11, 120, -36, 77, -30, 46, -107, 35, 119, -36, -36, 54, 63, -93, 29, 125, 18, -50, -95, -39, -98, 68, 75, 86, -113, 52, 115, 124, -118, 69, 31, -10, -89, -8, -90, -30, -70, 121, -46, 107, 20, 46, -18, 54, 110, 12, 14, 66, -92, 113, -77, 121, 56, -66, -99, -21, 66, 120, 78, -41, 109, 28, -78, -121, 102, 90, 94, 11, 103, -21, 109, -110, -109, 124, 55, 105, 29, -128, 33, 17, 46, -121, 48, 79, 68, -105, 60, 118, -1, -22, -6, -108, -100, 2, -35, -73, -93, 55, -49, 124, -85, -11, 123, -47, -83, 78, 15, 50, -69, -94, 124, -100, 47, -87, 35, 83, 0, 79, 11, -19, -84, -61, -91, -68, 17, -98, -125, -102, -123, 64, 6, -84, -97, -11, 36, -46, -57, -39, 72, 112, 16, 118, 120, -100, 114, -82, 58, 32, 48, -78, 119, -51, -43, 72, -123, -103, -10, 44, -105, 83, -84, -74, -51, 97, 64, -115, 22, 109, 53, 17, 78, 97, -66, 69, -46, -94, -61, 9, 39, 123, -64, -70, -110, -69, 61, 95, -79, 20, 5, 28, 0, 79, 49, 18, 9, -128, 69, 101, 127, -29, -37, -95, -50, 20, -65, -65, -43, -84, 31, -9, -52, -87, -6, 54, 99, 1, 25, 113, -112, -72, 87, 5, -42, -4, -52, 20, 7, -124, 2, 9, -9, -47, -73, 84, -85, 112, -110, -61, -83, -4, 65, 100, 62, 87, -46, -107, 72, 56, -28, 32, -53, 31, 90, -86, -9, 75, -95, 31, -70, -14, -27, 81, 54, -21, -126, 84, 85, -27, -112, -117, -3, 58, 25, 39, 113, 16, -47, -78, 30, 56, 39, 39, 93, 93, -29, 118, 67, -115, 60, 54, -103, -118, 84, -33, -21, 67, -92, -86, 71, -108, -16, 89, -97, -27, -67, 25, 14, 85, -31, -26, -36, -115, 21, -102, 77, -90, 65, -112, 54, -123, 62, 80, 51, 98, 123, 78, -38, -38, 37, -102, -79, -60, -51, 37, -16, -8, 30, 76, -110, -91, -73, 45, 75, 120, -21, 6, 2, 23, -44, 124, -16, -54, -110, -125, 101, 3, 88, 64, 9, 87, 76, 9, 62, -12, -88, -48, 121, -88, -114, -30, 104, -15, -17, 34, -35, -7, -4, -109, -95, 44, -9, -35, -24, -64, 65, 3, -109, 58, -118, 97, 42, 78, -27, -24, 33, 15, -59, 42, 12, -76, -37, -14, -99, 86, -107, 74, -96, 51, -125, 63, -73, 72, 38, 5, -44, 102, 35, 24, 7, 75, 67, 109, -98, -61, -116, 64, 122, -69, 103, 58, 31, -56, -26, -25, -76, -39, -56, -21, 116, 67, -55, -94, 56, -48, 90, 125, 81, -82, -122, -46, -89, -3, -121, -22, 14, -114, -40, 28, -23, -103, 79, -128, 70, -83, 30, -19, 108, -5, 60, 37, -69, -124, -13, 100, 22, 67, 126, -98, 3, 66, 120, 11, -112, 54, 101, -85, 2, -111, -114, -84, -51, -78, -15, 41, 19, 60, -107, -8, 19, 7, -89, 79, 23, 121, 121, 84, 66, -51, 26, 71, 35, -67, -3, 18, 114, -72, 100, -70, -44, -64, -20, -30, -19, 50, -104, -39, 117, -9, 12, 48, -11, 100, 126, -66, 31, 24, -28, -113, -62, -26, -124, -119, 9, 60, -14, 15, -73, 51, -126, 82, -17, -118, -39, 4, -125, 81, 71, -62, 12, 61, 49, -27, 15, 77, 25, -44, 49, 121, -12, -58, 95, -48, -53, -99, 38, -58, 115, -95, -93, 31, -115, -6, 43, -71, -103, 71, 60, 24, 126, 39, 10, 91, -70, 58, -77, 120, 65, 45, -75, 40, -48, 62, -81, 99, 66, 36, 85, 62, 122, 126, 5, -41, -21, 78, 119, -87, -72, 18, 101, -112, -5, 77, -96, 57, -24, -111, -78, -128, -63, -97, 98, 82, -63, 45, 111, -70, 49, -26, 28, 3, 20, 72, -25, -109, -23, -20, 83, -122, 25, -7, 23, -79, -34, 40, 13, 43, -35, -113, 32, 25, -127, 50, 87, -112, -41, -14, -92, -101, -101, 24, -58, 117, 79, -69, 58, -49, 103, 73, 86, -48, -73, -95, -26, 115, 3, 51, -127, -16, 14, 99, -7, 57, -8, 11, 5, -23, -4, -106, 33, -3, -117, 125, 81, 53, -63, -11, -81, 63, 53, -92, 112, -82, 121, 63, -81, 92, 84, 49, -97, -35, -47, 110, -99, 92, 22, -19, 7, 21, 104, -120, -16, 126, 84, -114, -73, -120, 106, 92, 83, 4, -63, -24, -17, -123, 108, 31, 50, 55, -19, -94, 17, 79, 31, 7, -92, 118, -15, -62, 107, -7, 18, 74, 120, 98, -54, 94, 91, 90, 30, -16, 87, -30, 117, -56, -49, 39, 73, 94, -128, 52, 19, -24, 34, -63, 6, 10, -48, -101, -114, 29, -18, -59, 49, -67, -47, -10, 44, 101, 35, -6, -75, -49, -125, -34, -75, 65, -35, 54, 120, -81, -110, -9, -30, 31, -8, -124, 95, 74, 61, -42, 123, -8, -103, 57, 113, 112, 10, -94, 69, 73, -43, 1, -31, 109, 38, 24, 33, -37, -37, 79, -37, 8, -22, -11, 75, -17, 34, -44, -79, -111, 107, 95, -122, -65, 114, 35, -64, -16, 83, -98, -61, -42, -3, -95, -87, 105, 37, 31, -58, 114, -22, -7, 110, 107, 88, 15, -94, -97, 31, -38, 55, -45, -35, -72, -111, 77, -79, -58, 86, 5, 51, -20, 123, -19, -77, 87, 109, 3, -82, -47, 43, 5, -77, -27, 118, -107, 54, -68, 73, 44, -19, 101, -127, 68, -77, -63, -19, 92, 48, -46, 17, 10, 60, 59, 120, -70, 13, -111, -24, -71, -24, 103, 103, 20, 19, -3, -14, 12, 33, 53, -10, -28, -53, -51, 79, 74, 87, -96, -123, 77, 28, 36, 38, -74, 122, -98, -27, -96, 87, -34, -125, 120, -123, 68, 61, -40, -79, -100, -118, 68, -31, 99, -95, -16, 9, 119, -96, 22, -28, 89, -6, -59, -7, -46, -10, 123, 46, -118, -28, 49, 117, -81, -70, -26, -58, -126, -92, -89, 103, 105, 53, 53, -125, -70, 50, 33, -44, -102, -121, -127, 17, -88, 25, 26, -10, -115, -21, 115, -35, 39, -18, -33, -27, -42, 77, -5, -76, -50, 7, 125, -126, -113, -11, -86, -15, 9, 12, 125, 61, -75, 114, -79, -11, 16, 55, -110, -92, 122, -123, 2, -3, 6, -118, 101, -119, -78, 46, -3, 90, 35, -93, 31, -34, -42, -55, -10, 63, -91, -39, -20, -6, -74, -19, -125, -97, -35, -124, 65, 82, 11, -12, -43, 17, -25, 63, -44, 97, 64, 122, -28, -8, 76, 94, -98, -22, 110, 97, -88, -1, -97, -127, 115, 87, 43, -126, 107, 113, 111, -40, -24, -76, 53, 8, -11, -100, 25, -15, 86, -74, 102, 54, 67, -36, -18, -95, 34, -14, 25, 119, 52, 22, 42, -119, 125, -63, 49, 112, -72, -30, 66, -22, 14, -118, -90, -108, 69, -72, 4, 71, 109, -49, 110, 118, 65, -115, 58, 31, 15, -27, -25, -77, -28, 70, 23, -61, 126, -51, -19, -88, 34, 123, 3, -57, -65, 86, -103, 70, 58, 29, -58, -48, -33, -67, 23, 35, -101, -39, 52, -53, 92, 75, -21, -42, -22, -118, -125, 16, 123, -79, 113, -47, 25, -119, -70, -127, 86, -7, 119, 74, -46, -3, 97, 63, -102, 116, -99, -73, 16, 114, -84, 124, 31, -37, 100, 79, -66, 43, -119, 28, -127, 1, 51, -59, 80, -1, 57, 118, 21, -3, 6, 4, -53, -121, 38, -125, -112, 71, 57, -68, -85, -81, 79, 30, 35, -11, 95, -88, 119, 118, -26, -65, -104, 97, 6, 102, 120, -46, 77, -16, 123, -76, 74, -88, -112, 106, 67, 98, -65, 31, 6, 102, -42, 55, -126, -37, 7, -93, -30, 108, 99, -80, 122, -32, 109, 53, 64, 79, -21, -71, 124, -45, 64, -31, 87, -41, -6, -88, 73, 84, -92, -2, -6, 6, -19, 58, 115, -33, 114, 91, -68, -109, -107, 9, 100, 103, -34, 55, 41, -80, 105, -36, 28, 103, -13, 22, 73, -44, 85, -80, -7, 124, -108, 57, -58, 40, -26, -60, -40, -107, -106, -64, -76, 34, 72, 81, -14, 17, -47, 60, -61, 116, -33, 78, -95, 85, 21, 64, 118, 49, -7, 49, 97, -41, 110, -59, -104, -122, -74, -116, -38, 68, 84, -6, -120, 82, -44, -101, -2, 105, -30, -14, -38, 17, -46, -122, 18, 38, -10, -122, 54, 103, 84, -3, 87, -116, -25, 26, -82, 45, 106, -48, -59, -57, 15, 108, -87, -58, 103, -117, -88, -50, 80, 54, -107, 53, -3, -3, -43, 2, -90, 110, -64, -56, 67, 107, -76, 88, -87, 82, 79, -116, -69, -40, 61, -84, 125, 86, 102, -15, 6, 24, 126, 52, -69, -63, 12, 68, 118, 97, 126, -102, 99, 52, -90, -65, 0, 110, 21, -66, -60, 38, 32, -58, 51, -7, 53, -35, 76, -23, -50, -80, -125, -103, -46, -4, -17, -1, -83, -126, -24, 2, 95, 66, -13, 98, -93, 124, 18, 106, 26, 87, 107, 63, -40, -73, 28, -104, -98, -82, 14, 70, 77, 81, -103, 57, 36, -50, 37, 9, -70, 81, -103, 27, -121, 80, 63, 120, -21, 81, 23, -82, -109, -67, 35, -75, -48, 8, -96, 85, 106, -49, 54, 51, 92, -109, -59, -36, 91, -119, 26, -39, 108, -59, 2, 48, 104, -40, 26, -53, -76, -21, -31, 16, -73, 106, -64, -5, -1, -70, 21, 108, -28, 53, 96, -80, -9, 106, -82, 13, 88, -51, 7, 119, 36, 111, 102, 106, -125, 122, 107, 106, 11, 127, 41, 27, -128, -85, 85, 97, -30, 29, 70, -116, 43, -3, 32, 72, 9, 125, 119, -56, -39, -6, -86, -85, -6, -118, 120, -114, -102, -10, 26, -81, 117, -83, 23, 93, -86, -57, -16, 81, 24, 31, 8, -34, 41, 22, -67, -100, 127, 87, 123, -23, -76, 54, 70, 114, -109, 48, 3, 11, 74, 15, 20, -47, 43, 123, 30, 47, -117, 18, 90, 32, -45, 49, 64, -108, -90, -1, 34, 103, 3, 118, -80, -4, 116, 97, 88, -67, -43, -115, 30, 7, -76, -80, 29, -70, 12, 88, 66, 74, -62, -86, -114, 34, -108, -70, -75, 106, 4, -17, 99, 6, -43, 13, -83, -8, -28, -22, -22, 31, 34, -26, 116, 56, 31, -90, 96, -43, -35, 7, 118, -56, 34, -115, 40, -29, -111, -124, -11, 41, 120, 116, -44, 84, -97, 54, -61, 91, 118, 21, -9, 8, 51, -1, 15, 40, -119, -32, 2, 114, -74, -82, -38, 109, -123, 15, -35, -108, -21, -88, -108, -108, 99, 64, -115, -97, 122, -43, -6, -82, -42, 111, 12, -64, -25, -49, 31, -16, 91, 109, -88, -24, 20, 29, 42, -45, -124, -98, -124, 36, 105, 92, -109, -79, 46, -9, -93, 89, 72, -102, -24, -89, 111, 68, -77, 120, 126, -105, 13, -123, 88, 51, 119, 125, -57, 86, -96, -106, 47, 87, -47, 6, 63, 98, -85, 14, -14, -116, 97, 120, 20, 4, -28, 40, 31, -91, -128, -98, 60, -119, -96, 74, 36, 31, -122, 60, 94, 66, 84, -123, 33, -112, -105, 97, 126, -1, 16, 23, -47, 116, 105, 36, -12, -109, 99, 80, -122, -120, 86, -82, -53, -51, -38, -16, 69, -87, 54, -71, -41, -68, -79, -17, -14, -114, -85, -111, -54, -127, -68, -39, -69, -37, -82, -6, -111, -13, 88, 96, -89, 125, 87, -52, 107, -48, 15, 83, 105, 23, 15, 11, 9, -103, -35, -73, 24, 58, 58, 83, -67, 94, 12, 117, 88, 42, -40, -35, 84, 100, 73, 73, -41, -72, -31, -127, -117, 124, 72, 5, 112, 82, 1, -59, 40, 0, 47, 120, 101, -19, -61, 122, -97, -114, 112, -81, 61, 18, -92, 26, -80, -104, 21, -28, -63, -122, -28, -28, -67, 78, 2, -96, 72, -99, -88, 34, 105, 85, -57, 11, -22, -24, -68, -128, -120, 28, -99, -88, -4, -73, 26, -22, 1, -18, -78, -75, -52, -103, 32, -105, 76, -128, -17, 96, -112, -84, -18, 78, -81, 45, 16, 108, -7, -106, -100, -37, 34, -119, -39, 70, -75, 89, -69, 36, 71, 127, -1, -85, 125, 17, -99, 58, 22, -66, -10, 81, -5, 51, 83, 117, -80, 57, 2, -68, 65, -86, -50, -102, 18, -114, 52, 90, 18, 62, -69, 125, 24, -37, 88, -97, -117, 44, 25, -81, 64, -60, -78, -33, -51, 89, 127, 15, 25, 57, -42, 77, -115, -123, 125, -39, 90, 24, 18, 92, 106, 46, -118, 55, -48, -56, -63, -75, -53, 75, -128, 102, -90, -3, 33, -114, -111, -110, -91, -16, -110, -31, 100, 86, 20, 62, -79, 61, 77, -103, -86, -30, 73, -40, 50, -24, -68, -17, -34, -4, -119, -102, -5, -17, 19, 110, -103, -43, 27, 15, 32, -104, -63, -117, -8, -82, -82, -5, 70, 6, 27, 30, 33, 36, 15, -59, 88, 21, -113, -66, -98, -82, -124, 126, 48, -106, 24, -47, 92, -117, -74, -101, 65, -43, -51, 49, -102, -110, 115, 50, -13, 92, 75, 14, -95, 66, -5, -106, -103, -37, 41, -104, 61, 71, -70, 111, -115, 94, -116, -120, -37, 97, -48, 92, -71, -39, -63, -11, 84, 77, -119, -14, -123, 89, 68, -62, -122, -109, 119, 96, -114, 18, 63, 101, 54, 40, 103, 59, 27, -83, 29, 96, -18, -57, -34, -68, -60, 85, -112, 74, 42, -99, 122, 127, -7, -57, -40, -95, -70, 97, -35, -123, -63, -10, 50, -58, 122, 32, 73, -38, 78, 111, -95, 98, 14, 92, -73, 120, -72, -36, 83, -85, 86, -18, -64, 23, -80, -1, 60, -127, 2, -24, 91, -8, -31, 40, -124, -85, 80, 84, -100, -93, -42, 39, -38, 94, 71, -12, -49, -60, -63, -28, 90, 59, 112, -16, -103, -57, 5, -118, -45, -3, 45, -44, -101, 69, -28, -121, 49, 37, -80, -38, -83, -1, -115, 21, -41, -49, 124, -48, -3, 121, -68, 29, -125, 5, 49, -4, -103, 74, 104, 55, 4, 105, 2, -19, 108, 106, 85, 39, 21, -57, 112, -66, 22, 126, -116, 98, -99, 0, 42, 74, 74, 121, -97, -12, 39, -108, -59, 76, -18, 1, 92, -117, -101, 60, 20, 30, -100, 71, -83, -20, 123, 103, -13, -123, -127, -128, -117, 50, -115, 72, -99, 107, -60, -91, 39, -127, 73, 66, 127, -37, 112, -45, 67, 91, 83, 26, -61, -69, -89, -84, -92, -65, -55, 97, 117, 108, 88, -88, 31, -72, 109, -82, -14, -39, 27, -110, -72, 27, 66, 61, 24, 45, -50, 35, -10, 78, -94, 97, 58, -100, 4, -38, -62, -107, -56, 89, 110, -70, 100, -110, 73, 28, 57, -21, 93, 81, 125, 15, 88, 22, 40, 88, -41, -100, -120, -124, 54, -84, 18, -16, 3, 12, -93, -37, 73, -112, -59, -23, -126, 119, 41, -26, -105, -21, 118, -62, 50, -107, -126, 78, 103, -114, -69, -90, -74, 51, -44, 49, 82, 58, -105, 53, -67, -126, -96, -121, -19, -106, 47, 126, 118, -45, -15, 54, -13, -14, 24, 1, -94, -93, 78, -19, 25, 71, -32, -62, 1, 12, 44, -115, -100, 37, 0, -101, 38, -51, 71, 29, 29, -74, 37, 65, 109, 1, 57, -19, -23, 123, 83, 63, -121, 30, 32, 76, 92, -58, -11, -70, 121, 29, 123, -51, 51, 80, -91, -86, 118, -94, -63, -125, -5, -49, 73, -58, 48, 81, -81, 53, -96, -102, 35, -77, -108, -19, 79, 103, -92, 57, -28, -91, 14, 111, -88, -123, -46, 92, -112, 22, -75, -30, -15, 102, 78, -35, 0, -12, 25, 41, 58, 43, -124, 53, 81, -54, -65, 124, -22, 116, 13, -12, -118, -73, -25, 66, -7, -72, 54, -81, -87, 21, 95, -62, -113, -87, 14, -115, 100, -85, 37, 87, 104, 66, 100, -126, 80, 27, -73, 121, 0, 94, 124, 31, -63, 97, 55, 26, 101, -93, 103, 101, 71, -20, -99, -122, 121, 44, -69, 6, 72, 81, -19, -85, 103, 98, 127, 62, 99, 65, 25, -125, 115, 30, 97, 101, -98, -20, -29, -6, -50, 85, 35, -42, -49, -46, -3, 47, -56, -126, -16, 11, 70, 115, -46, 111, 112, -24, -11, -92, 42, -68, -9, -127, 4, -127, 122, -116, 55, 113, -85, -124, -43, 35, -119, 114, -42, 58, 54, -8, 96, -90, 49, 29, 82, -72, 47, 63, -26, 66, -98, -39, -61, -72, -38, 25, 87, 20, -57, 60, -127, -51, -47, 58, -114, 19, 55, -110, -97, 62, 34, -85, 22, -49, -19, 23, -40, -23, -32, -1, -88, -26, 54, 109, -113, -43, 44, -85, -98, -71, -86, -60, -43, -69, -108, 55, 119, -119, -104, -101, -41, 109, 20, 27, -25, 22, 49, 19, 111, 121, -58, -18, 11, -127, 83, -68, 30, 100, -125, -101, 102, -92, 1, -86, 93, 75, 51, -58, 116, 127, 42, -90, -37, 64, -124, -1, 28, 127, 74, -111, 18, 77, 103, -106, 71, -6, -93, -14, 96, -40, 43, -113, -66, 85, -24, -97, -96, -127, 45, 53, 125, 109, 74, 65, -72, 36, 99, -58, 117, 50, -86, 54, 29, -81, -82, -71, 121, 39, 81, 111, -27, 42, -82, 6, 125, 109, -56, 40, -107, 96, -90, -55, -53, 94, 64, -51, 84, 91, -26, -124, 22, -10, 72, -63, 2, 114, 101, -72, 18, 42, 19, 106, 103, 120, 81, 66, -2, -18, 36, -56, 8, -123, 33, -90, -26, 117, 27, 111, 16, 107, 55, 112, -34, 9, -49, -54, -4, -100, 18, 44, -57, -49, 84, -126, -25, -19, -32, -7, 26, 67, 121, 71, -78, -56, -36, -6, -67, -76, -16, -54, -93, 34, -57, -38, 22, 93, -101, -51, -85, 8, 113, 4, 13, 102, -119, -123, 40, 69, -16, 77, 82, -48, 66, 1, -48, 60, -76, 115, -78, 109, 109, 60, -18, -104, -33, 59, 86, 118, 10, -109, -19, -32, -111, -47, -3, -11, -32, -5, -121, -39, -125, 106, 82, 31, 65, -18, 18, 117, -23, -99, 123, -28, 82, -16, -74, -71, 45, 4, -72, -34, 69, -28, -53, 105, -87, 67, -77, -35, -60, 51, 111, 114, -102, 0, 111, 55, -127, -127, 72, 104, -110, -14, 61, 47, 102, 99, 12, 82, 32, -99, -69, -8, -96, -112, 0, 6, 85, 25, -77, 30, -78, 9, -72, -83, -74, -50, 102, 12, 114, -23, 16, 24, 108, -2, 0, -118, -98, 61, 8, -78, -11, 100, -73, -118, -83, -127, 16, 2, 49, -102, -25, 108, 43, -123, 106, -84, 36, -81, -64, 99, 98, 92, 116, -6, 26, -47, -40, -120, -121, -70, -115, -43, 65, 21, -72, -48, 66, 68, -56, -22, 8, 49, 108, 72, 84, 49, 56, 21, -17, 103, -94, 9, 117, 116, -3, -15, 17, 76, 68, 89, -82, -61, 87, 5, -90, -102, 113, -21, 34, -33, -15, -57, -17, -91, 53, 24, 3, 29, 76, 13, 20, 80, 71, -114, 95, 23, 82, 48, -42, -7, 29, -91, 86, 54, -62, -111, -71, -110, -106, -76, -115, -80, -31, 57, -46, -99, -91, 10, 60, 14, -47, 20, 102, -1, -105, 11, 25, -75, -92, -28, 86, -100, -31, 58, 93, -75, -50, 97, 58, -18, 40, -109, -20, 60, -31, 49, -75, -61, -34, -42, -107, -3, -23, 88, 12, 67, -105, -101, 9, 110, 99, -51, 43, 82, 103, 35, -73, -107, -22, -37, -81, -35, -31, -34, 19, 35, -33, -127, 49, 109, 117, 107, 109, 58, 9, -5, 75, -127, 13, 54, -19, 123, -104, 63, -107, -48, 108, 48, -47, -64, 106, 104, 65, 114, -122, -1, 45, 15, 13, 21, -102, 95, 77, -120, -76, 121, 2, 121, 47, -31, -40, 68, 33, 108, 53, -56, -79, -23, 79, 124, -23, 91, -112, -4, -128, 96, -105, -60, 122, 125, 14, -112, 124, 35, -109, -114, 82, -49, 96, -73, -99, -50, 98, -105, 78, -125, -29, -50, 97, -42, 47, 8, 28, 63, 47, 112, -69, -125, -76, 95, 85, 7, -21, -84, -11, -12, 21, -88, -110, -51, 100, 79, -27, 115, 110, 54, 90, -110, 27, 122, -35, 31, 106, 30, -109, -4, -111, 106, -65, 18, -35, -61, 104, 121, -33, 82, 6, -125, -10, -75, 120, -43, 7, -23, -46, -105, -35, 101, -77, -1, 67, -26, -25, -115, 70, -65, -45, 10, -118, -112, -90, 46, 118, 94, -104, -60, 122, 36, 82, -67, 3, -66, -72, 19, 96, 21, 87, -51, 11, 3, -34, 113, -64, -95, -113, 45, -73, 42, -40, 68, 10, 57, 29, 78, 40, 8, 32, -92, -107, 88, -65, 29, -63, 44, -78, 17, 86, 50, -53, 99, -122, -94, -118, 17, -31, 117, -11, 39, -118, 102, -69, 43, 10, -116, -38, 39, -53, -2, 100, 31, -94, 71, 38, 1, -81, 1, 116, -14, -11, 46, -98, -87, 21, 30, 22, -93, -111, -91, 87, 36, -66, -118, 2, -117, -19, -71, -62, -107, 98, -96, 48, -62, -29, 63, -71, 16, 14, -2, -52, -19, -108, -69, -24, -39, -39, -103, 34, -80, -65, -125, -20, -96, -6, -115, -92, -30, -127, 93, -50, 42, 78, 58, -7, -98, 12, -43, -45, -23, 65, 42, 22, 98, 86, -60, -30, -115, 3, 33, 41, 81, -99, -70, 111, -95, 69, -95, -36, -17, -34, -53, 84, -114, -76, 38, 60, 3, -60, -105, 100, -49, -14, -95, 74, 25, -81, -99, 98, 93, -4, 88, 58, -8, 92, -99, -89, -86, 98, -99, -76, -42, 32, -76, 91, 127, -63, -47, 17, -102, 61, 90, 74, -108, -89, -92, -65, 30, 87, -101, 95, -92, -43, -17, -107, -22, -58, 39, -35, 73, 81, -47, 56, 4, 65, 15, 106, -64, -110, -18, 91, -57, -94, 102, -28, -7, -96, 54, 9, 26, 59, 79, 113, -16, 23, 14, 81, -42, 15, 48, -52, 92, -103, 68, 6, 13, -128, -76, 52, 63, -88, -70, 33, -118, 61, 14, -36, 111, 75, -58, -111, -71, 3, 28, -81, -114, 90, 46, -88, 58, -34, 104, 66, 88, -89, -60, 85, -36, 97, 59, -90, -106, 103, 107, -60, -65, 90, 42, 32, -111, -88, -103, 85, 119, 83, -84, 45, 0, 46, -55, 82, -82, -50, -87, 4, -121, -92, 33, -88, 63, 117, 51, -32, 49, 18, -55, 99, 107, 10, 22, -122, -74, 37, -53, -20, 97, 19, 15, -83, 31, -108, -74, -22, -28, -13, 103, -7, 44, -79, 42, 70, -20, -53, 25, 1, -3, -91, -105, 25, 47, -123, 3, 55, -18, 24, -32, -58, 71, 75, 90, 79, 40, 117, 125, -53, -56, -99, 105, 44, -15, -73, 67, -60, 57, 77, 34, -100, -113, -45, 37, -62, 33, 28, -9, 86, 76, 46, -94, -69, 124, 55, 66, 51, -20, 111, -80, 117, -94, 67, 8, -21, 54, 81, -30, -89, 91, -123, 22, 15, 102, 91, -60, 47, 3, -7, 76, -112, -101, 52, -83, 71, -19, -21, -67, 71, 53, -120, 98, -20, 49, -36, -106, -44, 66, -82, -35, -83, -17, 24, 45, 80, 29, 75, 43, 36, -79, -60, 123, 16, 77, 75, 41, 68, 43, 85, -10, 27, -3, -36, -76, -124, 29, 27, -63, 80, -114, 38, 103, -75, 9, -72, -12, -86, 11, 52, -66, 28, 111, -24, -75, -28, -83, 7, -115, 6, -47, 109, -17, -104, -69, -36, -35, -115, 11, 112, -88, -38, -100, 36, -69, -57, 25, -55, 24, -32, 117, 1, 111, -50, -89, 108, -10, 47, 65, -23, -117, -8, 87, -79, 104, -58, -51, 38, -124, 72, 2, -85, 75, -78, 121, -57, -45, 67, 89, -107, 61, 94, 93, 52, 22, 39, 13, 21, -109, -40, 80, 76, -36, -70, 23, -126, 108, 121, 40, -123, 51, 18, 57, 76, 31, 44, 68, 29, -38, -100, -67, -90, -9, -104, 41, -38, 79, -4, -19, 6, 118, 96, -26, 98, -91, 8, -2, 7, 114, -14, -124, 95, 42, 77, 80, 38, -84, 24, -100, -63, 106, 42, 67, -72, -97, 110, -66, -11, 69, 71, 0, -48, 98, -128, 21, -45, -7, -75, -126, -120, 55, 96, 52, 77, -78, -122, -51, 69, 64, -98, 87, 92, -11, 11, -113, -20, 29, -108, -56, -18, -5, -2, 123, -54, 71, 44, 36, -3, 76, 116, -51, 77, -24, -107, -126, 18, 10, -95, -5, 112, 115, 28, -102, -54, 66, -114, 107, -62, 116, -3, 48, 110, -25, -40, -33, 125, -117, -20, 5, -57, -10, 114, -64, 14, 7, -65, -87, -55, -110, -12, 95, 11, -17, -123, 111, -21, -110, -19, -52, 0, 106, -11, -109, 28, -16, 75, 37, -39, -34, 88, -20, 11, 113, 70, 26, -93, -59, -7, -44, 38, -126, -70, -98, -38, 91, 35, 70, -5, 121, 99, -103, 56, -12, 77, -59, -14, -67, 100, 2, -108, 21, 108, -77, 68, 9, 125, -57, 64, -106, 83, -71, -10, -18, -108, -72, -86, 63, -27, -93, -39, -3, -36, -3, -62, 38, 22, 84, 29, 81, -38, -60, -48, -115, -124, 30, -60, 13, 114, -97, 95, 108, -90, -76, 8, -75, -39, 7, -113, -73, 6, -77, -55, 99, 91, 7, -12, 8, -65, 23, -26, -76, -121, 91, -94, 16, 17, 4, 96, 42, -80, 58, -39, 111, 54, -64, -66, -13, 89, -81, 61, -108, 104, -110, -53, -50, -5, 16, -118, 32, 107, -41, -63, -104, 72, 69, -42, -26, -64, 30, 54, -26, 61, 61, 113, -62, 98, 79, -11, 60, 89, 60, -126, -67, 103, -74, -111, 36, -13, 1, -40, -11, 47, -16, -25, 35, 69, 27, 11, 21, 86, -22, -12, 93, 120, -95, 64, -100, -46, -36, -67, -29, 54, 35, 124, 105, -2, -11, 25, -68, -18, 84, 106, 83, 4, -62, 126, 38, 22, -79, -113, 79, 83, -15, -64, 106, -107, -74, -118, -53, 120, 17, -79, -64, -45, -33, -56, 7, 2, 2, 22, -38, 69, -34, -92, -73, 7, -82, 73, -19, 106, 86, -70, -66, -117, 115, -12, -83, 80, -86, 28, 52, -9, 119, -59, 52, -117, 13, 94, -19, 0, -81, -102, -2, 48, 47, 36, -125, 50, 35, -57, -122, 102, -21, -36, 120, 11, -86, -123, -38, 83, -2, 82, -121, 60, -8, 27, 67, 68, 41, 41, -72, 68, 38, -122, 83, 7, -69, -61, -9, -45, -52, 50, 97, 45, -2, 48, -43, -17, -40, -7, -68, 32, -53, 46, -41, 112, 24, 13, 36, -53, 81, 104, -58, 96, 3, 94, 5, -126, -114, -7, -43, 86, -82, -29, -102, 113, 102, -53, -15, 57, 46, -17, 6, -29, -41, 112, 99, 54, -92, 28, -66, 44, -128, -108, 99, -56, -121, -116, 53, 27, -75, 57, -15, 17, 20, 36, -17, 43, 79, 38, 75, -34, -90, 45, -119, 120, -16, -70, 36, -103, -5 );
    signal scenario_output : scenario_type :=( -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 74, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -108, 127, -128, 127, 127, 127, -10, -128, -22, 127, -128, 127, -128, 102, -128, -128, 118, 127, 127, -128, 127, -128, -128, -128, 127, 127, -88, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 6, -95, -128, -128, 127, 127, -101, -128, -128, 127, -128, -128, 127, -109, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -114, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -87, 127, -128, 60, 127, 127, -128, 127, -128, -128, -128, -128, 11, 65, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 79, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -49, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 33, 127, -97, -128, -128, 127, -128, 127, -128, -128, 127, -26, -128, -128, 127, -128, -128, 127, -128, 0, 127, -128, 127, -128, -70, -128, 127, -90, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -52, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, -128, 79, 127, 127, -128, 78, 127, -65, -128, 127, 113, -128, 127, -53, -128, 127, -68, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -100, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 37, -128, 127, -111, -128, -128, 127, -128, 127, -97, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 47, -128, -7, 127, -128, 27, 127, -128, 127, -128, 49, 127, -128, -128, -128, 127, 127, -128, -42, 127, -128, 39, -128, 127, 17, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -22, 127, -128, -128, 127, 90, -128, 127, 127, 127, -60, -128, 42, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -109, 127, -128, -128, -58, -39, 127, -128, 127, -128, 127, -128, 12, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -43, 8, 127, 127, -128, 127, -128, -108, -128, -128, 127, 127, 127, 127, 127, -44, -11, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -50, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -88, -128, 127, 127, 11, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -107, -128, 127, 127, -128, -128, 127, 96, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 74, 127, -128, 108, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -119, 27, -128, 127, -128, 127, -128, -128, 54, -128, -128, 127, 127, -128, -128, -128, 127, -128, -80, 127, -128, 127, -128, 127, 127, 86, 127, -128, 127, 127, -128, 127, 127, -128, 127, 109, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -95, 127, 103, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -98, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -6, -128, -128, -123, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -6, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -109, 127, 127, -128, 127, 127, -69, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -118, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -68, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 37, 127, -128, 127, 127, 127, 127, -128, 127, -128, 87, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -76, -58, -103, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 57, -128, 127, -128, -128, 127, -128, 127, -11, -128, 127, -36, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -8, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 100, 127, -128, 127, -128, -128, 127, -128, -66, 127, 127, -128, -112, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 2, -128, 127, -100, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -60, 127, -128, -128, -128, 127, 127, -6, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 85, 127, -85, -128, 127, 127, -128, -128, -128, 127, -128, 127, 42, -128, 127, 127, -128, 127, 127, 127, -128, -128, -54, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 97, 127, -128, 127, 31, 11, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -33, 127, 48, -2, 127, -122, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, 55, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -23, 127, 127, 127, 64, -128, 127, -128, -128, -13, -128, 127, 127, -128, 7, 127, -128, 127, -128, 127, 127, -93, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -53, 127, -128, 127, 59, -128, -128, 78, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 79, 127, 64, 127, 127, 127, 127, -128, -26, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -106, 15, 127, 64, -16, -128, 127, 127, -128, 127, -16, -128, -128, -128, 127, 127, -128, 127, -128, -128, -117, -128, 127, -128, -28, 127, -128, 127, 127, -128, 127, 127, 127, 29, 127, 127, -128, 127, -128, -128, -128, 15, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 1, -17, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 78, 127, -117, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 63, -128, -102, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 66, 127, 127, -128, 127, 127, -128, 127, -128, 88, -128, 127, -128, 127, -128, 68, 127, -128, -122, -128, -128, -128, -128, -128, -121, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -118, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 11, 127, 127, -128, -128, 127, 127, 127, -128, -128, 17, -128, 127, -128, -42, -128, 58, 127, -128, -128, 75, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 60, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 54, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 76, -128, -128, -128, 127, -128, -12, 127, -128, -85, 127, -128, -128, 127, -8, -128, 127, -128, 127, -128, 127, 43, -128, -21, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -100, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -8, 127, 127, 127, 6, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 34, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 100, 127, -128, -128, 59, -128, 127, -128, 127, -128, -68, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -55, -128, 127, -128, -128, -128, 119, 93, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -2, -128, -128, 127, 127, -128, -128, 127, -36, -21, 127, -24, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -117, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, 88, -71, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 26, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -76, -128, 127, 127, 127, -88, 127, -128, -128, -112, -128, 127, -128, 127, -128, -128, -128, -128, 112, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 119, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -95, -128, -128, -128, -75, 127, -128, -128, 127, 70, -128, 127, 127, -128, 127, 127, -55, -128, 127, 127, -128, -21, 127, -128, 127, 127, -128, -128, -128, -128, 13, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -68, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 28, -128, -128, -128, 127, 127, -128, 76, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -43, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 22, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -95, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -45, 127, -128, -128, -128, 127, 127, 92, 127, 127, -128, -128, 127, 127, -127, 127, -128, -6, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -49, -128, 88, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -11, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -88, 127, -128, -8, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -118, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 95, -128, 127, -128, 127, -128, -128, -128, 127, -128, 49, 127, -128, -128, 127, 127, 127, 127, -128, 27, 127, -128, -128, 127, 114, 127, -128, -128, -111, -128, 127, -128, 118, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -29, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -86, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 81, 127, -128, -128, 127, -128, -128, -128, 127, -73, 0, 127, -128, 127, -128, 127, -128, -128, 54, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -27, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 21, 127, -128, 127, 127, -128, 127, -128, 37, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -44, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 10, -128, -128, 127, 127, -12, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 73, 112, 127, -128, -128, -128, 127, 59, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 121, 13, -128, 127, 127, -128, 127, 127, -128, -128, 127, 103, -128, 127, 127, -128, 127, -128, -128, 127, -128, 68, -128, -128, -128, -128, -128, -128, 127, -128, 127, -79, 106, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -79, -128, 127, -54, -128, 127, -128, 127, 127, 127, -114, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 8, 127, -128, -128, 127, -128, -128, -113, -128, 38, 127, 15, -128, -128, 127, -92, -128, -128, 127, -128, -128, 111, -128, 127, -128, -128, 127, -128, -128, -96, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -78, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -21, 127, 21, 127, 127, 127, 127, 127, 127, 127, 127, 15, 127, 127, -66, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -92, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 39, 127, -128, 127, 68, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 26, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -64, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -91, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -108, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 92, -128, 127, 124, 127, -128, 127, -128, -128, 127, 32, -128, 127, 127, -128, -128, 127, -15, 127, 112, -128, -128, -128, -128, 127, 127, -128, 127, -87, -128, -119, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 57, -128, 127, -128, 127, 127, 18, -128, 127, 127, 127, 127, 127, 127, -128, 127, 71, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 100, 127, -128, 95, 127, 127, 92, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -79, -128, 127, -128, 127, 127, -128, 127, 127, 6, -128, -29, 127, -128, -128, 127, -128, -128, 73, 127, -50, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 78, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -31, 127, -128, 127, -128, -117, -128, -128, -128, -128, 127, 127, -128, -128, 127, 91, 79, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 90, -128, 63, -128, 127, -128, -128, 127, 78, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 108, 127, -128, 127, 85, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 33, -128, -128, 127, 127, -128, -128, -53, 127, -128, 127, -128, 127, -128, -128, 127, -128, 108, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 101, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 42, 127, 127, -128, 127, -128, -128, 71, -128, 43, 117, 28, -128, 127, -128, -128, 127, -24, -128, 127, -128, 127, -128, -128, 127, -128, -128, 111, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 26, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -13, 127, -128, -128, -113, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 80, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -90, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 116, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -92, -128, 15, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 98, 127, 127, -128, -128, 127, -128, -128, -128, 114, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 93, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -8, 36, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -66, 127, 127, 127, -128, 118, 127, 33, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 93, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -22, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -10, 127, 127, -70, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 26, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -34, 127, 3, -128, -128, 127, -128, 127, 127, -128, 107, 81, -123, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -18, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -85, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 114, 127, -128, 127, -5, -128, 127, -128, -128, 127, 127, -29, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 23, 127, -79, 127, 127, -52, 90, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -76, -128, 127, -128, 127, -128, 127, -128, 127, 127, -16, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 79, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 80, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 76, -128, 87, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 100, 29, -128, 127, -86, -128, -128, -128, -128, 127, 127, -128, -93, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 76, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -49, -128, -128, -44, -50, -123, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 71, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 79, 127, -128, 3, 127, -128, 127, 127, -128, -3, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -111, -128, 127, -128, -128, 37, -128, -17, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 10, 127, -128, -128, 68, 8, 127, -128, 127, -128, 127, 127, -87, 127, -128, 86, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -121, 127, 34, -128, 127, -128, 127, -128, 127, -128, -128, -107, -128, -128, 127, -128, 127, -128, 127, 127, -12, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 15, 127, -128, -73, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -70, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, 16, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -60, 127, -37, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 59, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -42, -128, -128, -128, -128, -128, -128, 127, 127, 59, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -24, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -86, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 102, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 73, -128, -128, 127, -16, -128, -128, 127, -128, 127, 106, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 60, 127, -100, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 73, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -39, 127, -128, 127, -128, 127, 127, -128, 127, 76, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -122, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -15, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 63, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -18, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -123, 127, 127, 127, -128, -128, -68, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 49, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -11, 109, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -106, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -107, 127, -128, 124, 127, -29, 127, -128, -128, 127, -128, 127, -128, 6, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 111, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -93, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 70, -128, 127, -31, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 118, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 98, -128, -128, -127, 127, 127, -128, -128, -128, -49, -98, 127, -128, 127, 127, -53, 127, 127, -13, 127, -128, 127, -119, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 64, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -16, 127, -59, 127, 127, 127, -128, 127, 127, -128, 74, 127, 45, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 36, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -59, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -13, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -48, 127, -128, 127, -106, 127, 127, 127, 127, -128, 127, -128, 13, 127, -128, -128, -128, -122, -128, -128, 127, 127, -69, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -23, 127, -128, 127, -128, -128, 127, -128, -2, 127, 127, -128, 86, 127, -128, 127, -128, 127, -128, -128, 127, 98, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -17, -128, 63, -128, 127, -128, -128, -128, -128, 127, 117, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 23, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -45, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 102, -128, -128, 127, 69, -128, 127, 127, -128, -16, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -60, -128, 52, 127, 127, -128, -128, 127, -128, 127, 127, 5, 127, 127, -128, -128, 127, 127, -128, -128, 127, -66, 127, -128, 127, -128, -128, 127, 32, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 0, 127, -128, 127, 10, -128, 127, -128, -128, -78, -124, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -96, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -68, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, 86, -128, 127, 127, 17, -128, 127, -128, 127, 127, 96, -88, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -113, -128, 127, 127, -128, 127, -128, 127, -64, 127, 127, -128, -128, -128, -122, -49, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 64, -128, 127, 127, 7, -24, -128, 127, 127, -128, -128, 127, -8, -128, -128, 90, -128, -128, -128, -128, -128, -128, -128, 127, -97, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 39, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -2, 8, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 76, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -100, 127, 127, -128, 127, -128, 127, -128, 127, -64, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -54, 127, -128, -128, 127, 127, -128, -128, 127, -109, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 114, 127, -128, 127, -43, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 59, -128, 127, 81, -128, 75, -54, 127, 127, 127, -128, 127, -128, 3, 127, -128, 127, -112, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 50, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -116, 127, -128, 127, -113, -128, 127, 127, -128, 127, -128, 127, 57, -128, 127, 127, 127, -128, -128, 127, -128, 103, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -50, -6, 127, -128, -128, 127, -128, -128, 75, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -81, 127, -34, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -87, 127, -15, -128, 127, -128, 127, -128, 124, -2, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 69, 118, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -59, -128, -128, -128, 127, -128, -45, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 119, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -34, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -3, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 103, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -52, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -17, -128, -128, 127, -128, 127, 127, -128, -128, 127, 32, -128, 127, -128, 127, 127, 12, 127, -128, 127, 127, -48, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -32, 127, 39, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -29, 127, 54, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, 76, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 3, -34, -128, 127, -128, 127, -128, -13, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 22, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -6, -128, -128, 122, -128, 127, -128, -128, -128, -128, -128, 127, -128, -69, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -95, -128, 127, -128, 127, 29, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -122, 127, -128, -128, 86, -128, -128, -128, 127, 75, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 0, 127, -128, -102, 127, -128, 127, -50, 127, 32, 127, -121, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 95, 127, -128, -128, -128, -128, -102, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -34, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 98, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 47, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 101, -128, 127, -128, 127, -50, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 96, 127, -128, 75, 18, -26, -128, -128, 116, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -6, -128, -38, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -117, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -36, 127, 127, -128, 127, 127, -128, 127, 127, 127, 101, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -8, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 13, 127, -65, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 53, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -63, 127, -128, 127, -127, 127, 127, -128, 95, 127, -128, 127, 127, 127, -128, -128, -128, -11, 127, -128, -90, 127, 127, -128, 127, 127, -128, -128, 127, 43, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 38, 127, 127, -128, -49, 127, -128, -128, -128, 127, -128, -128, 127, -31, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -47, -79, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -16, -128, 127, -128, 127, -128, 127, -128, 127, -98, -128, -128, -128, 127, 127, 127, -128, 127, 127, -98, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, -23, -128, 37, -128, 127, -128, -128, 127, -128, 127, -128, -128, -100, 127, -128, -128, -2, 58, 127, -128, 98, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -53, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 63, 127, 48, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 8, 127, 127, -3, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -34, 127, -128, 127, -128, 117, 127, -73, -128, 127, 127, -128, 127, -128, 38, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 107, 127, -128, 127, -128, 127, 127, 127, -119, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 65, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 0, -128, 127, 127, -128, -15, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 114, 127, 127, -128, 85, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -74, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 123, 127, -128, 127, -128, -59, 127, -111, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -109, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 50, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 69, 0, -128, 127, 127, -128, -92, 127, -128, 127, -128, -128, -128, 127, -128, 127, 1, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -64, -108, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -24, -128, -128, 96, 127, -128, -28, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 63, -128, -128, 86, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 95, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -38, 127, -128, -128, -128, -128, -128, 127, 127, 24, 127, -128, 127, 0, -128, -43, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 78, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 27, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 28, 127, -128, 127, -128, 127, -71, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 53, -128, 127, 127, -128, -128, -128, 127, -128, 127, -29, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -75, 123, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -91, 127, 127, -128, 127, -128, 127, 90, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -98, -128, -128, -10, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 54, -93, 127, 127, -128, 127, 127, -128, 127, -128, -29, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 2, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -98, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -88, -128, 5, -128, 127, 127, -128, 127, 127, -128, 127, 28, 127, -50, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, -54, -128, 127, 127, 127, -128, 127, 127, -128, 127, -11, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -109, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 44, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -21, 127, -128, -98, -128, 127, 127, -128, 127, 127, 124, -128, 127, 127, -100, -128, -128, 7, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 112, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -38, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -98, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 16, 127, -128, 127, -128, -128, -128, 127, -128, 44, -128, 127, 127, -128, 127, -128, 80, 127, -50, 127, -128, -7, 127, -128, -128, -15, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -118, -128, 127, -128, 107, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 39, -48, -128, 127, 127, -128, 52, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 90, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -15, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, -71, 58, -128, 87, 127, 127, -128, -128, 127, 127, 127, -128, -75, 127, 127, -128, 127, 127, -48, 127, -128, -128, -128, 127, 127, 127, -128, 127, 54, -128, -128, -128, 93, 127, -128, 127, -128, 127, -58, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 121, 127, -128, -128, 127, -128, 127, -128, -128, 127, -27, -128, -128, 127, 111, -128, 127, -128, 127, -128, 127, -128, -128, 127, 76, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -73, -97, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 31, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -80, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -112, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 97, 127, 112, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 91, 127, -128, -128, 127, 127, 127, -114, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -75, -128, 127, -128, -128, 127, -128, 127, 13, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 52, -128, 101, -68, -128, 127, -128, -128, -128, 114, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -97, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 102, -128, -16, 127, 127, -128, -128, 127, -108, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -65, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 53, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 26, -66, 127, 127, 127, -128, 127, 54, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 60, 127, 127, 121, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 13, -44, 127, -128, -128, 127, -7, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -81, 127, -128, 127, 127, -128, 127, 71, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -101, 127, -128, -128, 127, -128, -6, 127, -128, -128, 113, 127, -128, -128, -128, 127, -128, -91, 127, -128, 127, 127, 127, -128, -128, 127, -103, 127, -128, 127, -128, 127, -128, 127, -128, -111, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -44, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -39, 127, 127, 127, 102, 127, -128, 127, 88, -128, -128, -128, -128, 127, -128, -128, -128, 127, -127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -38, 127, 127, -128, 127, 127, -128, -128, 127, -52, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -57, 43, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -85, 127, -128, -66, 44, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 90, -128, -128, -128, -128, 127, -128, -8, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -3, -128, -128, -128, -128, -85, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 43, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 76, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -6, -128, 127, 43, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -54, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -92, -53, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 34, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 86, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -95, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -11, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 42, -42, 127, -128, 127, -128, 127, -128, 127, -128, 127, -86, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 29, 127, 15, 127, -128, -128, 127, -128, 48, 32, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 111, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 54, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 85, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 96, -128, -123, -128, -128, -128, -128, 127, 91, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 28, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -90, 127, -128, -27, -128, -128, -128, 53, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 109, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 38, 37, -128, 127, 127, -128, 127, 127, -128, -52, 127, -128, -128, -128, 127, -128, -128, -11, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 10, -128, -128, 127, -128, -128, 127, -128, 0, -128, 127, 127, -95, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 68, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -65, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, -118, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 32, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 55, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -112, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -24, 71, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -5, -128, 127, -128, 127, -65, -128, 127, -128, -128, 57, 127, -128, 127, 127, 127, 127, 49, 127, 127, 68, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -1, -128, -128, 127, 127, -21, 127, -128, 70, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -117, -128, 127, -71, -128, 127, -128, -128, -91, -128, 127, -128, 127, 26, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -69, 127, 127, -112, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -43, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -22, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -7, -128, 127, 127, -128, -1, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -90, 127, -81, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -85, -128, 127, 127, -128, 127, -128, 16, 127, 127, -128, -128, 127, -128, -128, -24, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 101, -128, 127, 85, -128, 127, -118, -26, 127, -128, 127, -73, -128, 127, 127, 127, -128, -93, 127, -128, 127, -128, 127, 127, -128, 127, 127, -114, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 18, 107, 127, 6, -128, -128, 127, 127, -128, 98, -128, 27, -128, -29, 127, -128, -128, -128, 127, -128, -42, 127, 127, 127, 127, 127, -108, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, -43, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -55, 127, -128, 127, 127, 127, 127, 127, 127, 127, 7, 127, 53, -128, -24, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 101, 127, -128, 127, -128, -124, -128, 127, -128, -112, 127, 127, -63, 127, -128, 127, 127, -128, -11, 127, 127, 106, 127, 127, -8, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -121, -128, -128, 127, 127, -128, 127, -128, 39, 127, 127, -128, 31, 127, 127, 127, -128, -128, -65, 127, -128, -21, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 85, -128, 127, 127, -127, 127, 87, -128, 69, 108, -128, -128, 127, 127, -128, 127, -128, 78, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 97, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 38, -128, 127, 127, 127, -128, 97, 127, 127, -128, 127, 127, -128, 127, 87, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 75, 127, 127, -128, -49, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 90, 127, -128, 127, -128, -128, 127, -128, -128, -128, -87, 127, -128, -128, -128, 10, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 98, -128, -106, 127, -128, 127, 127, 127, 127, -128, 127, -45, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -32, -128, 127, 127, -128, 57, 127, -128, -128, 48, -128, 127, 127, -128, 107, 107, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 54, -128, 127, 127, -128, 26, 127, 127, -128, 33, -100, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 74, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -76, -50, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -87, -128, 127, 16, -128, 127, -112, -128, 127, 127, -128, -128, -69, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -32, 96, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 106, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 85, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -57, 127, -128, -36, 127, 127, 127, -64, -128, 127, 127, 106, -128, -32, -98, -58, -128, -128, 127, -1, -128, 66, -128, -128, -128, 122, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 112, -128, 127, -128, -128, 127, -128, 127, -128, 32, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 117, 127, 127, 127, 127, -128, 127, -128, 34, 127, 127, 31, 127, -80, 127, 31, 127, -128, 127, -128, 127, 45, 127, -128, -128, 127, -128, 127, -128, -128, 127, 15, 127, -128, 127, -128, -128, -128, -121, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 24, -128, 108, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 109, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -96, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 93, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -93, -128, 127, 127, -128, 69, 127, 127, 127, 127, 127, -128, 31, 127, -128, 127, 127, 127, -128, -26, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 63, 127, -128, -117, 127, 127, 127, -128, 127, -128, 112, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -113, 117, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 15, 127, -128, 127, 127, -128, 127, -128, -128, -128, 28, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -74, 127, -128, 127, 127, -128, 127, 127, -8, -128, 127, 127, -128, -128, -128, 127, -128, 127, 57, -128, 127, 127, -128, -128, -3, -128, -128, 127, -128, 127, 0, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -114, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -76, -128, 127, -128, 127, -128, 127, -128, 6, 127, -128, -128, -128, 127, 127, -128, 127, 97, -128, 127, -128, 98, -106, -128, 127, -128, 127, -128, 86, 127, 127, 26, -128, 127, -128, -68, 127, -128, 127, -128, -78, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -100, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 22, 127, -128, 127, -128, 127, 127, -128, -128, 11, -128, -128, 127, -128, -128, -128, 127, -128, 127, 55, 127, -69, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 53, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 76, 127, -128, -128, 127, 17, 127, 127, 39, -128, -128, 127, -128, -128, 127, 57, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 101, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 86, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 114, 127, -128, 127, -128, 127, -100, -128, 127, 127, 127, -128, 127, 127, -5, -78, 127, -128, 127, 127, 24, -128, 127, 127, 64, 16, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -66, 127, 127, -128, 3, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 113, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 42, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 121, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 88, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -53, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -81, -128, 127, -128, 127, 127, -128, 127, -128, -31, -128, -128, 127, -97, -128, 127, -68, -128, -128, -128, 127, 113, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 45, -128, -128, 127, -128, -128, 127, 108, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -34, -128, -128, 127, 127, -128, -128, -128, 23, 127, -128, 127, -128, 71, 127, -128, -128, -128, 127, 65, -128, 127, -128, 127, 127, -59, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 81, 127, -128, 127, -128, 127, -128, -128, 127, 119, -128, -128, -128, 127, -128, 18, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 57, 127, -128, -24, 127, 127, 127, -128, 127, -128, -128, 123, 127, -128, 127, 127, -128, 127, 127, 127, 127, -91, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 49, 127, -128, -128, 127, -128, 114, -128, -128, 127, -128, 127, -128, -128, 112, 127, 127, -128, -128, -128, 127, 127, -108, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 38, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 17, 127, -128, 127, -128, 114, 127, -128, 127, 127, -128, 127, 127, -128, -128, 96, 127, -128, -128, -128, 127, 124, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 96, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 24, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -90, -50, -128, 127, -128, 127, 127, 127, 127, -54, -128, 127, -128, -128, 127, -128, 127, -113, -128, 113, -128, -128, -128, -55, 127, -128, 127, -33, 127, -128, -128, 127, 127, 127, 127, -112, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -91, 127, 127, -91, -128, -128, -128, -128, -128, -128, 74, -128, 127, -128, 70, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -12, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 17, 127, 127, -128, 127, -128, 127, 127, 127, 44, 127, -128, 127, -128, 127, -128, 127, -80, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 95, 127, 127, -128, 127, 127, -128, -128, -128, -128, -29, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 114, -128, 127, -128, -128, 127, -128, -128, -128, 127, 29, -128, 127, 127, -128, -128, -128, 59, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 21, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 108, 127, -128, 127, 48, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -53, 127, 79, -118, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 73, -128, -128, -128, 127, 127, 117, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -29, 127, -128, -128, 127, 127, -128, -128, 34, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 102, 127, -28, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 97, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, 109, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 21, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -38, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 29, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 0, 127, -128, 127, -98, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 7, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 114, 127, -128, 127, -128, -74, -128, 127, 127, -128, -128, 127, 127, 69, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 124, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 21, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, 75, -128, -128, 127, 28, -128, 127, -128, -128, -128, -128, 17, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 3, -128, -69, -128, 127, 127, 127, 127, -128, 127, -128, 127, 92, 127, -128, 127, 127, -128, 127, 127, 127, 127, -16, 127, -128, 127, -128, 127, 127, -128, 127, 68, -128, 127, -119, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 101, -128, -128, -26, 127, 127, 127, 127, 127, -128, 127, 127, -71, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -78, 127, 127, -128, -128, 127, -128, 127, -101, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 106, -128, 127, 127, 10, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 26, 127, -128, -128, 127, 91, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -71, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 38, 127, -63, 127, -128, -128, 127, 127, 70, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 70, -128, 127, 121, -128, 127, -128, 127, 127, 127, 36, -128, -128, 127, 127, -128, -128, 127, 127, 37, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -78, -98, 127, -128, -128, 127, -128, 127, -128, -128, 38, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -64, 127, -128, -128, 127, 127, 54, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -80, 127, 127, -128, 127, -128, 7, 100, 127, -128, -128, -97, -128, -128, 127, -128, -128, 127, -128, -128, 63, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 70, -128, 127, -128, -128, -100, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -22, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -2, 127, 127, -128, 127, -128, -128, 95, 127, 127, -128, 127, 45, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 90, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -37, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 5, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 92, 127, 127, 127, 127, 127, 127, -128, 96, 127, -128, -128, 127, 127, -128, -128, 127, -117, 127, -128, -128, 127, -128, -128, -128, 127, -128, -79, -128, 95, -128, -70, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -121, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 123, -128, 127, 63, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -91, -128, -66, 127, 127, -128, -128, 127, 127, -128, 60, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -103, -71, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -108, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 79, 64, -95, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -118, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -6, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -108, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -33, -128, -109, 127, -128, 127, 127, -128, 127, 18, -128, 127, -128, 127, 127, 1, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 18, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -113, 127, -106, -128, 57, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -32, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 63, -128, 127, 127, -128, 127, -128, -128, 127, 127, 26, -128, 127, -128, 127, 127, -128, -2, -112, 127, -128, -128, -128, 127, 127, 127, 127, -26, -128, 127, -128, 55, 127, -128, -128, 127, -128, -128, -87, 127, 127, -128, -128, 127, -128, 127, -70, -128, -128, 127, 127, -128, -128, 70, -128, 86, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -102, 127, -128, 127, 127, -128, -73, 127, -128, 127, 127, -128, 127, -23, -128, 127, -128, 127, 127, 127, -128, 127, -78, -128, 127, -128, -128, 127, -128, -16, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -116, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -68, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, -44, 127, 127, -24, -128, -128, 127, 127, -128, 127, 127, 127, -60, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -59, 127, -128, -74, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -116, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -26, -128, 127, -128, 127, -128, -128, -50, 127, -128, -96, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 49, 127, 127, 78, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -13, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 106, 127, 127, -128, 127, -128, -128, 127, 95, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, 119, 127, 127, 127, -128, 127, 127, 127, 127, -10, 127, 22, 127, -128, 127, -128, 127, 64, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 88, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 60, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 5, 127, 127, 127, 127, 127, -128, -128, -128, -128, 111, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 117, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 97, 127, -128, 127, 127, -128, -128, 127, -128, -65, 127, -128, 80, -128, -101, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -42, 127, 127, -58, 127, 127, 127, 127, -128, -117, 76, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -116, -128, 127, -128, 127, -128, -37, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -7, 127, 10, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 2, -128, 127, -128, -128, 127, 127, 127, 36, -128, 127, 127, -128, 127, -73, -128, -128, 127, -128, 127, -128, 127, -128, -71, 127, -128, 127, 127, -128, 127, -128, -111, -128, 22, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 101, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -85, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -98, -128, -7, -128, -128, 127, 127, -128, 127, 127, 127, 127, -17, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -16, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -6, 127, -128, 127, 127, 127, -36, -95, -128, 127, -128, 127, -128, -36, 127, 127, -128, 3, 127, -128, 127, 127, -48, 93, 127, -128, 127, -128, 127, 127, -128, -69, -128, 127, 127, -128, -128, 127, -128, 127, 64, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 96, 127, -121, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 13, -128, 127, -36, -128, 127, 64, -128, -128, 127, 127, -128, -128, 127, -116, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -7, -128, 127, -128, 127, -128, 33, 127, -128, 127, 36, 127, -128, -128, 127, 95, 13, -128, 127, -128, 127, 127, -128, 127, 27, 127, -128, 127, -128, 127, -128, -79, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 121, -128, 127, 111, -128, -128, -128, -128, 127, 127, -128, 127, -50, -128, 127, 127, -128, -128, 127, 127, -128, 127, 93, -128, 127, 127, -128, 44, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 50, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 102, -128, -128, 127, 127, -128, 127, 33, -128, 127, -128, 127, -34, 127, -128, -85, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 90, 127, -128, -128, 127, 127, 127, -128, 65, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -85, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 21, -128, 127, -128, 127, 127, -128, -59, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -63, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 31, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -109, 80, -128, 127, -128, 127, 127, -128, -128, 50, 98, -128, -128, 127, -128, -79, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -81, -128, 127, 127, 127, 127, 127, 127, 27, 127, -127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -103, 127, -128, 127, -53, -128, -128, -128, 60, -128, -128, 127, -128, -128, 127, 100, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -26, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 50, 127, 127, -128, 127, 127, -128, -128, 127, 87, -128, -128, 127, -128, 127, -128, 80, -128, 127, -128, -128, 127, -128, 127, -93, 127, -128, 127, 127, -98, -128, -28, 127, -128, -128, 127, -128, -128, 1, -128, 127, -128, 127, 127, -128, 44, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 98, -128, 127, -128, -128, 127, 127, -49, -128, -21, -128, -128, 127, -128, 127, -57, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 2, -128, -128, 127, -96, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 114, -128, -47, 127, 127, 127, 127, -76, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 93, 127, -128, -128, 127, -128, -128, -128, -128, -128, -98, 127, -128, 127, -128, -128, 127, 0, -58, -128, 127, 127, -128, 127, 127, -128, 127, 127, 85, 127, -128, 78, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -21, 101, 127, 127, 92, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -97, 127, -39, -37, 127, -128, 52, -128, 127, 127, -128, 34, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -49, 127, -17, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 92, -128, -128, 127, 127, -128, -128, 127, 64, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 52, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 2, -128, -128, -128, 127, 127, 127, -128, -128, 109, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 103, 127, -69, -128, -128, 127, 127, -128, 127, 127, -128, 127, -91, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, 31, -128, 127, 127, 127, 13, 127, 127, 127, 127, -128, -128, 17, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 49, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -2, -128, 127, -15, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -69, 127, -128, 127, -128, 127, -39, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -22, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 97, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -101, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -75, -128, -128, 127, -128, -128, -1, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 18, -128, -128, 127, 127, 27, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -43, 55, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -60, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -78, 127, -38, -128, 127, -128, 28, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 71, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 123, -54, 127, -128, -90, -128, 86, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 44, -128, 127, 127, 127, 117, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 32, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -101, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 79, 127, -128, 127, 106, 127, -128, 33, -128, -128, -128, -18, 53, 127, 127, -128, 127, -128, -128, 127, -128, -36, -128, -128, -128, 127, -32, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 93, 127, 127, 127, -128, -128, 127, -36, 31, 127, 127, -128, 127, -128, 127, 127, -128, -128, 6, 127, 53, 127, 127, 127, -45, 127, 127, -128, -52, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -98, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 58, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -2, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 117, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -102, -48, 127, -128, 127, 127, -128, 127, -128, -128, -68, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -97, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 65, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -121, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 39, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -96, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -52, -34, -128, 127, -128, 127, -128, 60, -128, -128, -128, -128, -128, 127, 127, 26, 127, -32, 127, -128, -128, -7, 127, 106, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -91, -128, -128, -128, 127, 127, -128, 57, 127, -128, -128, -128, 119, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -109, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 36, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 22, 127, -128, 127, -128, 127, 127, 127, -63, 127, -128, 127, -128, 127, -128, 100, 127, 127, 127, 81, -128, 127, 127, -128, 127, -128, 127, -128, -29, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -70, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 36, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 45, -128, -128, 127, -128, -128, -128, 127, -45, -128, -128, 127, 127, -128, 127, 127, -128, -111, -101, -128, 127, -128, -128, 10, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 73, 127, -128, -128, -128, -111, 127, 127, 127, -74, -128, 127, 127, -128, 127, -128, 127, -128, -112, 127, -128, -128, -85, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 11, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -50, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -86, -128, 69, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -43, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 1, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -78, -128, -31, -12, -128, 127, 73, 127, -5, -128, 127, 127, -128, -128, -128, -57, -128, 127, 127, 81, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 49, 127, -5, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 33, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -127, 127, 93, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 12, 127, 127, 127, -128, 127, 69, 127, -128, 127, 127, -128, 127, 119, -128, -128, -128, -128, -73, -128, -128, -128, -128, -128, 127, 127, -128, -50, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 60, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 44, -128, -128, 127, -128, 127, 127, -128, 127, -128, 59, -128, -128, 127, 127, -128, -128, 127, -128, 38, -128, -128, 127, -128, -128, 127, -68, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -47, -128, 127, 127, 127, 96, 127, 127, 127, -128, 127, -128, -128, -18, 127, -128, -28, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -11, -91, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 117, -128, 127, 127, -33, 127, -128, 127, -1, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 101, 10, -128, 127, -128, 127, -128, 127, -128, -63, 127, 127, 127, -128, -2, 38, 127, -128, 127, 127, -128, -128, -128, 127, -60, -128, 127, -63, 127, 127, 127, 127, 127, 52, -128, -49, -52, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 81, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 69, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 93, 127, 127, -128, 127, -128, 127, 27, -128, 127, 127, -128, -128, 127, -128, -103, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 45, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -47, 21, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -50, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, -58, -128, 112, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -103, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 50, -128, -128, -128, 127, 127, -128, 127, -128, 11, 127, -128, 127, 127, 127, -128, 127, -74, -128, -27, -128, 127, -128, 37, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -78, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 121, 127, 42, -128, -128, 127, -128, -128, 127, 127, 47, -128, 127, -128, 127, -128, -43, 38, -128, -128, 127, -32, -128, 127, 111, -128, 127, -128, 127, -78, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -108, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 93, 3, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -33, -128, 88, 100, 127, 127, -128, -112, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 0, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -124, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -124, 127, -128, 127, 127, -128, 127, 127, 42, -128, 127, -128, 127, 127, -128, -128, 127, 58, -128, 127, -128, -128, 127, -128, -128, 127, -128, 95, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 69, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -80, -128, 127, -34, 127, 127, 127, -128, 127, -5, -128, 127, 118, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, -11, 127, 127, 127, 127, -128, -36, 127, -128, -69, -128, 127, -128, 127, -128, -32, -128, 127, -128, -128, -11, -79, -128, -128, 127, -128, 123, 127, -128, -128, 127, -128, -128, 87, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 23, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 22, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 102, -128, -128, 127, -128, -128, -128, -128, 64, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 59, -128, 127, 127, -128, -128, 127, -128, -128, 127, 66, -128, 127, -128, 53, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, 33, 127, -27, -128, 127, -128, -7, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 109, -50, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -90, -128, 127, -128, 127, -128, -128, -128, -66, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 101, -128, 127, -128, 127, -128, -128, -8, -128, 127, 127, -128, 127, 127, -128, -128, -54, -128, 127, 31, -128, -49, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -109, -128, 38, 127, -128, 127, 45, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 85, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 116, -128, 127, -128, -128, 127, 127, -128, 127, 16, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -3, 109, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -2, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, 127, -22, -128, 127, -113, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, -128, -48, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -18, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 2, -128, 127, -128, -128, 127, 127, 127, 127, -128, 2, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, -52, -128, -128, 127, -128, 107, 127, -128, 127, 127, -128, 127, 127, -128, 127, -11, 127, -128, -80, 127, -128, -128, 127, 127, -128, 127, -128, -128, -34, 127, 127, -86, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -66, 127, 127, -128, 127, -128, 127, -128, -128, -24, 53, 127, -128, 127, -128, 127, -128, -128, 68, -128, -128, 127, 103, 127, 71, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -32, 127, -128, 95, -91, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -47, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 88, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 68, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -28, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 1, 127, -128, 15, 127, 127, 127, 127, -128, -128, -7, -128, 127, -128, -128, 6, -128, -128, -128, 127, -128, -128, 70, 17, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -44, -128, 127, -63, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 50, -128, -128, 127, 127, -128, -128, 127, -128, 78, -128, -87, 127, -128, 127, 60, -128, -128, -128, 127, -128, -59, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -81, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 117, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 53, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -2, 127, 127, -128, -128, 127, 127, 58, 127, -128, 127, -128, 127, 79, -128, 47, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -90, 127, 127, -128, -128, 127, -128, 127, -27, -128, 127, -128, -128, 127, -128, -128, 127, -128, 54, 127, -2, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 102, -50, 127, 127, 127, -128, 127, -128, 127, -128, 127, -74, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -97, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -22, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 31, -128, -128, -128, 76, -128, -128, -121, -128, -128, -128, 12, 127, -85, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -75, 127, -128, -128, 127, 127, -128, 127, 53, -128, 127, -128, -128, -128, -128, -128, -107, -128, 127, 127, 127, -128, 127, 127, 127, -97, 127, 101, -128, -128, 127, -128, -128, 121, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -124, 21, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -109, -128, 100, -128, 92, -128, 127, -128, -128, -36, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 69, -128, -50, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -50, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, -66, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 54, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -93, 127, 127, -128, -128, 127, -128, -128, 127, 103, 127, -128, -128, 127, 127, -128, -128, 127, -10, 127, 127, 78, 127, 127, 103, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 16, 0, 127, -128, -98, -128, -128, -128, -60, 24, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 63, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 49, 127, -128, 127, -128, -128, -128, -128, -29, 127, 127, -128, 127, 127, -128, -100, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -76, -128, 127, 127, -128, 127, -128, 127, -128, -119, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 8, 127, -128, -128, -87, 127, -128, 127, 127, -10, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 22, -128, 127, -128, 127, -128, -128, 127, 16, -128, -128, 127, 90, 127, -128, 53, 127, -128, -128, 127, 127, -128, 127, 127, 127, -8, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 45, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, -63, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 59, 127, 66, -128, 127, 127, -128, -128, 127, 127, 127, 127, 23, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 73, 127, 127, -128, -128, -128, -128, 127, 44, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -27, 127, -128, -52, -128, 127, -128, 127, -128, -48, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 31, 127, 127, -128, -128, 127, -128, 127, -128, -88, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -26, -128, 127, 127, 127, 127, 127, -8, 127, 127, 127, 127, 127, -128, 127, 127, -49, -128, 127, 127, -1, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, 53, 8, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -81, 127, 33, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -119, 127, 127, -128, -128, -128, 127, -36, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -102, -31, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 108, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -37, -128, 39, -7, -128, -128, 127, 127, -128, -128, 22, -128, -128, -128, 47, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 33, 127, -128, 127, 127, -128, 127, -128, -55, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -113, 127, 48, -128, 127, -128, -128, 127, 127, -128, -26, -128, -128, -128, 127, -128, 39, 24, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 74, -128, -128, 127, 127, -128, -73, 127, -128, -128, -128, 127, -128, -59, 127, -128, 127, 127, -128, -128, 127, 127, 127, -8, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 63, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 114, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 116, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 63, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -88, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 64, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -11, 127, 127, -128, 127, 127, 15, -128, 127, -128, -128, -128, -102, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 57, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 114, -128, -128, 127, -128, -128, -37, 127, -128, -128, 127, 55, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 50, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -96, 127, 127, -128, 106, 127, 127, -128, 127, 127, 127, -128, -128, 127, -95, 127, -2, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -119, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, 68, 127, -128, 127, -128, 127, 49, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -103, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 58, -128, 127, -128, 127, 127, -128, 127, 93, -128, 127, -128, 91, 127, -5, -128, -91, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 106, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 3, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -101, -128, 127, -128, -128, -128, 127, -128, -128, -128, -124, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 48, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 75, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 98, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 47, -128, 127, -128, -128, -128, -65, 127, 127, 127, -128, -128, -54, 127, 127, -128, -128, 127, -128, 127, -124, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, -39, -128, 127, -128, 127, -128, -128, -23, 127, -128, 127, -128, 127, -71, -122, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 49, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 74, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -45, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 34, 127, 127, -128, 127, 127, -10, 38, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -71, -128, 127, -119, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 53, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 92, 45, -128, 74, 127, 127, -128, 127, 42, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -33, 127, 103, -128, -128, 127, -128, 127, 127, 127, -64, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -81, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 114, 127, -128, 127, -128, 127, 127, -128, -128, 127, -5, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -81, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -68, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -2, -128, 127, -128, 127, -128, -106, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 0, -128, -128, -58, 55, -128, 127, 127, 127, 45, -128, -128, 127, 127, -128, 127, -96, -128, 127, -128, -128, 127, -128, -11, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -53, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -17, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 49, 127, -128, 127, 45, 127, 127, -128, 127, 127, 106, -128, -128, -49, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -34, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -17, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -7, 103, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -101, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -42, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 86, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -71, 127, -128, 127, 96, -15, 127, 127, 127, -128, 127, -128, 127, 127, -128, -22, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -102, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 12, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 26, -128, -128, 127, 15, 127, -128, 17, 127, -128, -128, 127, 127, -128, -128, -128, -128, -63, -128, 127, -128, -128, -128, 68, 127, -31, 127, -128, 127, 127, -128, 1, 127, -128, -128, -128, 54, 127, 127, 127, 58, 127, -128, -128, -128, 127, -128, -128, 127, -128, 79, 127, -128, 127, 88, -128, -128, 127, -128, -128, 127, 127, -47, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 114, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, -24, 127, -128, -128, 127, 127, -128, 127, 127, 101, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -50, -128, 127, 127, -128, -86, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 53, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 5, 127, 127, 127, 127, 127, 127, -3, 127, 127, 127, 127, 127, 127, -128, -128, 127, 34, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -60, 127, 127, -128, 127, -128, -128, -128, -24, 127, -128, 127, -128, 95, 119, 127, -128, -128, -128, -128, -118, 127, 44, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -2, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 13, -128, 127, 127, 39, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -103, 127, 6, 127, -128, 127, -3, -128, 52, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -90, 127, -128, -128, 68, 127, -128, -44, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -50, 127, -128, 127, 127, -114, 127, 127, 127, -128, -81, 127, -128, 127, 127, -128, -114, 127, 127, 127, 127, 127, 22, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 98, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -101, -128, 127, 127, 44, -128, 127, 127, -128, 127, 106, -128, 127, -128, 127, -128, -128, -65, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -24, 127, 127, -128, -24, 127, -128, 127, -128, -128, 127, 127, -44, 127, 127, -128, -128, 127, 127, -128, -78, 127, 43, -128, 127, -128, 108, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 32, 127, -128, 127, -128, -76, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 86, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 34, 127, 127, -128, -128, 127, -128, -128, 127, 127, -87, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -11, -128, -128, 127, -128, -128, -128, -128, -128, 6, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 55, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 98, 127, -128, 127, -128, 127, -128, 95, 127, -128, 74, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, -106, -128, 127, -128, -32, 127, 127, 127, 98, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -23, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 112, 127, -128, -128, 79, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 29, 127, -58, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 90, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -29, 127, 127, -128, 127, -128, -128, -128, -128, 88, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 13, 127, 127, -128, -128, 127, 80, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -13, 127, -101, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 101, 127, -128, 127, 127, 127, -128, -71, -128, -31, 86, -128, 127, 127, -128, 127, -128, 127, 102, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 101, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -113, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -81, -128, 127, 127, -128, 127, -128, -128, 127, -128, 118, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 76, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -22, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 33, 127, -128, 127, 127, -128, 127, -27, -128, 127, 127, 95, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -27, -128, 127, -128, 127, -128, -128, 127, 127, -128, 68, -128, -128, -128, -128, -128, -128, 127, -128, -22, 127, 68, 127, -128, 127, -128, -128, 127, -128, -78, -128, -128, -128, 127, -128, 127, 5, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 92, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -118, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 11, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -17, -128, 0, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -44, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 106, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 26, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -93, -128, 127, 127, -124, -128, -128, 127, 48, -128, 127, 127, -37, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -121, -7, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -74, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 98, -49, 127, 127, -12, 127, 8, -128, 127, 127, -27, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 33, -128, 11, 127, -128, 127, 127, -128, 127, 122, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, 44, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 112, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, 76, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -53, -128, -63, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -93, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 33, -128, 127, -128, 127, -128, -128, 127, 127, 86, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 21, -128, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 90, 127, 127, 127, -23, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -28, -128, -128, 127, -128, -128, 127, 127, -26, 127, -128, 122, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -15, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 43, 127, 127, -128, 127, 127, -128, 127, 127, -128, 78, 127, 127, -73, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 24, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 107, -101, -128, 3, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -93, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 52, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -2, -128, 127, 127, -128, 127, -128, -128, 37, 127, 127, -128, -128, 127, -128, -52, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 23, -128, 127, 127, -128, 127, -128, 127, 127, -128, -106, 127, -128, 127, -28, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 7, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 59, -128, 127, -128, 127, 127, -128, 127, -18, 127, -128, 127, 127, -128, 80, 127, -70, 127, 127, 127, 127, -128, 127, -128, 127, 127, -60, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 88, 127, -128, -57, -128, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 75, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 90, -128, -1, 127, 22, -128, -128, 127, 127, -128, 127, 127, 97, 127, -128, 127, 127, -128, 127, 124, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -54, -128, 127, 127, -128, -128, 107, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -106, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, -1, -128, 127, -34, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -69, -128, -128, -128, 127, 47, 127, 127, -23, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 11, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -124, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 16, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 12, 127, -128, -128, 127, -49, 127, -128, -71, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -123, 127, -128, -128, 127, 97, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -7, 127, 127, 127, -128, 127, -128, 60, 1, -128, 127, 127, -91, 127, 127, -128, 127, -128, 127, 127, 69, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -75, 127, -23, -128, -128, -45, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 23, -29, -128, 127, 127, -128, 127, -128, 127, 127, -128, -1, 127, -128, 127, -128, 80, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -92, 127, -128, -128, 127, 127, -128, -128, 127, 87, -128, 127, -128, -128, -102, -43, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -70, 127, -128 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
