-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            -7, 42, -6, 90, 86, -23, 27, 31, 77, 85, -67, 26, -109, 112     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -48, 88, 40, 0, -81, -67, 102, -108, -125, 40, 114, 53, -93, 56, -78, 26, -19, -128, -57, -113, -5, -61, -21, 117, 72, -82, 101, 65, -35, -113, 94, -95, -34, -42, -123, 64, -17, -26, 7, 7, 83, -76, 117, -63, 119, 60, 127, 2, -29, -81, -26, 91, -1, 5, 76, -112, -78, 116, 85, 74, -66, 63, -117, -19, -102, 60, 108, -66, 28, 0, 59, 127, 59, -8, 50, 31, 30, 30, 54, -106, 68, 42, -114, 83, -58, 25, -40, -61, 6, -81, 72, 12, -84, -128, -64, -9, -60, -93, 35, 52, 10, 1, 44, -123, 36, -27, 82, 20, 16, -37, 80, 98, 127, -69, -18, 47, 18, -87, -100, 115, -110, 32, 41, -99, 26, 98, -25, -26, 75, -19, 6, 110, -123, -43, -86, -45, -95, -6, -105, 75, 29, -69, -113, 57, -75, 97, 73, -71, -23, 85, 40, -49, -10, 81, 7, 74, 61, 126, -59, 3, 0, 75, -24, 41, 54, 39, -4, -113, 45, 95, 52, 16, -38, 4, -119, 82, 85, -33, -55, 17, -102, 42, 127, 26, 92, -17, 103, -45, -63, -15, 88, -90, 32, 18, 31, -65, -8, 27, -37, -101, 15, -62, 26, 18, -42, 79, -126, 95, -81, 81, -31, -93, 124, -3, -66, -37, 66, 35, 59, 94, 53, 89, -78, 118, -35, 32, 98, 109, -74, -23, 78, 85, 105, 93, 21, -99, -29, 64, -54, -90, -43, 35, -80, -53, -68, 31, -120, 37, -81, 77, 58, -65, 67, -14, -114, -37, -45, 4, -66, -98, 5, 67, -71, 51, 110, 42, 55, 78, 4, -123, -9, -94, -28, -58, -71, 56, 124, -25, -56, 71, -38, -40, 80, 102, -121, -23, 47, 5, 9, 25, -118, 118, -58, 25, 27, 37, -125, 85, -20, 90, 78, -49, 6, -107, -43, -113, 53, 50, -109, -11, 4, -5, 52, 17, -113, 70, 77, -8, -33, 86, 85, -41, -119, 26, -99, 55, 5, 30, -78, -2, 87, -117, 93, 55, 76, -88, -91, -70, -112, 2, -53, -108, -97, -95, -123, -90, 6, 83, -53, 94, 36, -121, -57, -41, -121, 58, -58, 108, 78, -101, 96, -51, -101, 13, 22, -57, 83, 46, -121, -91, 99, 41, 58, -51, -41, -117, 6, -6, 72, 46, 90, 108, 93, -72, 55, -102, -71, -4, 62, 79, 109, 55, 107, -21, 95, 76, -50, 106, -97, -42, 66, 44, -70, 13, -21, 61, 90, -80, -44, -14, -79, 66, -69, 14, 109, 112, -47, -52, 67, 100, -28, 0, 17, -43, 115, 117, 34, -57, 35, 69, -99, -40, 72, 92, 103, -74, 81, -42, 113, 37, 46, 113, -1, -50, 58, 0, -46, 119, -122, 3, -61, -38, -28, -128, 18, -58, -38, -117, 71, -10, -27, -122, 41, 41, 41, -77, -124, -104, 108, -126, -127, -95, -108, -88, 25, 60, -32, 119, 95, -64, -84, -67, 106, 90, 79, -61, -37, -99, -41, 72, 33, -4, -111, -38, -13, 82, -112, 53, 85, 98, 32, 41, 2, 2, -101, 116, -12, -86, -73, -38, -34, 99, 124, 52, -9, 60, -77, -16, -127, -56, -37, 17, -48, 63, -18, 17, -3, 85, -12, 77, 32, -16, 41, -11, -74, 39, -55, -25, -52, 70, -20, -40, -41, -109, -14, -127, -49, -42, -104, -23, 77, 100, 42, -17, 110, 58, -67, 94, -2, -84, -33, 75, -68, 25, -21, -44, 107, -66, 12, 33, -78, -127, -51, 92, 45, 74, 114, -93, 90, -50, 39, 91, 60, -69, -60, -64, -61, -13, -14, 76, 67, 117, 66, -34, -122, 41, 91, 67, -91, 46, 21, -126, 111, -7, -118, -11, -96, 22, -104, 77, -91, 82, -104, -89, 45, -81, 117, -51, -60, -21, 118, 59, 101, -120, 56, -114, -55, 38, -80, 17, 40, -15, 100, 31, -92, 59, 118, -101, -41, 110, 38, 80, -114, -39, -56, -101, -62, 23, 51, 66, -28, 101, -14, 96, -25, 94, -82, 109, 87, 87, -25, 84, -109, 25, 106, -70, -27, 25, -95, 32, -127, -111, -35, 10, -7, 47, 74, 28, -60, 39, 1, 92, -46, -90, 70, -100, -103, -118, 3, 106, 11, 110, 73, -24, 32, -117, 17, 75, 124, -106, -43, -74, -27, 13, -122, -127, -30, 91, -69, 3, -10, -6, -88, 32, -117, -3, 86, 13, 90, -79, -38, 6, -40, -17, 40, 124, -97, -9, 120, -106, 1, -70, -7, 27, 103, -93, 114, 82, -12, -77, 38, -89, 110, 38, 3, 19, 74, -98, 50, 55, -90, 51, -81, 7, -111, 106, -52, 9, 1, -20, -93, -75, -12, 77, -100, -99, 103, 118, -118, -123, 112, -92, -76, 67, -119, 15, -60, -50, -8, -115, 44, 33, 47, 35, -97, -60, -31, -40, -119, 39, 46, -45, -65, -5, 51, 18, 104, 21, 67, 95, 91, 93, 96, 75, 83, 26, -21, 44, -46, -54, -125, 78, 115, 13, -76, 43, 29, 34, -111, -4, 38, -5, 97, -36, -55, -104, -32, -11, -122, 53, 50, 7, -89, 103, 82, 113, -81, -5, 48, -40, -105, 107, 81, -51, -84, -35, -64, -93, -77, -91, 29, -36, 113, 22, -97, 36, -57, 23, 16, -63, 103, 21, 74, 36, 26, 50, 50, 117, -100, -18, -73, -72, 77, -81, 22, -23, -125, 97, 36, -27, 113, -8, -50, -90, -116, 70, 36, -47, -50, 15, 95, 79, 105, -3, -74, 23, -44, 92, -21, 59, 20, -114, -7, -10, -38, 27, -11, -108, -72, -20, 61, -112, -88, 82, 49, 2, -124, -76, 87, 15, 27, -1, -128, 68, 33, -47, -86, -126, -120, -48, -12, -113, 34, 22, 97, -82, 113, 101, 71, -61, 19, 34, 42, 70, -29, 113, -35, -15, 32, 64, 26, -51, 21, 110, -78, 46, 1, -79, -87, 1, 47, 1, -98, -48, 13, 52, -114, -34, -25, -78, 74, 95, -16, 21, 62, -61, -105, 68, 124, 41, -106, -49, 48, 88, -67, -73, 90, 67, 33, -91, -8, -26, 33, -6, 18, -67, 116, 65, -113, 36, -98, -20, -28, -23, 73, 101, 104, 74, 19, -2, 108, 26, -8, -61, -26, -76, 12, 50, 41, 94, 18, -52, 18, 14, -112, 50, 15, 31, -30, -77, 0, 28, 125, 51, -65, 15, 31, -55, 91, -103, -33, -104, -41, 57, 0, -123, 29, 42, 126, 105, -48, -3, 66, 126, -45, 115, 125, 29, 11, 47, 108, -104, -91, -126, -37, 62, -73, 92, -32, -37, -43, -124, -121, 55, -5, 75, 22, 88, -74, -16, -114, 98, 20, 81, 118, 28, 84, -18, -25, -46, -99, 21, -27, -49, -116, 108, -123, 47, -10, 88, -71, -77, 125, -96, -102, -72, 30, 78, -21, -71, 31, 43, -29, 2, 31, -64, 80, -113, -25, 87, -68, 84, 107, -76, -10, 55, 33, 50, 46, 87, 41, 57, -102, -87, 114, 98, 20, -118, -23, 121, 51, 31, 97, 89, -54, -40, 0, 14, 47, -114, -115, 54, -88, -1, -59, -109, 75, -48, 59, -46, 113, 27, -111, 3, 19, 12, 62, 86, 50, -128, -22, -9, -21, 104, -67, 77, 115, -92, -14, 48, -119, -1, 88, 115, -67, 0, -113, 50, 102, -82, 113, 115, -26, 108, -71, -125, 25, -45, -109, -109, -63, -118, -73, -9, 117, 90, -111, 24, -119, 110, -77, 79, 107, 30, -95, -85, -16, 7, -124, -76, 111, -81, -17, 105, 57, 69, -74, -71, -37, -21, -84, -24, 30, 16, -94, 69, 85, -80, 26, -12, 103, -84, 28, -28, 1, 98, 8, 7, 75, 102, 114, -9, 118, 94, 121, 84, -22, 106, 85, 107, 34, -104, -74, -9, -13, -120, -121, 6, 52, -118, 94, -7, 7, 121, 40, 40, 5, -9, -73, 101, -52, -60, 49, 43, 122, -6, -52, 97, -30, -53, 28, 13, -94, -9, -119, -80, 56, 72, 52, -125, -93, 112, 55, 102, -37, -84, 28, 33, -26, -85, 87, -92, -25, 72, 62, 31, -112, -114, -126, 27, 63, -58, -94, -92, -55, 14, 39, -22, -50, -34, 91, 2, 37, 119, 122, -89, -18, 21, -107, -127, 125, 53, -76, 85, -89, 27, -8, 123, -109, -90, -54, -79, -45, -89, -121, -58, 0, 104, 127, -7, 60, -119, 22, -32, 49, -10, -90, -85, 53, 40, 38, -116, 40, -34, -35, -82, -75, -13, -50, -55, 84, 123, -25, -15, -117, 101, 70, 74, -7, 115, 119, 67, 49, 11, -38, 14, -11, 47, -113, 22, 60, 46, 126, -12, 27, 99, 62, 54, 99, 75, -61, -3, 17, 116, -120, 65, -40, 37, -128, -25, -81, 80, -63, -70, -127, -71, 100, 53, 15, -53, -89, -30, -78, 122, -103, -124, 90, 57, 83, 9, 36, -9, 80, -54, 53, -33, -34, 97, 65, -99, 76, -2, 104, 101, -88, 100, 36, 70, -23, -118, -51, -100, 123, 47, 67, 64, 19, -53, -109, 97, 89, 7, 26, 9, 92, -104, -107, -37, 23, 61, 5, -16, -77, 85, 111, -10, 118, 7, -16, -33, -70, -24, 107, -28, -91, -12, 123, 9, -124, -52, 93, -75, 39, -11, -100, 121, -104, -103, 32, 83, 46, -37, 107, -20, -88, 11, 59, -30, 6, -7, 32, -23, 96, 27, 79, 105, -71, -58, 51, 3, -116, 35, -104, 121, 49, -8, 107, 68, -108, 5, 96, 64, 60, 120, 64, -20, 121, 85, -125, 19, 35, 46, -95, 17, -67, -72, 98, 25, -94, 92, -78, 73, -92, 92, -37, -80, 1, -67, 78, 80, 38, -40, 49, -48, 83, -103, -36, -98, 72, -98, 59, 45, -78, -108, -124, -28, 14, 103, 58, -5, 49, -71, -56, -90, 123, 47, 88, 66, 42, -107, 49, 5, 14, 76, -78, 70, 26, -2, 88, -103, 55, 34, 65, -102, -91, -60, 108, 73, -99, 64, -76, 74, -33, -36, 74, -90, 49, 86, 9, -37, 121, 99, 8, 7, 45, 28, 44, 103, 5, -92, 120, -54, -50, -14, 52, 71, 125, -98, 94, 61, 72, 85, 87, -1, 54, 0, 105, 67, 14, 106, -24, -33, 47, 45, -54, -102, 6, 114, -49, 33, 52, 32, -41, 69, 116, -25, 106, -16, 65, 27, -60, -33, 42, 29, -47, -112, 41, -98, -27, 101, 72, 121, 111, -53, 69, 64, 108, -78, 126, -105, -10, 76, 40, 102, 127, 115, -42, 118, 11, -118, 67, 52, -121, 60, 32, 22, 29, -7, -72, 9, 7, 64, 48, 119, 36, -122, -87, 26, -15, 107, -49, 100, 127, 51, 14, -14, -111, 18, -64, -20, -58, -32, -125, 92, 102, -102, 123, -42, -128, -122, 127, 44, -52, 74, 30, 25, -44, 96, 41, 45, 16, 104, 8, -115, -112, -118, -65, 43, -70, 65, 16, 111, -93, -123, 40, -118, -4, 99, 64, -117, 39, 61, 56, -29, 102, 0, 52, -72, -23, -26, 90, 75, -116, -99, 105, -20, 26, 63, 33, 20, -35, 49, 84, -43, -40, -93, 58, 16, -51, -27, -106, 64, 124, -15, 69, -24, 96, -96, -113, 52, 115, 10, -21, -116, -30, -64, 20, -84, -65, -109, -117, 61, 57, -32, 46, -103, 8, -9, 38, 13, -91, 82, 28, -8, -48, -112, -58, 5, 9, 113, 60, -23, 50, 8, -87, 3, 6, 25, 70, -26, 30, -30, 44, -71, 112, 71, 83, 9, -83, -88, 19, 89, 36, -123, -103, 102, 86, 74, -95, -30, 29, 104, 64, 38, 122, 31, 118, -123, 104, -88, 89, 30, 72, -74, -35, 63, -52, 122, -109, 2, 72, 42, -59, 98, 24, 82, 116, -103, -26, -115, 96, -14, -40, 22, 44, 82, 11, -99, -59, 47, 46, 65, -3, -75, 59, 56, -12, -86, -38, -95, 67, -114, 23, 13, 58, 113, -13, 35, 73, -100, 108, 83, 46, 123, 31, 77, -60, 70, -50, 26, -55, 65, 38, 12, 20, -122, -28, 43, -36, 73, 3, 30, 82, 115, -128, 25, 33, -10, 122, 124, -78, 127, 48, -27, 19, -43, 105, 90, 31, -32, 48, -60, 18, 71, 102, 31, 28, 19, 78, 75, 122, 117, -95, 29, 108, -91, -58, -77, 13, -118, -111, 32, -67, -49, 42, -28, -22, 25, 24, 35, -98, -18, -66, 102, 93, 48, 54, 64, 99, -7, 10, -18, -19, 117, -61, 63, 80, 20, 123, 12, -26, 124, 62, -64, -22, 72, 13, 94, 18, -117, 1, 90, -124, 50, 52, 106, -113, -110, -94, 91, 104, 108, -20, -51, -106, 18, -18, -62, 117, -63, 45, -8, -85, 78, 93, -84, 84, -24, -55, 38, 1, 53, -45, -110, -96, -11, 103, 28, 19, 36, 70, -24, -15, 117, 110, 95, 125, -8, 114, 37, 101, -96, 55, 58, -84, 94, -120, -118, 45, -17, 11, 82, 52, 40, 117, -62, -98, 2, 13, 125, 101, 85, 0, -114, -76, 59, 79, 109, -103, 9, 35, 3, -81, 33, 98, -53, -88, -75, 74, -115, -25, 29, 3, -31, 114, 108, -53, -27, -104, -56, -11, -64, 6, -105, 116, -24, 64, -98, -110, 71, 94, 79, -26, 42, 50, 15, 104, 21, 32, 116, 67, -120, -65, -46, -25, 70, -127, -54, 51, 80, -34, -8, -65, 83, 92, -9, -72, -126, -2, 104, 20, 53, -127, -20, -36, 16, 78, 25, -73, 115, -91, 110, -122, 86, 29, -17, -33, 90, -35, 82, 24, -20, 5, -72, 66, -92, -66, -9, -108, -32, 99, 101, -119, 26, -87, 75, 83, 54, -70, -14, 122, -23, -67, 121, 46, -5, -84, -128, -75, -52, 22, -21, -35, -1, 40, 71, -36, 91, 86, 6, 19, 22, 21, -54, 38, 87, 0, -128, -13, -102, 43, -99, -96, 28, 46, 36, -68, -114, -68, 21, 67, -121, 26, -30, -59, -97, 6, -4, 116, 8, -59, -105, 10, -50, -121, -60, -36, -95, 40, 33, 127, -29, 85, -61, 120, 105, -23, -43, 96, 99, 15, 39, 19, -60, -110, 2, -72, 23, -21, -35, -119, 4, -8, -35, 54, -126, -109, 47, 30, 56, -13, -20, -2, 32, 51, -118, -57, -112, 90, 92, -2, 29, 34, 68, 7, 50, -25, -98, 77, -106, 86, 76, -43, -85, 18, 87, 97, 8, -43, -70, -18, -106, -66, -25, -94, 8, 15, -92, 0, -108, 55, -11, -41, 22, -82, -24, 93, 23, 123, 114, 24, -118, 37, 39, -57, 95, 106, 82, 93, 32, 47, -8, 88, 5, -47, 36, 1, -10, -3, -49, 29, -49, 31, 102, -46, 72, -58, 4, -94, -45, 35, -115, -19, 34, 63, 103, -8, -82, 13, 91, 61, -105, -70, 115, 14, 43, -12, -24, -14, 56, 127, -115, 36, -20, 45, -50, -96, -102, -16, -96, 1, 72, 60, 54, -96, 61, -43, 42, 29, 86, 17, -12, 91, -20, 99, 72, -25, -101, -74, 94, -58, -117, 8, -81, -122, -15, -49, -9, 85, 29, -6, -84, -78, -22, -79, -49, -104, -87, 12, -122, 90, 106, 29, -43, -49, -108, -40, 28, 125, -93, 61, 68, -6, -67, -48, 53, -93, 5, -115, -120, 70, 22, -36, 33, -111, 17, 73, 49, 45, 103, 47, -73, 126, -120, 55, -83, 70, -59, 15, 107, -36, -100, -46, -64, 47, -124, 31, -96, 77, 3, -32, -73, -37, -30, 29, 36, -121, -10, -109, -81, -89, 2, 28, -73, -53, -36, 107, -50, 13, 50, 45, 118, 19, 111, 52, -106, 54, -103, -100, -18, 101, 75, -45, -97, 106, 61, 39, 109, 115, 80, 66, -2, 79, -5, 59, 82, -82, 30, -9, -52, 86, -9, -52, 14, 12, 55, -79, -113, 60, 19, -127, -107, -46, 126, -29, 102, -56, 68, 91, 72, 96, 45, 83, 92, 63, -110, -128, -55, -61, -19, -84, -71, -48, -127, -18, 62, 54, -96, 126, 110, -40, -56, -59, -86, -82, -104, 104, 69, -117, 19, 85, 85, -38, 84, 40, 0, -52, 98, -45, 57, 5, -86, 92, 90, -33, 93, 49, 14, 120, -111, 121, 42, -34, -79, 24, 108, -18, -29, 14, 67, 47, 125, 16, 44, 98, -88, -118, -122, -26, -28, -15, -43, 77, -48, 22, 120, -35, -9, 26, 40, 14, 11, -29, -51, 89, -101, -18, 49, 99, 6, 119, 43, -8, -85, -83, 126, -110, 42, 26, -123, -30, 37, -117, 47, -100, 14, 42, 99, -104, -106, 56, 60, 41, -23, 36, 21, 102, 49, -13, -110, -77, -72, 42, 73, 116, -5, -6, 95, -49, 25, 60, 22, -18, -60, -45, -118, -34, 53, -87, -111, 35, 95, -25, 19, 0, -81, 96, 4, -71, 86, 108, 30, 96, -32, -50, 48, 23, -64, 111, 109, -53, -109, 6, -12, -122, -71, 37, -108, 87, -58, -118, 89, -49, 101, 77, 43, -21, -76, -31, 84, 68, -71, -70, -87, -21, 119, 55, -5, -6, -81, 35, -90, 77, 84, 69, 3, 2, 118, -119, 74, -54, -33, -16, -92, 113, -44, -78, -86, 124, -100, 62, -10, -125, 127, -30, -27, -16, -24, -60, -116, -14, -108, -48, -50, -75, -80, -86, -63, 52, -73, 19, 23, 105, 88, -39, -41, -123, -85, -33, 18, -128, 94, 123, 11, 9, 78, 56, 17, -58, 1, 20, 62, 16, 9, 83, -121, 41, -95, -95, 85, -93, -127, -86, 114, 103, 69, -32, -6, -127, 24, 76, -51, -62, -11, 54, -81, 19, -128, 81, -115, 71, 110, -55, 100, 75, -95, -66, -102, -34, -20, -113, -57, -92, 123, -110, -31, -31, -20, -66, 39, 8, -41, 20, -82, -4, -94, -100, -64, 29, 86, -31, 87, 110, 72, 37, 88, -102, -40, 39, -91, 102, 94, 110, -102, 3, 124, 85, -47, 47, -10, 114, 49, -45, -77, -22, -53, -17, -12, -72, -124, 73, -35, -64, -29, -97, -7, 48, 59, 96, 75, -10, 1, -20, -72, 97, 92, -114, 114, -98, 50, 23, 32, -104, -103, -110, -108, 74, -92, -56, -49, -87, -28, 35, 62, -34, 104, -119, 119, 46, -58, -120, 36, -44, -2, -52, 87, -111, -54, 84, -54, 123, 123, -30, 64, 86, -92, -80, 21, -40, -115, 104, 47, 50, 126, -40, 41, -85, 37, 26, 44, -44, -8, -4, 120, -48, -9, 52, 46, -37, 38, -61, 25, -16, 42, -29, 43, 119, 54, 9, 31, -128, 10, -15, -119, -13, -17, 120, -72, -39, -128, -56, 46, -1, 46, -24, 64, 60, 10, -108, 68, 66, -110, 16, -61, 109, -31, 96, -117, 84, 79, -75, 37, -106, -29, -48, 47, -103, 100, -62, -12, 80, 18, 4, 10, -95, 35, 109, 2, -58, 123, -4, -11, 32, -7, -17, -117, 20, -8, 46, 119, 63, -106, 118, 104, -30, 68, -57, -91, 82, 53, 76, -84, -107, 72, -47, 112, 60, 90, 79, 126, -127, -50, 87, 92, -123, 5, -32, -50, -67, -108, -97, 90, -21, -59, 15, -11, -35, -9, 108, 15, 95, 117, 95, -47, 127, 63, 50, -103, -94, 35, 118, -8, 40, -108, 85, 14, -4, -73, 39, -44, -127, 58, 45, -103, 79, 20, -91, 35, 105, -32, -40, 44, -90, -12, 69, -114, 75, 57, -127, -83, -61, 63, -63, 40, 20, 85, 49, -32, -26, 38, 20, -73, 33, 127, 53, -77, 89, 69, 19, -51, -118, 84, -39, 83, 78, -14, -99, 26, -122, -104, -42, -74, -25, -40, 83, -51, -79, -112, 31, -76, 17, 18, 73, -33, 26, 70, -43, 15, 76, -84, 20, -41, -33, -35, -9, 123, -34, 12, -15, -71, 101, 70, 64, 53, 72, -13, 121, 101, -90, -85, 63, 110, 46, -127, -55, -96, -91, 10, 111, 3, 125, -97, -45, -117, -36, 95, -33, 118, 2, -57, -24, -113, 33, 92, -54, -83, -30, -33, 69, 17, 115, 76, -127, 89, -45, 91, -30, -13, 47, -94, 102, 39, -95, 11, -73, -126, -109, 84, 22, -59, 48, -46, -38, 22, 104, -7, -127, -39, 22, 56, -73, 109, -116, 102, 8, -3, 69, 29, 54, 43, 28, -80, -60, 50, 15, -128, 88, 13, 9, -105, 36, 74, -91, 101, -42, -58, 25, 87, 51, 47, 44, 107, 94, 74, -8, 4, 64, 109, 36, 97, -1, -103, -95, -109, -7, -26, -22, 7, 64, 49, 90, 118, 1, -105, 60, -88, -35, 110, 57, -74, -80, -10, -84, 124, -3, 106, 92, 46, -93, 118, 53, -87, 118, -19, -106, -96, 127, -57, 92, 124, -127, -74, -1, 33, -87, 95, -40, -23, -80, -76, -106, 94, 9, 78, 107, 99, 97, 26, -29, 73, -65, 59, -120, -111, 90, 58, -61, 38, 53, -35, -93, -22, -44, 102, -76, 10, -128, 73, 12, 74, -14, -1, -121, -17, 23, 4, -107, -71, -41, 62, -42, 53, 103, 79, -60, 91, 108, -101, -46, -54, -47, 12, -36, 90, 99, 1, 35, -112, 75, 44, 17, -83, 16, -101, 102, 81, 75, -2, 73, -1, -101, 33, -40, 73, 67, 71, -100, -126, 97, -46, -91, -105, 98, 119, 73, -18, 107, 21, -93, -106, -55, -10, 19, 49, 83, 70, 58, -2, -1, -62, 2, -26, -19, 96, -34, 20, -80, 40, -66, 61, -58, 119, 6, 75, 11, 5, -79, -122, 67, -61, -102, -35, 80, 85, -53, -54, 5, 21, 75, -113, 38, 77, -61, -25, -88, 17, -38, -18, 125, -55, 27, 33, -71, -119, -25, -13, 116, 49, -39, -100, -98, 40, 46, -64, -94, 26, -97, 51, -34, -52, -91, -99, 79, 84, 73, 19, -57, -102, 77, 39, -1, 59, 29, 117, 88, -25, -65, 21, -56, -86, 25, -9, -10, -49, -112, -29, 109, -111, 23, -115, 49, 94, -88, -33, 53, 8, -77, -13, -93, -31, 17, 19, -29, -90, 87, -74, -127, 19, 61, 69, -9, -109, 61, 0, -34, 27, 105, 7, 31, -13, -85, -94, -97, 33, 2, 69, -88, -80, 6, 69, 89, -114, 16, 95, 46, -59, -45, -86, 96, 4, 60, 85, 38, 78, -72, -20, 107, 68, 87, -92, -81, -28, -57, -7, -49, -106, 91, -118, 113, 53, -80, -89, -23, 63, -31, -58, -15, -51, -81, -75, 56, 25, 70, -122, 28, -83, -122, -121, 51, 102, 80, -19, -104, -115, 74, -10, -93, 91, 63, -49, -106, 97, 56, -123, -104, -88, -69, 38, 23, -90, -70, -14, 87, -75, 57, 67, 61, -23, 123, -18, 23, -16, 40, -29, -62, 32, -75, 15, 114, 102, 88, -97, -103, -68, 121, 79, 118, 7, -103, 94, 24, 14, 9, -55, -106, -81, 102, 115, 9, -10, -46, -47, -38, 86, -61, -55, 36, 104, 24, 87, 103, -108, -106, 42, 83, -86, -85, 122, -7, -44, -120, 10, -59, 40, -89, 125, -49, 47, -30, 70, 108, 77, 6, 44, -96, 65, -80, 6, 50, -65, -107, -46, 125, 107, 1, -88, -93, 64, 106, 80, -81, 69, -1, -125, -22, -20, 35, -98, 57, -120, 48, 4, -52, -4, -67, -21, 116, 28, -124, -85, 120, -103, -20, 72, 32, 35, -32, -63, 94, -96, 19, -18, -70, 76, 45, -76, -116, 103, 0, 65, 105, -3, -96, -117, -104, 31, 23, 26, -110, 59, -119, 99, 20, 2, 103, -45, -17, 44, 6, -10, -51, 28, -13, -56, 109, -53, 111, -101, 35, 32, -67, -47, -30, -121, -89, 13, -101, 80, 73, 118, 77, -119, 41, 102, -17, 30, -3, 112, -24, 82, -15, -42, 111, 110, -80, 40, 39, -115, -12, 5, 120, 127, 121, -110, 96, 67, 80, -80, 54, -57, -37, -109, -15, 32, -38, 14, 27, -101, 39, -126, -64, 94, -54, -119, 13, -31, 45, 34, 6, -10, 56, 69, -121, -97, -14, 83, -21, -95, -51, 32, 71, -53, -101, -16, 62, 41, -90, -51, -63, 19, 24, -94, 31, 93, -49, 12, -120, -116, 31, 113, 30, -12, 77, 42, 117, -2, 87, 26, -121, -85, 101, -74, -17, 17, -34, -110, 28, 39, -1, -11, -38, -78, 24, -53, 97, -35, 97, -90, 97, -126, -38, 36, -94, 107, 37, 103, 2, 85, -19, -73, -14, -12, -8, -40, 33, 78, -3, 103, -99, 106, 11, 109, -74, -40, -73, 29, 1, 66, -62, -16, -56, 44, 127, 121, -16, 118, -78, 76, 35, -41, -63, -76, -90, 122, -14, -61, -51, -60, -36, -105, -33, 75, 111, 40, 24, -107, -6, 53, 38, 9, -81, -120, 57, -92, 94, 39, 120, -34, -62, -45, 54, -79, 107, -68, 20, -127, 115, -91, 53, -16, 93, 6, -51, 99, 35, -20, 33, 79, -118, -75, -55, -44, -76, -119, -76, 22, 67, 95, -63, 70, -22, -6, -123, -88, -71, -102, 120, 100, -80, -110, 91, -116, 0, -112, 18, -68, -67, 112, 23, 127, -57, -121, -68, -115, 24, 64, -53, -25, -127, -38, 94, -21, -4, 46, -13, -56, -128, -9, 21, 53, 33, 98, -119, -10, -41, -12, -44, 14, 100, -14, -44, 58, -14, 54, 98, -78, 113, -119, 70, 69, -81, -19, -87, 9, 75, 32, 76, 53, 81, -120, -102, -14, 15, -6, -13, 64, -20, -105, -91, -90, 1, 113, -52, 126, -43, -62, 8, -39, -2, 71, 109, 124, 93, 57, 88, 4, 18, 36, -16, -117, -113, -41, 103, -53, 52, 28, 2, -22, 57, -114, -77, 52, -6, 124, -9, 96, 47, 37, 57, -28, -45, 24, -15, -19, -81, -69, 7, 76, -95, -98, -120, -4, 82, -92, 15, -55, -85, -83, -37, -122, -38, 95, 16, -101, 48, -21, -128, -76, 87, 43, -86, -56, 18, -42, -28, 110, -88, -9, -43, -25, 50, 65, -107, 45, -54, 67, 29, 96, 31, 49, -91, -12, 8, 18, -104, 57, 9, 59, -119, 66, 39, 30, 14, 55, -126, -6, -49, 2, 59, 127, 4, 117, -27, -112, -128, -114, 48, 57, 59, 111, -1, -70, 35, 65, 51, -125, -71, -77, 93, 2, 39, -3, 22, 76, 30, -37, 91, 13, -32, 77, 75, -102, -92, -35, 23, 49, 98, 15, 109, 84, 114, 87, 76, -38, -20, 15, -42, -74, 58, -82, 50, -85, -72, -100, 39, -113, 68, 106, -111, -22, 96, 89, -113, -51, 100, -92, 46, -74, -112, 83, 51, 107, 70, -112, -55, -49, 43, 101, -29, -67, 99, 80, -4, 98, 13, 32, 96, -50, -10, 125, -50, -7, 36, 46, 106, 104, -104, 72, 119, -82, 82, 0, -8, -5, 93, 94, 106, 81, 12, 13, 54, 78, -101, 7, -4, -100, -52, -103, 104, 77, -56, 21, 47, -93, -96, 68, 127, -68, 111, 75, -1, -89, -51, 21, -107, -55, -72, 70, 36, 32, -39, 54, -93, -59, 6, -63, 124, -29, 57, -87, 95, -78, -92, 3, -86, -21, 23, -16, -73, -110, 35, 43, 1, 116, 12, 118, 31, 69, 66, 62, 35, 110, -79, 52, 3, -44, -64, -57, -6, -89, -66, -124, 126, -3, -65, 72, 86, -50, -23, -46, 89, -84, -113, -27, -54, -60, -91, 72, 10, 126, 19, 113, 91, -126, 112, -51, -88, -64, 107, 120, 38, -84, 77, -72, -57, 111, -98, -56, 93, 13, -111, -95, -61, 111, 12, 91, 12, -30, 117, -98, -15, 102, -122, 91, 69, -62, -80, -30, -90, 118, -23, 29, 94, 21, -70, -27, -18, -33, 17, 102, -105, 59, -69, 33, -28, 43, 116, -99, -87, -51, 7, -18, -28, 20, 58, -9, 104, 86, 51, -30, -114, -15, 29, 84, -74, 54, -39, -99, 105, -75, -78, 93, 123, -126, -56, 2, 100, -45, -44, 96, 21, -74, -2, -91, 11, 79, -93, 121, 81, 66, 81, -85, 114, 50, 102, -95, 113, 24, -50, 64, -70, 92, 49, -98, 62, 27, 97, -23, 83, -13, 110, -85, 62, 31, 2, 55, -115, 114, 93, -77, 2, 57, -53, -28, -89, -70, 113, -104, 35, -66, 103, 94, -25, -5, 45, 32, -104, -74, 124, 5, -82, 61, -41, -64, -120, 1, 21, -70, 1, -86, -23, 27, 127, 38, 46, -57, 65, 0, -26, 80, 75, -83, 68, -112, -33, 120, 84, -50, -57, 58, 72, 17, -124, -83, -128, -108, -41, 73, -125, -88, 75, 70, 20, 84, 9, -12, -54, -106, 114, 1, -105, -106, -41, 0, -65, -118, -70, 88, 46, -104, -114, 65, -50, 87, 101, -65, -88, 85, 17, 103, 100, 48, 99, -15, -5, 55, -105, -120, 55, 76, -71, -125, 37, 49, -75, 25, -76, 97, -66, -108, -7, -118, 21, -1, 124, 70, 121, -36, -60, 99, 17, 99, 62, 110, -56, 78, -86, -78, -122, -120, -118, -75, 21, -43, 81, 39, 55, 62, -88, -34, 41, 126, -8, 108, 10, 71, -13, -116, 88, 20, 88, 75, -128, -4, -98, -97, -70, 25, -78, 119, 75, 14, -125, 25, 88, -74, -106, -21, -63, -118, -115, -76, 36, -105, 4, 28, -23, -12, 38, -19, -29, 86, -42, -3, 43, 77, 22, -104, -53, -16, 59, 33, 19, 66, 82, 127, 86, -23, -18, 65, 0, -26, 102, 97, -117, -4, -102, -31, 57, 73, 0, -18, 6, -101, -43, 110, 19, 32, -8, 25, -3, -33, -99, -67, -41, -81, 118, 54, 85, 62, 29, 111, -36, 30, -5, -113, 58, -6, -56, -104, -87, 30, 27, 27, -66, -119, -51, -119, -109, -65, 13, -114, 53, -27, -47, -75, -75, 96, -81, -77, -65, 83, -126, 114, 49, 81, 16, 65, 84, 116, -57, 9, 4, -47, -86, 116, -92, 73, 24, 13, 109, -121, 116, -76, -54, -77, 32, 119, 111, -111, 90, -30, -109, 52, 107, 110, -90, -36, -119, 70, -1, 84, 98, -86, 3, 113, -115, -79, 121, -3, 87, 40, -25, -37, 64, -70, 98, 81, 89, -72, -81, -16, -16, 75, 28, 67, 23, -66, 50, -28, -65, -66, -114, -14, -1, 95, -119, 41, -58, -58, 40, 105, 3, -7, -70, 39, -89, -100, -103, -98, 0, 6, -22, -108, 87, -53, 61, -60, 21, 100, -29, -99, -51, -51, 31, 34, -49, 15, -98, 97, -24, 103, 83, -65, -89, 5, 89, -52, 83, 121, -24, 55, -62, 29, 25, -124, 2, -79, -32, 73, -114, -81, 28, 36, -28, -112, -48, -65, -30, 90, -46, 66, -15, 110, -87, -88, -28, -43, 84, 83, -79, 113, 99, 84, 49, -14, 51, -67, -15, -91, -73, -7, 111, -25, 51, 38, 58, -60, -46, -30, 38, -67, 123, 31, 96, -107, 36, 48, 117, -59, -54, 53, 37, 103, 35, -38, -67, -105, -13, -21, 80, -36, 22, -48, -29, -27, 70, -77, -4, 68, -43, -12, 2, 117, -18, 65, -25, -2, 104, 88, -56, -3, -45, 33, -39, -124, -34, 116, 97, 44, 25, -33, -31, 91, -42, -85, 101, -6, 53, -77, 35, 39, -19, -88, 55, 120, -64, 30, -2, 20, -109, 52, 103, 2, 99, -96, -63, 4, -57, -74, -2, 55, -28, -25, 100, 88, -68, 24, 98, 76, 79, 73, 12, -108, 26, 101, 113, 1, 67, 46, -5, 86, -35, -67, -80, 67, -102, -2, 56, 32, -51, 48, -40, -40, -76, -14, 70, 5, -17, 105, 79, -9, 46, 98, -124, 17, -100, 72, 0, -126, 109, -58, -90, 88, 117, -61, 87, -99, 94, 49, 114, -63, 92, 54, 44, 125, 113, 115, 122, -38, -64, -58, -44, -116, 35, 54, 127, -15, 63, -117, -108, 13, 88, 116, -89, -33, -91, 69, 0, -41, 104, -60, 111, -66, -52, 25, 43, 26, 80, -120, 108, 84, 8, -61, -30, -58, -63, 4, 49, -34, -2, -39, -100, -63, 53, 94, -12, 50, -58, 55, -19, -53, -73, -16, -102, -97, 19, -52, -80, -52, 82, -103, 36, 34, 33, -83, 29, -3, -84, -89, 72, -103, -44, 102, 98, 108, 76, -50, -77, -68, 36, 39, -98, -20, -24, -97, -66, 67, -31, 11, -48, -27, -85, -96, 40, -80, 101, 85, 61, -100, -62, -23, -77, -102, -34, 99, 91, -74, 105, -74, -119, -13, 71, 1, 45, -55, -58, 104, 6, 39, -89, -14, -97, 126, 58, 58, -79, -56, -118, -86, -34, 123, -65, -7, 77, 94, -48, 67, 104, -126, 92, -41, -82, 13, 3, -53, 110, -99, -97, 54, 68, 95, -121, 0, -42, 87, 57, -24, -66, 119, 123, -27, -41, -76, 79, 66, -73, 20, 61, -112, -101, -25, -121, -25, -33, 37, -68, -102, -106, 71, -40, -39, 77, -51, -120, 43, 54, -107, 28, -37, 31, -13, 50, -81, -74, -50, 63, -70, -17, 124, -20, -124, 86, -45, 42, -58, -111, -21, 114, -102, -1, -29, -56, 106, -56, 35, 93, 61, -76, 24, -22, 93, -57, 50, 52, -66, 45, 116, -5, 62, -83, -117, 28, 100, -72, 107, 60, -37, -93, -88, 18, -30, -122, -73, -25, -62, 30, 115, 67, 123, 81, 15, -127, -7, 49, -7, 19, 75, 53, -5, 27, 52, 102, -122, 92, 18, -18, 43, 127, -90, -6, -13, 78, 4, 127, -11, -4, 63, 114, 43, 62, -88, -90, 63, -81, -62, 49, 56, 49, 50, -104, -55, 41, 36, 112, -112, 25, 127, -110, -101, -115, 122, -5, -66, 85, 81, -83, 44, 20, 115, 121, -91, 96, 10, 107, 122, -63, 122, -47, -97, -5, -16, 75, -89, 111, 41, -24, 83, 103, -44, -13, 63, -22, -22, 94, 7, 7, -105, -72, 78, -80, -1, -40, 113, -86, 34, 55, 99, -80, -87, 10, -61, 1, 35, 38, -91, -114, 14, -26, -104, -118, -43, -17, 31, -98, -12, 89, 70, -13, 89, 114, -121, 116, 75, -26, 83, 74, 120, 69, -88, -30, -123, -80, 56, 75, -43, -10, 0, 73, 58, -115, 16, -113, -13, -42, 32, 53, 102, 64, 57, -29, -56, -93, 97, 63, -45, 81, 61, 106, -21, 71, -48, 111, 40, -55, 3, -113, -61, 82, 54, -51, 23, -23, 84, -22, 89, -21, -125, 103, 4, 89, -70, -4, 28, -81, -101, -125, 85, 102, -14, -30, 3, -35, -48, 18, 52, 30, 5, -71, -72, 36, 9, -50, 15, 117, 85, -13, 62, -15, -113, -36, 39, 75, -51, -38, -30, 74, -52, -126, -71, -22, -93, 26, -69, -58, -100, -71, -104, -128, -30, 116, 99, -65, -122, -97, -85, -49, -51, 41, 48, 115, 43, -81, -66, -59, -33, 96, -20, -57, 26, -9, -114, 41, 33, -41, -23, -1, -121, 104, 40, -84, -81, -75, 98, -122, 112, -58, -36, -13, 87, 19, 59, -98, -37, -14, -128, -127, 12, -122, 86, 35, -45, -86, 99, -127, -55, 55, 79, 71, 120, 32, -42, -112, -32, 67, -81, -115, 52, 105, -117, -83, -121, 53, 68, -70, -30, -26, 61, 119, 126, -68, 55, -46, 79, -101, 113, 77, -34, -73, 37, 38, 72, -11, 6, 115, -48, 86, 107, -99, 54, 107, -20, 83, -75, 22, 108, 5, 94, -2, -69, -82, -100, -94, 96, -124, -16, 127, 113, -113, 80, 92, 114, -123, -7, -121, 64, -57, 79, -76, -33, 82, 81, 39, 76, -11, -46, 47, 126, -10, 110, 1, 20, -120, 30, -20, 50, 16, 86, 84, 81, 87, 71, 28, -79, 11, -96, -95, -86, -39, -31, 122, -73, 81, -98, -51, -23, 58, 16, -1, 9, -41, 81, 65, 63, -93, 60, -90, 53, -1, -57, 69, 93, 1, -16, 120, 13, 90, 23, 6, 7, 9, -5, 80, 25, 93, -103, 109, -84, 38, -33, -57, -74, 47, 82, -49, -97, -66, 10, -4, 115, 43, -85, 126, 98, 122, -38, -51, -17, -11, -85, -73, -57, -101, -97, -1, -61, -23, -114, -2, 63, -119, -64, -57, -92, 65, -103, -92, 1, -33, -98, -21, 67, -25, 35, -31, -15, -8, -121, -84, -68, -97, -122, -124, 36, 85, -89, 41, 97, 70, -77, 56, -9, -3, -63, 22, -27, -84, 28, -75, 109, 117, 106, 50, -49, 111, 39, -51, 38, -41, -114, -42, -32, -128, 46, 14, -26, 45, -48, 16, -56, -64, -88, 16, 82, 111, -12, 66, 26, -41, -6, -106, 51, 65, 120, -90, -42, 91, -38, -15, -108, 36, -50, -91, -82, 5, 113, -49, 98, 0, -105, 9, 7, 120, -48, 65, 49, -111, 18, 109, -69, -66, 83, -91, 7, -29, 64, 3, 78, 40, 120, 10, 49, -58, 66, 77, 30, -121, 90, -52, -12, 13, 118, 66, 109, 78, -40, -65, 43, 86, 86, -36, 125, -28, -116, 20, -63, -29, 19, -86, -40, 111, -58, 126, -113, 15, 37, 106, -36, 58, -72, -117, -26, 124, 3, 102, -56, 49, 116, -6, 32, -69, -28, -39, 19, 108, -7, 57, -2, -41, 20, -70, -127, -81, 90, -98, -98, -92, 32, 59, -88, -124, 125, 93, -63, 119, -54, 54, -88, 110, 60, -6, 72, -85, 53, 118, -55, -79, 124, -123, 95, -60, 37, 13, -113, 103, -83, -56, -123, 67, 35, 90, 33, 101, -28, 67, 84, -66, -2, 116, 50, 33, -75, 76, 40, 119, -89, 97, 11, 14, -12, -39, -57, -54, -74, -91, 33, 70, 55, -41, 102, -32, -114, 4, -58, 57, 53, 0, 70, -97, -54, -20, 108, -121, -9, 22, -91, -39, 109, -84, -105, 125, 112, -111, -98, 24, 30, 108, -85, 3, 54, 100, -73, 25, 99, 29, 36, 10, -3, 122, 8, 62, -46, -79, 92, -67, -47, 52, -56, -9, -76, 81, 0, -46, -38, -96, -47, -50, 97, -17, -34, -102, 63, 107, -50, -113, 126, -77, -50, 125, 82, -87, 7, 80, -27, -55, -123, 116, 84, 111, 47, 17, -67, -23, 73, -71, 62, 17, -111, 120, -16, -110, 43, 11, 39, 65, -45, -42, -59, -94, 81, 115, 55, 11, 73, -52, 45, -30, 127, 18, -2, -47, -90, -110, -127, -39, -123, -56, -21, -103, -57, -123, -12, -127, -80, -77, 73, 92, -60, -13, -68, -119, -60, -116, 48, -71, 24, -128, 83, 2, -7, 116, 105, -114, 89, -83, -121, 80, 43, -90, -25, 48, -124, -92, -16, 8, -12, 14, 92, -4, 107, 4, 81, -96, -4, -26, -110, 12, -47, 48, -30, 72, 8, -53, 40, 60, 7, 21, -26, -49, 46, 68, 66, -124, 36, -71, -125, -47, 52, 0, -1, 35, 76, 93, 38, 61, -43, -48, -71, -18, 127, -12, -102, 73, -29, 24, -114, -126, -2, 25, -12, 7, -126, -65, 44, -107, 46, 53, 127, 17, 84, -99, -106, -26, -56, 77, 59, -54, -94, 56, 93, -52, 25, 90, 25, -122, 57, 55, 112, -61, 64, 2, -92, -125, -103, 61, -81, -85, 78, 34, 24, -108, -7, -29, -107, -123, -24, 101, 102, -66, -93, -121, 27, -77, 118, 3, -36, 97, -122, -3, -35, 54, -63, -105, 86, 30, -105, 71, -12, 104, 45, -73, 40, -41, 95, 81, 3, -25, 68, 30, 91, -104, 74, -77, -4, 25, -66, 69, 87, -100, -103, 68, -37, 107, -10, 90, -84, -2, -104, -73, -46, 37, -28, 43, 25, 68, 17, -116, -24, 66, 37, -50, -99, 38, 23, 80, 54, -64, -39, -98, -70, 68, 69, -27, -36, 25, 20, -50, -51, 100, -36, -53, -32, -115, -101, 68, 73, -113, -30, 122, -48, -59, 12, 93, 83, 119, 68, 22, 120, 25, 120, 22, -117, -65, 29, 40, 126, -117, 13, -42, -110, -54, 82, 60, -41, 32, 126, -56, -62, -27, -25, -79, 39, 56, 93, -13, 60, -2, 27, 74, -16, 47, -127, -119, 89, 23, -52, -117, -61, -115, 111, -122, 71, 11, 1, 18, -53, 66, 8, 27, -119, 127, 56, 21, 35, -71, 117, -30, 94, 122, -52, 36, -67, 91, 45, -97, -51, 30, -102, -116, 32, -98, -37, 42, -86, 74, -43, -27, -86, -71, 97, -116, -20, -7, 73, -30, 81, 77, 114, -58, 104, 8, 119, -124, -126, 47, -39, 51, -33, -125, -12, 107, 29, -4, 41, -125, 28, -50, -79, -85, -57, -17, 84, -71, 106, -126, 90, -89, 51, 20, -18, 72, -76, -77, 38, 50, 16, -1, -48, 52, -42, -34, 103, -35, -76, -100, 97, 66, 98, 53, 98, -20, -95, 50, 76, -22, -1, 102, -56, 29, 79, 94, 5, -26, 15, -7, -86, 36, 96, 10, -97, -37, -76, -122, -110, 57, -54, -90, 76, 33, -126, 46, 111, -85, 10, 57, 6, 71, -88, 6, -88, -54, -113, 126, 64, -118, -87, -91, -120, 24, -8, 3, 117, 47, 39, -105, 63, 82, 115, 72, -74, 3, -32, -9, 96, 15, 98, -83, 113, -12, 73, 76, -115, -60, 39, 101, -25, 105, -65, -104, 10, 108, 11, -4, -38, 118, -57, -36, 54, -48, 44, -62, 23, 4, 111, 102, 123, -107, -117, 106, 51, 25, -105, -101, 54, 10, 105, 20, 13, 37, 8, -12, 52, 116, 25, 88, -91, 38, 42, 72, 94, -33, -15, -57, -64, -24, 121, -68, -117, -7, 46, -98, 78, -57, 72, 97, 43, 22, 121, 30, -118, 89, -54, 84, 52, -97, -106, 53, 96, 16, -125, -115, 0, -120, -72, -80, 6, 126, 62, 116, -115, -25, 55, 109, -103, 111, 80, -17, -64, 13, 31, -27, -91, -125, -54, -99, 3, -15, -25, 14, -99, -14, -98, -101, -2, -75, -32, 123, 122, 117, 4, -88, -57, 85, 20, 50, -40, 41, 47, -15, -112, -119, -83, -1, -23, 10, 66, -28, -60, -104, -8, 67, -108, -124, 104, 122, -43, 28, 103, 2, 81, -93, 54, 27, -9, 99, -125, -22, 119, 50, 27, 121, -56, -4, 88, 59, -42, -7, 38, 89, -41, 74, 123, -85, -61, -28, -127, -27, 41, 95, -15, 100, 124, 120, 102, -109, 126, 62, 19, -33, 77, -119, 8, 105, 122, 7, -51, 101, 64, -49, 18, 22, 10, -42, -39, 102, -39, 46, 0, -41, -77, 45, -48, -76, 77, 55, 56, -96, -119, -46, -82, 2, 11, -95, -100, -43, -23, -85, 102, 39, -73, 116, -111, -102, -53, 10, -120, -94, 80, 112, -103, 54, -88, -80, 36, -100, -34, -102, 97, 98, 84, -106, -10, 33, 82, 122, 78, -112, -9, 87, 90, 23, 71, 38, -40, -13, -25, -39, -42, 103, 6, 89, 33, -6, 110, -76, -48, -64, -2, -3, 31, 31, 98, 108, -44, -127, 39, -52, -5, -54, 76, -128, -97, -118, 105, -38, -22, -27, 43, 59, -15, 81, 72, -2, 30, -40, 4, -104, -33, -90, 7, 57, 46, 67, -93, 76, -120, -79, 68, -118, -1, -96, 86, 85, 58, -114, -10, -54, -70, -66, 96, 50, 107, -56, -1, 74, 42, -51, 87, -84, 4, -106, -64, -36, -14, 15, 64, -103, 61, -127, -96, 74, 73, 47, 78, 51, 40, 50, -1, 70, -107, -109, -51, -69, -123, 67, 90, 127, -35, -103, 64, -79, 115, 107, -98, 79, 55, 94, -50, -26, 86, -6, 51, -63, 33, 9, -121, -70, 42, -45, 74, -55, 98, -82, -64, -108, 42, -109, 48, 25, -66, -22, -42, 86, -125, -102, -87, -65, -34, -45, -90, -93, -32, -77, 0, 54, 90, 73, -29, -77, -103, 86, 110, -77, 61, 41, -68, -113, -102, 42, 120, -98, -27, 38, 98, -116, -64, -66, 125, 60, -60, 70, 47, -92, 104, 102, -124, 123, -45, -15, 100, 45, 116, 73, -123, 48, -48, -11, 30, 113, 127, -5, -87, -119, -57, 59, 88, 125, -127, -39, -96, -26, 59, 83, -128, 37, -82, -12, 12, -121, -64, 49, 26, -26, -61, 19, 49, -13, 14, -58, -36, -33, -65, -12, 47, 44, 85, -127, 46, -25, -109, 22, -29, 34, -70, 44, 127, 63, -15, 102, -40, -20, 7, -69, 22, -8, -128, 59, 57, -17, 77, -53, 125, 110, -103, -46, 95, 102, -12, -104, 24, 79, -17, 107, -60, 90, 110, 35, 25, -108, 57, 43, -104, -121, -107, 33, -103, -49, -23, -20, 48, 64, 60, 77, 50, -92, -82, -20, -22, 54, -127, 66, 110, -18, -81, -59, 25, 63, 56, 74, -8, 10, -54, -110, -23, 101, 19, -3, -16, -117, 16, 90, -105, 50, 79, -84, 123, 110, -123, -128, 31, -41, -18, -108, -100, 62, 10, 27, 96, -25, -93, -13, 29, -104, -31, -7, 33, 82, -117, -16, -124, -56, -125, 76, 86, 114, -61, -72, -128, 10, -94, 77, -92, -23, -31, -19, 17, 74, -74, -28, 11, -19, 117, 98, 30, -12, -128, -12, 51, -35, 79, 123, -111, 80, 4, -3, -77, -79, 12, -5, -78, 119, 86, 41, 22, -63, 49, 29, -80, -10, -48, -54, 71, -18, -97, -100, 123, -36, 35, 113, -79, -103, 28, -125, 56, 52, -1, -92, -7, -127, -36, -25, 124, 66, 27, 9, -9, -22, -36, 47, -76, 84, 118, -45, 43, -113, -28, 38, -52, 102, -44, -1, -113, 60, -28, 23, -51, 49, -86, 25, -38, 35, 54, 89, -16, -17, -110, -3, -62, 41, 33, 88, 109, 7, -49, -53, 82, 74, -55, 1, 84, -25, -101, -66, -109, 109, -117, -73, -58, 27, -124, 88, 107, 79, -24, -68, 44, -38, -71, 85, 38, -127, -54, 123, 7, 12, 49, 125, -13, -28, -18, 88, -58, -93, -81, -107, -75, 40, -29, 15, -108, 41, 121, 123, 4, -11, 85, 8, -124, -73, -79, 122, 44, 118, 33, -114, 3, -3, 62, 106, 23, -85, -14, 36, 4, -124, -18, -6, 24, -53, 17, -33, -7, -102, 78, -93, 76, 46, -72, -22, -38, 110, -97, -47, 73, -44, 108, -109, 41, 66, 50, -112, -104, 69, -54, -86, -61, -119, -120, -48, -21, 9, 108, -39, 82, 101, 48, 66, -1, -33, -10, -90, 72, 31, 85, -73, -107, 100, -58, -70, -23, 6, -61, 18, 4, -127, -113, 75, 119, -87, -13, -116, 38, -73, 84, -14, 50, -108, -84, 12, 46, -114, 106, -17, -29, 28, -124, -86, -29, -71, -37, 118, -28, -12, 120, -121, 74, -59, 37, 80, 74, -19, -41, -52, 4, 125, 61, -20, -75, 44, -96, -37, -101, 35, 44, -9, -117, -89, 5, -26, 0, 84, 86, 116, 117, -57, 46, -114, -2, -22, 64, 117, 52, -27, -111, 31, -62, -44, 113, 91, -11, -51, 36, -100, 92, -25, -35, -54, -24, -6, -54, -42, 110, 40, 110, 122, 32, -35, -62, -24, -12, 49, -100, -120, -97, -117, 6, -4, -40, -87, 9, -126, 69, -62, 30, -63, 80, -123, 84, -31, 127, -106, 52, -83, 125, -89, -41, -6, -71, -99, 77, 69, -60, -120, 110, 94, -81, -3, 42, 23, -103, -54, 115, 28, -64, 72, -53, 119, 118, 124, 54, 22, -39, 64, 86, 89, 125, -128, 47, -81, -111, -125, -68, -36, -28, 117, 32, -56, 6, 1, -8, 74, 91, -59, 86, 73, 32, -32, -86, -36, 26, -115, -91, 40, -24, -126, -16, -50, 26, -6, -72, -102, -76, -31, 36, -103, 109, -114, -41, 68, -107, -42, -110, 117, -27, -108, -108, 97, 63, -20, -74, -43, 86, 117, 4, -106, -44, -75, -116, 98, -63, -15, 65, -70, -4, -19, -5, -29, 28, -53, -50, -101, -72, -42, -83, 65, 78, 4, 103, -96, -9, -22, 81, 13, 121, -101, 2, -42, -73, -57, -44, 66, 83, -60, 15, -99, 31, -51, -40, -70, -113, 102, 19, 0, -38, 18, 77, 23, 67, 31, -111, 52, -52, -77, 52, 113, 121, 32, 110, 35, 95, -51, 72, 104, -77, 22, 48, 2, -4, 85, 108, -100, 45, 32, -32, 56, 15, -1, 62, 101, 100, 66, -29, 53, -105, 62, 29, 16, 87, -17, -120, -97, 52, 100, 88, 103, -15, 117, -100, 15, 56, -44, 38, 66, 47, 64, 64, -32, 15, 13, -48, 104, 3, -96, -88, -3, 91, -18, -20, 125, 101, -11, -7, -79, -39, -71, 110, 74, -34, -16, -10, 41, 18, 111, -24, 10, 35, -120, 34, 115, -1, 79, 4, 78, 2, 8, -48, -29, 46, 95, -105, 67, 30, -8, -66, 108, -9, -41, 85, -86, 99, -23, -69, -78, -40, -121, -29, 125, 10, 117, 45, -28, -23, 90, 122, -53, -118, -115, -10, 89, -19, 23, 42, -24, 78, -70, 47, 61, 95, -49, -14, 114, 88, -73, 89, -127, -71, -63, -59, 94, 69, -9, -102, 49, -99, 29, -113, -96, 120, 20, 126, 57, -77, 79, -23, -58, -48, -48, -56, 122, -55, 103, 70, -33, -127, -52, -14, 12, 15, -71, 108, -88, 9, 77, -33, 28, -25, -113, -68, 6, -86, -29, -51, 107, -36, 58, -96, -14, -39, -116, 28, -40, 83, 125, 74, -99, -81, 32, -10, -109, 119, 125, -114, 10, 20, -97, -64, 67, 25, 49, -59, -122, -83, 91, 43, -107, -70, 69, 92, -112, 60, 94, -19, -45, 91, 76, 88, -7, -6, -125, -23, 78, 86, 95, 9, -101, -86, 121, -120, 49, 66, 24, 13, -85, -29, 51, -21, -40, -79, -118, 127, 7, 21, -13, 41, 44, 43, -79, 4, -124, -121, 80, -15, 15, 8, 124, -101, 23, 21, 124, -67, 7, -41, -127, -70, -110, -13, -70, -3, -51, 12, -60, 55, -101, 28, -115, 23, 90, -31, 127, -88, -16, -108, 110, -62, 76, 122, -8, -62, 67, -70, 115, 118, -97, 12, -100, -86, 90, 50, 41, -124, -48, 100, -118, 7, 94, -8, 120, 63, -121, 83, 24, 30, -58, -121, -34, 35, -80, -19, 102, -40, -71, 50, 75, -39, 117, 61, 49, 97, 37, 98, -91, 47, -2, 39, -24, 109, 14, -96, -30, 109, 7, 62, -50, -56, -92, -77, 16, 74, 29, 36, 6, 30, -6, 72, 58, 82, -73, 19, -112, -112, -122, 81, -49, 95, 95, 103, 122, -55, -79, 57, 96, -9, 6, -62, -111, -42, 121, 77, 99, -75, -65, -117, -5, 59, 90, 22, 93, 10, -19, 2, 45, -29, -27, -32, -55, 51, 46, 125, -46, -61, 9, 101, -102, -21, 53, 77, 72, -5, -117, -122, -19, -109, 49, 46, -86, -73, 105, 37, -78, 100, -29, 43, 76, -3, -39, 95, 79, -15, 35, -54, -60, -52, -46, 82, 58, 84, -95, 28, -49, -68, 44, 82, -79, -87, 3, -116, -50, -70, -89, -11, -26, -62, -16, 35, 17, -121, -74, -73, 78, 79, 124, -78, 69, -60, 122, -84, 18, -20, -70, -104, 57, -52, -82, 118, -24, 119, -26, -54, -103, -32, 3, 69, 8, -16, 96, -10, -122, -38, -65, -45, 112, 68, -59, 117, 72, -57, 22, 96, -118, -125, 63, -18, -97, 48, -85, -31, -76, 100, -4, -117, -81, -28, -76, -121, 68, -14, -75, -64, 80, 36, -126, -83, 94, -28, 77, -107, -67, -24, -4, 64, -22, -34, -70, -45, 51, -24, 93, 14, 104, 109, 8, 80, -27, 107, -57, 99, 70, 91, 58, -93, 120, 51, 30, -8, 72, -80, 43, 97, -126, -13, -89, -16, -121, -98, -104, 35, 30, 8, 87, -64, 18, 21, -49, 15, -9, 91, -56, 47, -66, -44, 69, -111, 104, -96, -4, -109, -87, 113, -118, 44, 42, 107, -32, 90, -49, 107, -37, 77, -88, 41, -90, 110, -70, 22, -1, -121, -116, -117, 115, 38, -86, -48, 125, -10, -103, 7, -43, -7, -119, -74, 71, -11, 77, -32, -113, -65, -19, -21, 78, -114, -76, 91, -89, -104, -56, -102, 115, -58, 108, 29, 25, -111, 112, 75, 1, -55, 121, 55, 2, 51, -37, 25, 24, -21, 46, -13, -107, 76, 1, -76, -114, -95, -33, 103, 81, -7, -116, -98, -124, 82, -35, 99, -3, 105, 91, -90, 124, -88, -38, 96, -14, 72, 85, -104, -9, 86, 29, -88, -20, 83, 73, -104, 55, 32, 15, 5, -111, 47, 107, -82, 35, 57, -89, 2, -60, -96, -6, 119, 54, -30, 79, 35, -64, -4, -23, -121, -111, -122, 112, -33, 127, -89, 125, 82, -14, 93, -101, -69, -11, -45, 23, 32, -6, 24, 62, 110, 57, 10, -58, -41, 82, -57, 47, -38, 83, 109, -80, 93, 106, 5, 52, 75, 125, -42, -35, 70, 98, -125, 94, -54, -10, -98, -108, 89, -110, -85, -29, 17, 116, 18, -100, -7, 81, 14, -104, -66, 3, 68, 48, -91, 49, 76, 100, 22, -23, -22, 108, -34, 52, 41, 92, -17, -79, -80, -45, -29, -57, 101, 59, -63, 58, 55, 104, -76, -38, 6, 109, -45, 1, -6, -104, -107, -91, 67, 127, -59, 15, -82, 20, -8, 25, 64, 63, -20, -33, 4, 126, 63, -58, 12, -25, -1, 81, -128, 15, 104, 41, -87, -95, -47, 53, -25, -101, -22, -109, -24, 33, -82, 100, -120, -6, -6, -22, 25, 118, 58, 78, -37, -74, 118, 5, -123, 62, 88, 95, -9, 52, 111, -86, 71, 113, 46, 23, 120, 0, 38, -40, 22, -42, 79, -127, 18, 80, 43, -109, -15, 66, -117, 49, -72, -66, -25, 49, -125, 46, -116, 37, 90, 43, 93, 84, 33, -60, -97, 75, -10, -7, 58, 9, 11, -121, 103, -115, -47, -10, -51, -11, 127, -35, -73, -106, -102, 4, -8, 116, -6, 77, 111, -53, -64, -91, 27, 49, -49, 44, 118, 11, -23, -9, -128, 19, -79, 30, 57, -42, 19, 34, 98, 43, -79, -94, 2, -20, -37, 62, -68, 29, -71, -50, 57, 3, 13, -52, -2, -61, 125, -46, 52, -74, 35, -102, -102, -101, -4, -24, -71, -7, -76, 23, 90, 33, 78, -39, 69, 7, 89, -52, -105, -91, -45, -39, -47, 16, -94, 3, 74, 111, 9, -20, 108, -17, -85, -60, 100, -93, 119, -91, 116, 101, 58, 6, -39, -11, 84, 38, 32, 124, 41, 12, 29, 49, 12, 89, 37, -2, -71, -125, 16, -90, 117, 21, -17, 32, 98, 69, -33, -38, 122, 51, -85, 124, 66, 20, 46, 67, -3, -94, 106, -5, 112, -6, -28, 52, -90, -79, -76, 66, 42, -128, 96, 50, -86, -112, -6, 91, 103, -10, 7, 124, -62, 4, 22, 110, -89, -24, -34, -14, 107, 22, 70, -35, 34, -18, -64, 87, 73, 64, -122, -3, 107, -56, -88, 105, 67, -10, 105, -92, -90, -80, 63, -1, -80, 36, -69, 90, 126, 85, 40, 30, -118, -95, -56, 125, -80, 27, 39, 112, 13, -94, -40, 6, -27, -48, 92, 71, 31, -6, 39, -128, -18, -104, 43, 102, -35, 61, 23, -26, 115, 78, -89, -63, 90, -77, 9, 14, -60, 59, -1, -14, -66, 60, 54, -64, 107, 87, 3, -60, 122, 93, -114, 47, -60, 81, 61, 96, 92, 107, 30, 71, -125, 2, -48, 100, -68, -38, 126, -87, -126, -81, 0, -80, 34, 56, 17, -33, -89, -7, -74, 13, -118, -100, 32, -36, 11, -49, -19, -86, -5, -31, -117, 54, -62, -1, 57, -51, -72, 75, -106, 123, -90, -16, 83, -22, -108, 93, 21, -28, -97, 124, 79, 41, 65, -78, 1, -97, -51, 121, 27, 42, -124, 7, -46, -11, 35, 18, -30, -70, -109, -3, -119, -115, -19, 91, 127, 105, 90, 68, -32, -20, 8, -14, -99, 78, 57, -10, 0, -57, 42, 95, 76, 82, -102, -128, -124, -16, 25, 32, -83, 48, 63, -63, -79, -101, 44, 80, -54, 90, 87, -75, 46, -15, 107, 126, 4, -45, -56, 125, -57, 13, -9, -104, 75, -72, 59, 70, 28, -73, 31, -98, 96, -44, 123, 103, 117, 116, 9, 64, 3, -53, 24, 54, 62, -9, 84, -81, -42, -73, 58, 127, 78, 80, -31, -126, -62, -19, -72, 88, -54, -34, -26, -124, -85, 61, 17, -113, -9, 10, -35, -20, -89, -41, 8, 9, 54, 118, -102, -79, -39, 17, 20, 81, 44, -4, 85, -69, -77, 73, -84, 40, 121, -31, 88, -7, -3, 55, -13, 2, 22, -113, -53, -128, 23, 97, -23, 52, 120, -100, -96, -104, 16, 110, -77, 52, -103, 55, 124, 68, -34, 48, -68, 111, -86, -111, 86, -75, -37, -113, -67, -19, -122, 101, 25, -81, 19, -83, 79, -25, 18, -27, 57, 102, 57, 99, -57, 89, -120, -102, 14, -51, 36, 88, -96, -12, -17, 99, 1, -124, 123, -75, -27, -70, -125, 6, -18, 124, 12, 84, 5, 63, 74, 14, 43, -7, 103, 122, 53, -21, -7, 88, -101, 15, 23, -79, -25, 1, -59, -77, -2, -86, 31, 3, 109, -38, 126, -32, -50, -49, -106, -47, 39, -97, -42, -106, -31, 41, 114, -6, 64, -44, 24, -121, 15, 96, -72, -78, 14, -96, -36, 28, 54, 103, 124, 78, -8, -24, -20, -80, -70, 120, 82, -92, 88, -51, 6, 53, -79, -7, 88, -60, -84, -119, -10, 97, 13, -4, -57, 42, -63, 1, -66, -13, 2, -108, 112, -82, 112, -37, 97, -121, -1, -15, 111, -4, -118, 95, -124, 85, -27, 123, -34, -97, 12, -112, -27, -34, 76, -95, 2, 25, 96, -38, 22, -64, -108, 120, 1, 37, 52, 23, -92, 103, -123, -85, 124, -110, 17, -5, 38, 19, -80, -25, -101, 62, -105, -122, -30, -77, -122, -42, -20, -106, -66, 94, 81, -108, -50, -92, 70, -67, 78, 45, -19, -121, -51, 47, -91, 108, 31, 125, 124, -13, -86, 104, -1, 63, 58, -103, 27, -53, -90, -35, -39, -105, 100, 6, -70, -14, 112, 48, -3, -9, 29, 41, -36, -111, 75, 119, 5, -28, -39, -67, -90, -34, -88, -21, -26, 127, 98, -109, -71, -5, -123, 50, -91, -123, -78, 81, -115, 62, 62, 33, -43, 9, -51, 87, -37, 75, 117, -38, 5, 30, 126, 86, -103, -118, -116, 68, -80, 71, -118, 114, -114, -9, -11, 121, 30, 28, -88, -83, 93, -110, 86, 8, -4, 83, 86, 5, -28, 66, 40, 29, -78, 83, 57, -2, -2, 72, -42, -6, -13, -40, -90, -48, 94, -51, -128, 43, 36, 97, -111, 83, 116, -46, 88, -72, 72, -20, 61, -125, 40, -98, -55, -9, 120, 101, -35, -93, -9, 40, 94, 106, -18, 6, 110, -30, 78, -26, 55, 16, -40, 124, 110, 125, 57, -117, 9, -81, -13, 47, 2, -50, -2, -88, 25, 33, -126, 28, -21, 53, -29, -85, -67, 18, -118, -7, 10, 27, -128, -12, -13, -91, 126, 54, 46, 72, -12, 71, 112, 36, -6, -112, -45, 77, -4, -61, 71, -33, 106, 115, -40, -78, -1, 109, 65, -126, -62, -45, -32, -61, -65, 44, -99, 4, -117, 25, -116, -125, -114, -22, 97, -4, -13, 36, 54, -9, 125, 38, -100, 102, 92, -116, 18, 79, -81, 44, 117, 10, 116, -75, -83, -90, 105, -49, -44, -124, 104, 110, 76, -71, -120, -54, -104, -94, -66, 50, 66, -51, -9, 90, 53, -94, 92, 121, 20, 102, 107, -46, 53, 6, 22, -104, -78, 5, -77, -117, 60, -77, 105, -114, 79, -95, -75, -49, -87, 99, -35, 54, -13, -16, 37, -127, 17, 17, -96, -2, -106, 27, 87, -116, -72, -68, -23, 53, -88, 40, -33, 127, 63, -23, -70, -105, -71, 48, 122, -24, -64, 76, -56, -80, -32, 30, 5, -36, -56, 12, 96, 77, 40, -72, -69, -10, -14, -26, 22, 89, -121, -65, -57, 123, 117, -90, 58, 8, 28, -39, 0, -56, 66, 0, 71, -18, 118, 60, -63, 24, -125, -8, 24, 126, 88, -1, -11, 63, 121, 2, 87, -91, -15, 115, 61, 102, 60, 64, 27, 116, -115, -7, -44, 28, -55, 83, -24, 3, -33, -28, 62, 73, -83, 0, 76, -64, -123, 88, 4, 118, 35, -39, -2, -118, -108, -126, -125, -69, 41, -61, -7, -66, 73, 104, 15, -6, -66, -32, -53, -40, -112, 34, -11, -74, -15, -119, -43, 62, 107, 25, 43, -64, -73, 53, -72, 95, -124, 33, 123, -30, -71, 62, -9, 126, 104, 63, 104, 78, 73, -6, -30, -66, -109, -22, -70, -61, 37, -111, -72, 86, -57, -30, 43, -93, -83, -127, -17, -97, -40, -29, -84, 125, 104, 112, 5, 81, -14, 101, 99, -106, 17, 90, -114, 83, 34, 123, -52, 126, -30, 83, 81, 54, 51, 32, -32, -18, 57, -112, -93, -14, 124, 42, 46, 95, -19, -23, -23, -86, -17, 64, 114, -127, -66, -65, -15, 49, 83, 10, 81, -85, 91, -105, 58, 111, -61, -85, -122, 22, 28, 53, -41, -30, -65, -74, 78, 116, 74, 70, -120, -113, -37, -15, 18, 48, 116, -111, 23, 35, 79, 113, -22, -15, -33, 64, -36, 43, 106, 1, 86, 24, -63, -88, 27, 86, -93, -84, -87, 81, 69, 111, 111, 67, 64, -92, -117, 47, -10, -34, 54, -91, 35, -34, 124, 100, 62, 0, 73, 107, -13, 122, 14, -65, -14, 33, 77, 63, -83, 11, -46, -17, -6, -104, 4, -54, -25, -6, 92, -114, 55, -60, 10, -125, 89, -84, 91, 115, -78, -81, 28, -115, -67, 55, 40, 44, -83, 10, -9, 83, -128, 111, -120, 89, -93, -27, -95, -45, -85, 98, -82, 19, -71, 114, -70, 106, -79, -38, 120, 111, -108, -108, 37, 77, 63, 121, -61, -111, -83, -46, -24, -112, -113, -2, -97, -3, 46, -119, 112, -22, -84, 85, 81, -82, -95, -49, -71, -58, -11, -30, 98, -105, -121, 94, -111, -7, -8, 37, -68, 46, -63, -23, 57, -91, -1, 76, 60, -19, 126, -63, -103, -32, -7, 57, -72, 46, -93, -6, 12, 4, 75, 119, 30, 81, -14, 28, 75, -12, -95, 94, 56, 38, -17, 88, -117, -43, -116, 29, -122, 30, -96, 85, -91, -70, 39, 116, 78, 21, 44, 81, -42, 71, -102, -37, -115, -111, -10, -87, -37, 31, -109, -109, 10, -101, -37, -23, 92, 79, 4, -4, -96, 64, 22, -96, 5, -86, -40, 1, 6, -122, 95, -6, -98, 14, -12, -95, 20, 68, -62, 81, 49, 4, -50, 36, -10, -74, -1, -68, -110, 42, -93, 2, -58, -76, -70, 74, -112, -70, -41, 24, 80, -126, 77, 73, 68, 85, -2, -3, 13, 48, -13, -106, -117, 92, -99, -37, 56, 37, -59, -3, -30, 7, 64, -11, -12, 63, -117, -42, 126, -75, -109, 115, -107, 100, -49, -114, 43, 21, -72, -29, 119, 81, -66, 62, -2, 19, 99, 100, 21, 10, 99, -64, 111, -78, 46, 24, -106, 25, 70, 3, -97, -31, -125, -44, 103, -22, 19, -107, -50, 55, -92, -109, 49, 31, -89, -110, -67, 119, -9, 86, -69, 77, -99, -16, -95, 27, 71, 41, 77, -116, 16, 84, -63, 21, 112, 110, 112, -51, -69, -44, 71, -52, -17, -127, -64, -65, -13, -122, 108, 27, -68, 95, -4, 38, -109, 49, -57, -51, 32, -22, -10, -20, -14, 91, -69, -115, 125, -45, 2, -23, -89, 87, 95, -80, 61, 79, -21, 39, -122, 0, -89, -18, -117, 59, -46, 96, 71, -53, -92, 95, -47, -113, 89, -119, -109, 1, 10, 101, -99, -59, 112, -31, -46, 102, 11, 60, -119, 55, 30, -113, 74, -14, -46, 19, -72, 32, 37, 71, 17, -16, 42, 15, -1, -31, -126, -38, 71, 110, 81, 69, 88, -24, -102, -30, 58, -53, 58, -123, 96, -79, 104, 99, 62, 8, 32, -93, 14, 63, -74, -125, -56, -114, 71, 58, 25, -97, -28, 62, 119, -11, 30, 35, 107, -113, -43, -126, -50, -121, -44, 96, -46, -24, 100, 66, 40, -78, 111, -63, -108, -48, -3, 29, 24, -84, 57, 113, 22, 111, -87, 117, 65, -32, -104, -21, -21, -59, 68, -78, 98, -112, -13, 17, 67, 72, -87, 21, -100, 99, -32, 12, -77, -67, -33, -96, 33, -39, 7, -94, -96, -40, -5, -21, -36, -39, -53, 47, 7, -46, -9, -52, 78, 99, -27, -75, 33, 60, 108, -64, 38, 6, 34, 74, -40, 71, 51, -111, -111, 4, 81, -104, 98, -98, 70, -32, -51, -88, -8, -78, -50, -56, -6, 85, -122, 109, -113, 87, 11, -128, -21, -69, -118, -30, -123, -40, -69, -57, 53, 80, -79, -116, 96, -109, -59, 16, -19, -61, -101, -87, 4, -57, 66, 110, -14, 13, -41, -62, -56, -52, -105, 127, 76, -90, -28, 22, -128, -49, -107, 67, -89, -41, 63, 75, -114, -22, -87, -82, -89, -16, 109, 115, 4, -115, -46, 57, -57, -106, -91, -105, -111, -87, -44, 46, 105, -53, -48, -4, -48, -48, 28, 62, -32, -56, 78, 124, -58, 115, -42, -28, -21, -91, 109, 31, 101, 0, 116, -119, -94, 125, 16, -123, -69, 45, 9, 19, 123, -42, -98, 55, 71, -49, 76, 3, 16, 6, 104, -119, 111, -95, 21, -93, 123, -5, 17, -94, -124, -13, 72, -114, -75, -30, 63, 77, -32, 98, 64, -77, -29, 109, -101, 57, -57, -7, -83, 104, 71, 120, -15, 74, -81, -22, -25, 125, -93, -128, -93, 4, -61, 71, -7, -123, 28, 76, -19, 90, -118, 42, 64, -44, 96, 78, -14, 109, 91, -36, -61, -97, 66, 23, -114, 22, 8, -33, -24, -125, -46, -76, 55, 105, -21, 120, 75, 80, 96, -43, 15, 31, 87, -44, -119, 74, -20, -26, -16, -79, -119, -100, 116, 45, -7, 41, -30, -1, 12, 5, 10, 64, 14, 78, 84, -29, 52, -109, -99, 36, 89, -33, -93, -62, -115, 2, -81, -108, -72, 12, -71, 28, -125, -104, 30, -41, -23, 51, 6, -1, 21, 53, -61, 118, 19, 20, -78, -128, -20, 121, -42, -101, -3, -112, 34, 83, 47, -87, 113, -89, 97, -42, 122, -9, -96, 76, -121, -17, -1, -75, 24, 50, -19, -100, -34, -56, 78, 97, 93, -95, -24, 93, 21, -127, 31, -72, -31, -127, -42, -17, -94, -25, 11, -13, -17, 62, 8, 27, 3, -106, -74, -106, 23, 63, -8, -70, 36, -127, 100, 5, -43, -41, -32, 115, -94, 0, -57, 41, -104, 38, 55, -32, -47, -53, 34, -21, -82, -88, -97, -70, 51, 35, -13, 65, 66, -127, -126, -65, 68, -27, -89, -114, -14, -38, 125, 115, 32, -82, 68, 113, 109, 2, 53, -83, -120, 54, 60, -70, -29, 63, -64, -111, -23, 20, 39, -110, -105, 99, -19, 87, -93, 22, 24, 14, -116, 44, -56, -52, 24, 19, -78, -45, 4, -100, 122, -35, 11, -90, 15, 34, -111, -68, 13, -49, -4, 79, 42, 4, 122, -95, 24, -71, 100, 98, 89, -28, -113, 9, -19, -39, -77, -50, -51, -3, 4, -47, -86, 127, -4, -108, -104, -9, -45, -104, -47, -116, -35, 0, 50, -54, -53, 23, 115, -16, 84, 81, -54, -68, 79, -6, -121, 9, -72, -56, -34, -37, -92, -122, -7, 91, 62, 104, 42, -108, -116, 102, -84, 68, -86, 45, 44, 35, -41, -106, -117, -1, 120, 34, 54, 78, -45, -40, -74, 117, -88, -28, -64, 78, 106, 52, -59, 117, 36, -28, -87, 35, 80, -75, 56, -63, -46, -66, 103, 87, -83, 11, 28, -33, -34, 104, 119, 10, -26, 18, 126, 127, -92, 78, -119, 125, -36, 15, 65, -54, 86, 70, -66, 69, 112, -68, -8, 4, 75, -68, -48, -11, 106, 24, -32, -44, 9, 95, 10, -40, -58, 127, -126, 37, 29, 65, 32, 1, -18, 71, 85, -103, -16, 32, 23, -123, 87, 95, 108, -124, 66, 108, 13, -30, 82, 105, 82, 69, 53, -109, 77, 16, 45, -54, 95, -38, 108, -53, -49, 54, -106, 54, 71, -61, 114, -49, 70, -28, -79, 103, 104, -67, 46, -59, 77, -66, 9, -116, 88, 4, 127, 46, 60, -68, -62, 48, -10, 104, -51, -74, -108, 30, -73, -30, 66, 48, 33, -113, -90, 79, 88, -8, 2, -71, 38, 31, 71, -15, 100, -42, 10, 34, -37, 7, -48, -45, -41, 60, 35, 102, 62, 121, 116, 13, -67, -5, -51, -9, -28, -41, -116, 42, -96, 86, 76, -95, -102, -29, -106, -101, 67, 18, 32, 22, -128, 74, 16, -4, 30, 61, -5, 61, -74, -28, 2, 111, 82, -78, -103, 56, 102, -60, -108, -67, 126, 27, 127, 21, -110, 69, -26, 74, 110, 71, -8, 27, 36, -93, 22, 122, 41, -116, -30, -78, 59, 75, -62, -83, -110, 53, 38, -31, 47, 110, -2, -72, 120, 124, -70, 108, -108, 73, -111, -58, -74, -18, 104, 38, 58, -48, 45, -12, 11, -60, -126, -31, 121, 84, 113, 94, -18, 78, -125, -109, 121, -119, -15, 124, 22, -92, 70, 61, -3, -44, -114, -113, 25, 78, -127, -122, -61, -77, 122, 86, 60, 45, -53, -40, 66, -70, -128, -126, -77, 66, -12, 77, 30, -10, 60, 3, -123, 87, 55, 55, -63, 83, -46, 39, 30, 39, 92, -63, -72, -111, 127, 103, 87, -94, -128, -42, -28, -44, 64, -20, 59, -75, -104, 37, 4, 33, -98, -91, 21, 75, 34, 0, 111, -70, -66, -65, -37, -11, 96, -113, -22, 119, -56, -33, -3, 113, 62, 65, 73, -40, 103, -63, -59, 103, -12, 51, -53, -60, -123, -19, 49, 28, 27, 7, -113, 113, -74, -112, -32, -121, -109, 47, -57, 29, -112, -96, -88, 18, -104, 55, 115, -28, 127, -98, -58, 124, 62, 32, -59, -72, -116, -61, 5, -73, -8, 38, -8, -64, 111, 123, 5, 52, 48, -36, -65, -44, -16, -100, -70, 107, -6, -4, 2, 106, 9, 41, 21, 104, -38, 42, -57, -92, 43, -5, -118, -61, -80, 67, 73, -29, 71, 123, 7, 103, 1, 110, -81, 52, -14, -21, -77, -126, -52, -32, -45, -35, 40, 103, -51, -35, -15, 100, -38, -16, 120, -98, -122, 80, 76, 122, 45, 20, -30, 15, 119, -96, -47, -118, 85, 94, 23, -86, 56, 5, -16, -21, -126, 9, -57, -45, 49, 124, -78, -75, 1, 66, -16, -30, -86, -125, 60, -70, -2, -20, 39, 20, -37, 97, -47, -76, -99, -105, -127, 83, 46, -15, 115, 42, -34, -65, -35, 88, -74, -59, 27, -50, -67, -89, -100, -97, -97, 33, -8, -101, 40, 56, -56, 47, 125, -48, 113, 104, -35, -60, -1, -19, -34, 14, 115, 94, 47, -20, 7, -105, 33, 17, -73, 60, 32, -10, 32, -93, -74, -13, 109, 45, 33, 70, -100, 59, -52, 46, -15, 44, -17, -112, 66, 91, 15, 39, -65, 88, -57, -82, 20, 75, 69, 105, 43, 49, 107, 79, -31, -97, 17, -63, -60, 49, 83, 66, -42, -103, 64, 29, -39, -101, 89, -9, -119, -72, 27, 16, 100, 15, -98, -17, 62, -48, -59, 86, 9, -81, 17, -65, 7, 86, -49, -3, 126, 125, -58, 126, -38, -51, -80, -34, -76, 78, 9, -18, 49, -4, 124, 125, 46, -8, 40, -48, -11, -43, 35, 96, 28, -19, -90, -85, -54, -51, -105, 34, -45, -5, 112, 82, 36, -76, 69, -72, 27, 28, 31, 85, -23, -55, 106, -123, 59, -56, 109, 97, 39, -17, 91, -53, -43, -102, 84, 122, -62, 81, -56, 48, -75, 100, -75, -34, -30, -96, -33, -85, -19, -30, -75, 39, 93, -93, -111, -45, 94, 30, -49, 22, 41, -126, -51, 40, 86, 108, 74, 73, 117, -92, 59, -20, -67, 35, -69, 19, 8, -73, -77, -93, -124, 89, -19, -61, 38, 98, 77, -11, 95, -60, 106, 85, -53, 57, -68, -91, 117, -95, 84, -1, -33, -63, -80, 53, -56, -43, 56, 119, 65, 90, 75, 69, 6, -56, -83, -27, 97, -120, -41, -108, 21, -100, -9, -17, 50, -7, 15, 14, -101, -62, 82, 46, -90, 105, -80, 58, -86, 51, 82, -105, 31, -69, -123, -36, -112, -62, -55, 20, -39, 39, 28, -109, -37, 97, 80, -30, -56, -101, -20, -105, 10, 20, 44, 0, -18, 56, 72, -40, -38, -69, 24, -8, -82, 82, 26, -74, 56, 71, -117, -17, -112, -25, 106, 112, 89, 92, 110, -16, -93, 53, 83, -94, 39, 44, -39, 89, -97, 88, 51, 91, 79, -23, 17, 88, 70, -106, 123, -44, 10, 53, 52, 35, 90, 19, 125, 68, 35, -127, -1, 59, -42, 77, -113, 95, -27, -85, -97, -114, -5, 30, -42, 94, -36, 90, 32, 109, -50, 62, 77, -42, 12, 100, 111, 31, 17, -25, -108, 14, 6, -40, 5, 14, 114, 37, 27, 0, -90, 63, -89, -108, -10, 6, -37, -66, -123, -13, -64, 1, -15, 42, 33, 43, 42, -77, 94, -58, 121, -86, -112, -90, 3, 24, -62, -128, 89, -110, -37, -32, -109, 117, -18, -126, -37, 112, 44, -104, -128, 95, -80, 54, 94, -52, 117, -93, -31, 89, 27, 106, 3, -84, 71, -88, 13, 126, -103, -59, -17, -62, -93, 52, 18, 127, -39, 8, 33, 127, -107, 68, 52, 26, -47, 117, 116, 70, 85, -35, -29, 85, -94, 89, -47, -56, 67, -78, 40, 91, -122, 80, 8, -42, -119, -59, -77, -65, 50, 123, -105, -105, -63, -54, 119, 6, 113, 109, -118, -39, 89, -104, 118, -75, -70, -18, -67, -37, 61, -65, -14, -30, -89, -29, 9, 91, -103, -108, 78, -2, -49, 43, -65, -99, -110, -123, 114, -110, 84, 53, -24, 23, 2, 68, 6, -44, 100, -11, 1, -55, 52, -99, 60, 43, 38, -6, 84, -57, 105, -86, 4, 35, -111, 21, -112, -63, 111, 90, -68, -32, 71, 87, 91, -49, -17, 75, 42, 46, 68, -128, -101, 44, 67, 12, -103, 100, -41, -73, -36, -87, -101, 103, -33, 121, 114, -7, 89, -94, -124, -15, 25, 78, -20, -111, -8, -58, -95, -90, 118, -69, -29, 76, -31, -105, 82, -2, -65, -51, 39, -113, 90, -105, -10, -42, -39, 19, 80, -77, 18, 25, 70, 42, 123, -117, 32, 81, -56, -125, -17, -40, -6, -51, -65, -47, -109, -55, 77, -36, 61, 104, -63, 101, 115, -51, 47, -109, -76, -15, -53, -23, -104, -16, -57, 17, 59, -126, 19, -61, 81, 59, -17, 21, 99, 26, 38, -85, 115, 122, -49, 116, -96, 18, -9, 21, -40, -80, -106, -113, -25, -1, -54, 17, 2, -35, -53, 118, 24, 71, -73, -29, -71, -89, 17, 94, 87, 6, 76, 20, -66, 84, -108, 52, 11, 67, -101, 69, -127, -120, 8, -71, 51, 2, 125, 6, -6, 53, -25, 32, 51, 119, 60, -19, -72, 47, 18, -122, -30, -116, -119, 3, -41, -42, 119, -29, -51, 46, -24, 93, 62, -54, 113, 76, 2, -1, -70, 68, -20, 70, -25, -28, 36, 99, 70, -79, -119, 91, 118, 83, -104, -55, -122, 2, 86, -60, 111, 111, 35, -91, -110, 23, -4, 51, -123, 99, -79, -55, 19, -118, -105, -90, 102, 18, 26, -7, -59, -97, -75, -52, -123, -95, -51, -1, 16, 91, 75, 79, -109, -75, 27, -32, -20, 9, 28, 89, 81, -11, 82, 120, -21, 102, 66, -122, -44, -30, 65, -47, -2, -119, 69, 109, 17, -123, 114, 69, 103, 127, 34, -72, 11, 31, 95, 119, 46, -60, -125, 114, 88, -14, 15, -83, 44, -70, 52, 88, -88, 97, 28, -6, -75, -118, 110, -60, 4, 104, 34, 3, 32, 127, -108, 108, -124, -10, 8, 9, 37, -72, -36, -8, 60, -95, -95, 67, -71, 113, 77, -73, -70, 12, 97, -22, -53, -104, 73, 43, 104, -32, 125, 87, 99, -85, 66, 48, 8, -40, -36, 62, 106, 5, 96, -114, 94, 110, -27, 54, -67, -35, -117, -48, -110, -10, 46, -20, 96, 71, 98, -30, 13, 79, -52, 69, -74, -124, -45, -79, -122, -48, 113, -82, -110, -60, 1, -35, -112, -68, -115, 80, -29, 86, 28, -67, 115, 102, 79, 105, -22, 43, -97, -39, -79, 10, 44, 50, 119, 73, 19, 23, -51, 107, -25, 101, -50, -9, 121, -96, -93, -122, 43, 1, -65, 117, -114, 29, -43, -50, -42, 46, 106, 84, 114, -14, 125, -20, -13, -128, 70, 75, -117, -74, 28, 41, 3, -46, -2, -112, -75, 39, -125, 4, 76, 92, 82, 91, 11, -40, -11, -44, -31, 44, 87, -26, 95, -33, 126, -62, -17, -49, -27, -2, 75, -96, -13, -9, 67, -29, -42, 56, 46, 90, 96, -44, -40, 118, 7, 41, -70, 115, -66, 60, 55, 105, -102, -80, 114, -51, -28, 24, -22, 127, 34, -70, 78, 30, 114, -127, 79, 20, 35, 22, -123, -118, 78, -74, 30, 20, -86, 122, 104, 28, 92, -66, 119, 57, 15, 62, -33, 19, -108, 37, -59, 92, -50, 59, -59, -14, 3, 126, 49, -75, 35, -73, 115, -33, -75, -36, 87, 15, -63, -68, 91, 8, -37, 66, -30, -17, 77, -91, 25, -26, 33, -17, -49, -47, 108, -58, -110, 105, 104, -29, 103, -128, 112, 57, 64, 79, -118, 42, 123, -124, 23, -96, -50, -84, 59, -118, 121, 11, 17, -106, 18, -18, -46, 59, 13, 25, -92, -62, -84, 101, 77, 35, -79, 53, 8, 51, -103, 53, 15, -121, -69, 26, -74, -37, 113, -78, -69, 107, 123, -66, -40, -124, 19, 119, 108, 81, 79, 100, 0, 108, -82, 107, 31, 97, 45, 106, 108, -47, -21, -8, 44, -79, 115, -114, -90, 115, 100, 125, -68, -57, -120, 4, -125, 123, -5, -10, 79, -71, 59, -61, 9, -64, -9, 34, 126, 12, 123, 82, 70, -65, -67, -45, 117, -74, 123, -121, 57, 121, 19, 75, 10, 33, 27, 126, 127, -17, -30, 7, 49, -108, -4, -92, 101, -60, 28, 102, -119, 81, -102, 36, -36, 93, -48, 20, 72, -28, 4, 78, 118, -47, -8, -59, 62, -52, 42, 37, -65, -12, 116, -107, 23, -50, -19, 1, -81, 84, 122, -47, -30, -10, 127, -20, 75, -28, -4, 84, 39, 41, -30, -68, -109, -42, 19, -119, -38, 41, -81, -67, 75, -21, -89, -81, 88, 56, -55, 51, -14, -79, 23, 72, -78, -114, 32, -104, -32, 33, 81, -56, 0, -11, 1, 89, -85, 112, 16, -41, 86, 45, 4, -106, -15, -80, -105, -55, 42, 124, -97, -62, -23, 23, -88, 3, -64, -29, 56, 16, 89, 43, 24, -19, -1, -66, 126, 64, 2, 102, 83, 54, 115, -124, 52, 105, 8, -67, 22, -90, -58, -92, 49, -47, 95, -21, 41, -122, 41, 22, 40, -119, -84, 118, 79, 53, -116, -100, 34, 61, -54, -41, -34, 101, 35, -69, 108, -89, -111, 22, -73, 104, 56, 114, -24, 5, 98, -32, 6, 97, 11, 18, -107, 55, 82, 118, 55, 125, -48, 88, 92, -21, -76, -15, 52, 112, 60, 40, 94, -95, -84, -94, 31, 94, 122, -89, -115, -108, -59, 2, 114, -23, 120, 59, -80, 39, 15, -100, -82, -83, 16, 32, -41, -50, -85, 26, 125, 124, -73, -71, 104, -10, 68, -82, -31, -122, 35, 2, -9, 46, 97, 94, -1, 105, -81, -2, -109, -28, -37, 20, 57, -98, -41, 91, 63, 86, 30, -67, 116, -65, -9, -14, -20, -80, -7, -11, 27, 30, 81, -53, 1, -99, 95, 21, 115, 21, -23, 15, 126, -19, -39, -116, -96, -111, 42, -102, -22, -126, -2, -18, -100, 93, 13, 0, 101, -59, 98, -91, -39, -51, 121, -60, -48, -42, 24, -28, 42, -90, 61, -33, -67, -95, -109, -12, 107, -73, 60, -62, -105, 13, -71, 38, 82, 4, 87, 77, 127, -100, -115, 110, 53, 46, 80, -35, -10, -117, -104, -83, 2, 60, 114, -79, 11, -78, 82, 77, -17, 10, 44, 62, 99, -20, 72, 53, -100, -17, -64, -68, -125, -54, -48, 98, 1, 7, -16, -60, 66, 63, -30, 32, 29, -103, -55, 67, -116, 115, 66, -98, 43, -83, 72, -18, 55, -9, -81, -110, 76, -104, -123, 124, -122, -49, -13, -54, -52, -85, -116, -69, -3, 31, -105, 96, -11, -66, -115, -59, -9, 64, 14, 45, -23, 71, -11, 42, -80, -83, -51, -2, 112, 116, -46, 18, 12, 81, 104, 93, -36, -109, 62, 69, -55, 13, 24, -14, 24, 125, 10, -39, -51, 9, -27, -25, 79, 95, -49, -108, -47, 88, 104, 99, 5, 58, -16, 52, -125, -26, -71, 60, -43, 14, -122, -48, 38, -34, -69, -106, 55, 72, 118, 37, -7, -3, -33, -80, -33, 64, -59, 45, 107, 82, -98, 118, -56, 56, 32, 0, 81, -114, -108, -28, -67, -43, -58, 95, -19, -18, 50, -111, 27, 75, -31, -109, -2, 70, -7, 30, -38, 30, -92, 13, -76, 88, 32, -126, 21, -60, 53, -61, 33, 66, -114, -108, -103, -106, -105, 108, -36, 116, -68, 117, -7, -46, 127, -59, -117, -107, 100, -124, 23, -40, 106, 118, 36, -65, -37, -127, 99, 103, -109, -117, 108, 126, -47, -28, -77, -8, -106, 104, -41, 124, -17, 34, 17, 111, -75, -90, 98, -53, 82, -104, 37, 77, 119, 81, 20, 5, -110, -26, -67, -29, 125, -68, -116, 48, 58, 46, -110, 8, 116, -62, -78, -118, 122, 115, -36, -109, -98, -3, 18, -121, -18, 101, 59, -110, -112, 29, -24, 27, -72, 85, 98, -64, 73, 114, 27, -106, 60, 61, -103, 104, 104, -87, -55, -65, -105, -104, 49, -60, -26, 97, 46, -125, -88, -1, -34, 68, 81, 87, -2, -64, -82, -98, -36, -121, -54, -69, 7, -89, -43, -14, 36, -104, 119, 108, -56, 13, 63, 55, -30, -125, 68, -43, 117, -82, -24, 8, 16, 127, -10, 39, 46, -76, -81, -122, 25, 65, 123, -109, -119, 95, -125, 23, 121, -95, -74, 113, 114, 16, -123, 19, -40, 61, 116, 40, -62, -127, -54, 88, 73, 71, -105, -6, -98, 14, 57, 68, -98, -90, 127, -13, 120, 59, 69, 17, 108, 5, -49, -109, 25, -60, 90, -18, -76, 5, 125, -88, -89, -89, -96, -44, -39, -3, -71, -85, -41, 5, -22, -53, 125, -32, 5, 73, 9, -127, -27, 108, 110, 67, -80, -34, -14, -31, 97, 99, 119, -16, -64, 102, 31, -62, -98, 37, -75, -87, 83, -120, 3, -106, 38, -6, 91, 50, 96, 59, 95, -62, 115, -64, -58, 95, -128, -126, -1, 0, -20, 51, 12, 93, 93, 84, 48, 36, -42, -11, -91, 39, -123, 88, -13, -75, -15, 72, 60, 30, 110, 63, -127, -4, -104, -56, -121, 89, 100, 108, -103, 57, -65, 65, 42, -51, -47, 42, -45, 42, -9, -75, 97, -61, 60, -118, -23, 117, -63, 48, 1, -20, -100, -70, 11, -13, -104, 69, 62, -4, 44, -115, 71, 54, -76, 28, -124, 54, 54, 3, 78, 57, -62, -101, -85, -81, -78, -92, 112, 99, 79, 33, 48, -103, -13, -100, -50, 24, 87, -60, -73, 54, -87, 78, -93, -50, 3, -96, 24, -18, 101, -93, -83, -15, -24, -61, 30, 104, -52, 16, -79, 102, -112, -107, 52, 113, -94, 116, 28, 116, -30, 46, 51, -80, -35, 117, -42, 93, -121, 64, -29, 78, -102, 125, 4, 99, -45, 7, -114, -39, 66, -58, 19, 37, -115, -5, 2, 14, -102, -54, -31, 98, -123, -91, 15, 119, 68, -30, -123, 90, 20, -39, -28, -67, 62, -9, 93, -21, -17, -76, 30, 8, 19, -1, -7, -22, 81, 112, -35, -1, 61, -45, -121, 6, 36, 7, -76, 94, -49, -78, 79, 96, 78, 90, 63, -4, 88, 48, -8, 44, 59, -23, 74, 96, -78, -121, -118, -97, -38, 116, 96, 83, 105, -5, 13, 68, 80, 126, 3, -24, 105, -22, -2, 23, 99, -43, -110, 76, -118, -9, 110, 51, 58, 122, 57, 83, -96, 71, 114, 66, 76, 61, 44, 35, 66, 86, -128, -101, 97, 17, -91, -61, -44, 118, -45, -22, 43, -126, -94, -96, 30, 70, -60, -120, -127, -117, -74, 41, 48, -90, -117, 126, -82, -65, -1, -43, 84, 110, -54, -123, 49, -9, 13, -46, -84, 79, -60, -106, -42, -16, -32, 86, 76, -12, -98, 101, 7, -15, -29, -91, 105, -46, -104, 84, -54, 62, 127, -4, -64, -115, -60, 98, -109, 13, -74, 44, -105, 4, 63, 117, -41, 24, 105, 83, -94, -54, -86, -14, 18, -5, 125, 33, -27, 70, 118, -70, -30, 123, -94, -118, -86, 5, 81, -3, 125, -57, -57, -82, 68, -97, -11, 29, 15, 47, 70, 110, 14, 117, 108, 72, -10, -117, -88, -107, -123, -9, 115, -35, -124, -58, -118, -84, 95, -112, -77, 67, 10, -41, 36, 86, -30, -123, -128, 59, 74, -84, 74, -124, -52, -14, 7, -4, 40, -100, 12, -2, -36, -106, 106, -74, 72, -63, -107, -112, 25, -39, -101, 112, 45, 20, -77, 36, -53, 106, -65, 72, -121, -11, -37, -117, 4, -122, -125, 122, -9, -20, -25, 84, 113, -40, 20, -99, -9, -26, -69, -7, 60, -112, 81, 83, 16, 27, 51, 65, -30, -23, -76, -125, -64, 80, 10, 90, -98, 11, -16, -122, -113, -37, 74, -104, 112, 125, 118, -124, -76, -46, 49, 107, -36, 21, -79, -94, -48, -106, -117, -6, 51, 17, 7, 118, -28, -32, -54, -43, -100, -116, 43, 17, -85, 58, 94, -103, 64, -86, 10, -100, 83, 67, -8, -114, 37, 3, 108, -98, 20, 88, -95, 67, 1, 93, -112, -48, -74, 68, -113, 106, 66, -101, 125, -116, -10, 105, 51, 100, 94, 127, 123, 80, -35, 64, 82, -24, -75, 78, 90, 26, 108, 96, -28, -5, -17, 113, 29, 89, 38, -32, -4, 91, 45, 16, 117, -64, 66, -114, 36, -32, -21, -9, -41, 13, 56, -1, -111, 98, -50, 120, -54, 69, -89, 103, 41, -123, -26, -117, 109, 96, 14, 88, 66, -22, -106, -2, -100, 1, -110, 37, 107, 16, 55, -10, -72, 117, -19, 125, -120, 93, -118, -88, -94, 94, 2, -74, 46, -69, -34, -120, 27, -80, 39, 117, -92, -124, -118, 1, -62, 45, -94, -50, -78, -52, -49, -5, -37, 26, 6, -58, -127, -71, 45, 57, 111, 48, -7, 36, 26, -66, -119, 22, 54, -123, 26, -114, 12, 71, -67, 125, 92, -8, 7, 2, -81, 78, 69, 74, -62, -25, 0, 74, -34, 112, -28, -23, -70, -81, 85, 105, -32, 80, -33, 95, 10, 62, 89, 125, 50, 29, 79, 9, 21, 86, 38, -30, -65, -41, -70, 75, 88, -116, 37, -6, 75, 111, -105, 38, 98, -96, 49, 5, -33, -102, 12, -112, 22, -35, -5, -111, -102, -49, -44, 77, 63, -95, 4, -4, -68, -6, 49, -112, -36, -18, -128, -31, 60, 49, 120, -90, 80, -53, 31, 44, 113, 9, 106, 114, -69, 54, -125, 25, -92, 44, -7, 92, -128, -82, -75, 61, 120, 14, 46, -111, -24, -117, -83, 27, 35, -53, 36, -128, -18, -99, -69, -1, 51, 6, 29, 79, 120, 106, 34, -128, -39, -29, -76, -91, 93, 51, -92, -11, 3, -120, -65, 32, 17, 81, 4, 103, 90, 26, 54, -110, 47, 67, 71, 81, -41, -115, -109, -19, 16, -30, -32, -46, -120, 11, 11, 107, -9, -91, -74, 121, 6, 71, 64, -100, 123, -103, 11, -8, -97, -101, 44, -33, -20, 45, 80, 82, -98, 38, -69, -79, -99, 62, 118, 9, -8, -120, -34, -122, -93, 113, -36, 6, 48, -52, 105, 112, 53, -50, -2, -28, 14, 46, 28, -32, -63, 42, 11, -77, -74, 63, -90, 81, -70, 50, 121, 116, -20, -115, 67, -108, 106, -120, -20, -8, 116, 12, 39, 35, -74, 48, 15, -25, 14, -53, 74, -39, -2, -124, -114, 21, 126, -36, -74, 47, 57, 43, 91, -74, -112, -123, 36, -59, -81, -65, -3, -44, -116, -119, 111, -26, 65, 32, 102, 0, -71, -53, 24, 30, -15, 34, 93, 48, -66, -30, -31, -101, -89, 5, 124, -116, -7, 32, -125, 94, -44, -5, 34, -33, -100, 22, -78, 93, 78, 108, -118, -58, -108, 125, -46, -50, -49, -99, -15, -32, 21, 77, 37, 125, 105, -71, -55, -75, 1, -126, -115, -67, 43, -52, -24, 63, -112, 5, -60, 111, -41, -89, 77, 97, 44, -61, 55, 35, -48, -44, -59, -53, 50, 56, -98, 34, -31, 53, 8, -71, 46, 122, -47, -35, 43, 64, 38, -45, -70, -118, 41, -50, 72, -39, -4, -34, 16, -65, -86, 69, -126, -47, 111, 100, -116, -112, 65, -19, 109, -90, -31, -93, -84, -105, 15, -34, 84, -68, -61, -128, 74, 71, -102, 68, 24, 56, 16, -54, -65, 65, 51, -70, 104, -112, 19, 24, 18, -55, 119, 69, 75, 52, 50, 108, 3, 26, 13, 47, -59, -122, 118, 122, -52, 124, -125, 49, 91, 23, 46, 61, 10, -87, -5, -119, 91, 111, -26, 104, -93, 42, -22, -39, 119, 28, 47, -61, -82, 119, 124, -87, -126, 37, 47, -102, -57, -90, 15, -127, -33, 120, -13, -82, 20, -59, -5, -71, -58, -95, 120, 69, 127, -124, -117, 109, -20, 19, -51, 74, 119, -37, -61, 48, -52, -43, 105, 123, 42, -9, -76, 41, -50, 12, -109, 37, -29, -32, 44, 41, -74, -4, 19, -38, -73, 12, 46, 47, 110, 66, -22, 101, 55, -116, -120, 98, -20, 49, -119, 89, 102, 124, -88, -93, 4, -91, -45, 9, -53, -28, -11, -108, -110, -121, -25, -44, 42, -71, -41, 67, 117, 48, -116, 104, -80, 85, -40, 81, 119, -97, 98, 27, -32, -104, 109, 87, 101, 49, -118, -6, 26, -72, -71, 10, 121, 16, -113, 37, 99, 10, -79, -53, -99, -126, 32, -43, 88, 28, 21, 26, 81, 24, -81, -117, 115, 11, -94, 9, -55, -78, -125, 124, 20, 84, 10, -74, -13, 33, 8, -25, 14, 22, 65, 39, -1, -87, 17, 48, -115, 14, -40, 122, -77, -113, 55, 86, -65, -5, -68, 50, 98, -6, -73, 119, 16, 3, 20, 32, -6, -62, 79, 98, -26, 79, -22, 83, -109, 8, -112, 103, -89, 104, -60, -78, -6, 56, -30, -45, 92, -81, -123, -102, -98, 114, 11, 27, 99, -113, -74, -49, -39, -116, 17, 120, 100, -51, 103, 81, 93, 27, -28, 73, 119, -116, -28, -113, 62, 85, -104, 113, -17, 86, -19, -13, 69, 98, 34, -72, 85, 106, -106, -15, -38, -104, 16, -95, 67, -78, -81, -9, 76, -84, -48, 40, 103, 71, -75, -31, -100, 120, 127, 17, -104, 52, -50, -124, -108, -71, -23, 123, -46, -78, -128, -69, 22, -59, 73, -51, 24, 1, -17, 113, -52, 97, -82, -14, -126, -17, 101, -3, -86, 10, -43, 96, 9, -89, 95, 59, 65, -85, -85, -65, -104, 80, -60, 77, -123, -92, 71, -108, 120, -6, -95, -34, 27, 47, -86, 10, 106, -80, -121, 48, -39, 113, -8, -128, 13, 86, 117, 125, 74, -25, -92, 101, -67, -111, -67, -107, 102, 2, 126, 61, 5, 52, -82, 44, 79, -112, 36, -113, -92, 41, -84, 64, 117, -102, 70, -37, 104, 2, 66, 15, 101, -7, 77, 122, 61, 13, 106, -23, -60, 29, 44, 77, -67, 96, -75, 80, 8, 74, 84, 4, 27, -55, 48, -124, 67, 42, 99, 96, 53, -11, -29, -103, -75, 5, 8, 120, -46, 47, -46, -116, 111, -11, 9, -72, -116, -110, 58, -123, 38, 112, -90, -107, -101, -118, -49, -83, -125, -107, -69, -66, -67, 9, 16, -32, 60, 125, -128, -100, 6, -32, -59, 8, 6, 33, 48, 75, -109, -112, 82, 27, 76, -12, 120, 70, 63, 7, -81, -16, 120, 87, -111, -45, -101, -22, 53, -66, -91, 14, 67, -61, 70, -79, 0, -41, -114, 62, 95, 124, 68, 56, 87, 8, 49, 127, 81, -118, -115, 118, -106, -36, 4, 64, 111, 29, 97, 53, -77, -123, 67, -68, -97, -21, -64, 54, 122, 96, 1, 22, -98, 65, 78, 14, 60, 58, 65, 63, 78, -57, 45, 28, -36, 24, -28, 57, -102, 11, -60, -73, -26, 63, -65, 14, 43, -40, 4, 67, -124, 8, 33, 79, 54, -70, 42, -55, 107, -74, -113, 62, 63, 112, -16, 26, 44, 18, 32, -102, 107, 113, -58, 6, 10, -119, 104, 93, -115, 67, 83, -102, -36, -73, 121, -21, 65, 48, -96, -45, -35, 88, 6, 12, -114, 77, -119, 82, 31, -112, -55, 3, -66, -117, 46, 73, 114, -101, -42, -126, 44, -93, -40, -109, 45, 36, 36, 94, -94, -122, -2, -4, 52, -9, -88, -46, 90, 32, 110, -36, -89, -98, -93, -100, -4, 26, 75, 72, -60, -110, 15, -16, -103, 48, -99, -1, 39, 109, -94, -99, 34, -90, -6, -34, 1, 57, -119, -19, -52, 69, -62, 119, 13, -19, -72, -112, 25, -72, 22, -19, 2, 70, 105, -64, 10, 53, -116, 55, 70, 126, -26, -119, 91, -6, 86, 37, -122, 121, 10, 109, -114, 4, -78, 36, -30, 4, 58, 115, -109, -48, -50, 56, 102, 117, 11, -121, -20, -97, -15, -35, 12, -6, -13, -2, -117, 13, -117, -48, -43, 72, 13, -74, -118, 70, -111, -59, 38, -69, -82, -84, 105, 20, -97, 50, -88, -51, -17, -118, -22, -127, 28, 97, -128, -11, 36, -12, 2, -48, 52, -91, 97, 103, 60, -59, 11, -61, 11, 102, 37, -104, 91, -43, -16, 16, 96, 36, -4, -29, 31, -67, 110, -123, 70, -37, 14, -50, 36, -50, 18, -48, -15, -11, -39, 108, -112, 65, -61, 109, 106, 46, -77, 24, 59, -8, -62, 30, -107, 123, 115, -26, -103, 65, 103, -88, 114, 126, -34, -54, 72, 22, -47, -103, 45, -88, 16, -18, -45, 86, -7, 68, 60, 109, 103, -55, 126, 31, 110, 60, 95, -99, -128, 124, -123, 27, 14, -102, 90, -54, 0, 78, -55, 92, -85, -77, 113, -82, 62, -13, 103, -52, -5, 46, 121, 18, -128, -19, 63, 71, 49, -44, 93, -74, -104, -63, -32, 106, -26, 11, -35, 28, -52, -111, -42, -1, -19, 109, 17, 121, 34, -5, 71, -78, 1, -112, -46, -2, -127, 63, -2, -21, 96, 46, -3, 117, -70, 79, 105, 47, 82, -100, -15, 125, -4, 78, 40, -28, -110, -49, 68, -23, 94, 64, 4, 39, -108, -91, -96, -67, -88, -108, 111, 109, -126, 61, -124, -119, 71, 103, -49, 107, -81, -93, 111, 126, 120, 4, 93, 106, -127, -63, -41, -110, 6, 70, -77, 89, -2, -54, 97, 0, 6, 48, 61, 36, 55, 57, 47, 87, -103, -43, 50, 41, 4, 120, 89, 46, -115, 18, 85, -25, 67, -83, 42, -95, -19, -99, 26, 56, 5, 103, -99, -73, 70, 75, -120, 14, 32, -22, 100, -77, 85, 17, -109, -128, 95, 16, -99, 29, -87, 13, -14, -53, 48, 16, 4, 15, 125, -118, 107, 108, 29, -84, -19, -24, 81, 65, -48, -17, -125, -91, 18, -45, -23, 100, -95, 80, -120, 89, 106, 72, 116, 104, -100, 18, 48, 59, 83, 120, 30, 23, 40, -97, 93, -78, -68, -108, 93, -74, 114, -84, -86, -123, -3, 51, 93, 83, -96, 90, -34, 66, -72, -12, 14, 85, -56, -57, 63, -87, 13, 46, -40, 97, 60, -47, 55, -15, 0, -84, -44, 41, -69, -81, 26, 119, 76, -107, 16, 62, -9, 107, 91, 9, -30, 25, 91, 91, 26, 123, 3, -26, -45, 82, 24, 10, 97, -20, 116, -90, 44, -119, 104, 118, -79, 59, 78, -38, -101, -14, -90, -17, -29, -74, 97, -127, 118, 44, 56, 72, 47, 20, 106, -122, -4, 96, -46, 29, 11, -33, -33, 72, 98, -74, 125, 62, -99, -26, 108, 29, -31, 100, -6, 26, -66, -16, -63, 68, -43, -56, -3, 98, -102, -64, -51, -51, 101, -72, 77, 25, -110, -49, -81, -2, -57, 33, -30, -104, 55, 85, 107, -10, -26, 83, 98, 68, 114, 10, 112, 34, -87, -84, -3, 34, 78, -10, 72, -116, 17, -69, 82, -10, 24, 62, -103, 73, -42, -49, -15, 119, 40, -59, -7, -117, -84, -102, -90, 57, -17, 124, 107, -106, -47, -115, -51, 107, -116, -105, -95, 9, -15, -56, 2, -121, 82, 124, -117, 22, 57, 27, -86, 58, -38, 24, -59, -24, -42, 100, -55, -17, -103, -16, 93, -66, -29, -87, -114, 61, -56, -14, -93, 78, 26, 96, -37, 40, 41, 4, 34, 95, -70, 100, -123, 111, -108, -14, 78, -113, 60, -70, -33, -65, 56, -4, -57, 86, -68, -58, 109, 65, -15, 89, 19, -106, 122, 39, 72, -14, 122, 107, 100, -77, -123, 108, -62, 32, 34, -100, 12, 56, -119, -112, -67, -112, 55, 82, -57, 126, 67, -108, -114, 39, 63, -110, -105, 120, -96, 55, 94, -61, -114, -113, 7, 105, 45, 56, -54, 74, 17, -90, -6, 55, 57, -104, -42, 33, -122, 22, 56, 45, -81, 127, 20, 127, -67, -32, 53, 71, -18, 101, -111, 18, 32, -42, -29, 101, -121, 100, -47, -34, -75, -90, 86, 116, 1, -97, 47, -62, -11, -4, 96, 6, 98, -17, 27, -7, 66, -101, -117, -102, -72, -126, 89, 90, -11, -91, 89, 29, 96, -4, -105, -32, -95, 58, -97, 97, -56, -7, 19, -79, -6, 90, 117, 64, 93, 122, -43, -5, 109, 6, 54, 74, -41, 86, 124, -37, 29, 85, 84, -46, -125, -98, 59, -113, -103, -118, -97, 92, 40, 41, -108, -100, 103, -113, 24, -98, -95, 5, -67, 110, 56, -47, 29, 38, -105, 0, 59, -50, -77, -77, 36, 115, -126, -103, -76, 16, -64, 55, 107, 9, -27, 66, -58, -59, 72, 71, -115, 76, 53, -26, 49, -121, -18, 5, 59, -26, -66, -98, -126, -79, -16, 94, -43, -62, -127, -70, -84, -114, -92, -115, 15, 126, -97, -118, 11, 39, 75, -119, -32, 59, -122, -31, 75, 87, -37, -112, -46, 116, 124, -98, -107, 30, 105, 97, -70, -62, 87, -30, -51, -4, 44, 83, 85, -100, -40, 118, 86, -85, 112, -10, -34, -119, 113, -41, -112, 19, -45, -37, -92, 120, 86, -73, -22, -128, -116, 127, 89, 40, 45, 21, 121, -25, 89, 88, 98, -4, -79, 4, 31, 103, -97, -108, 68, 21, -72, -66, 27, -97, -104, -48, 23, -77, -43, 18, -38, 43, -33, 81, -84, 84, -86, -124, 25, 117, -7, -43, -126, -4, 51, 44, 125, 80, -93, 112, 62, 113, -100, 13, 77, -38, 10, -99, 26, -57, -81, -26, -90, -36, -67, -60, 6, 28, -44, 23, 64, 61, -72, 77, 109, -34, 24, -12, -102, 35, 80, -14, -101, 60, 40, 59, 106, 54, 56, -93, -118, -61, 46, -30, 104, -65, 123, -32, 117, -21, 45, 114, -103, -17, -67, 113, -94, 95, 22, -4, -3, -77, -53, 65, 117, 28, 63, 23, 83, -107, -75, 127, 24, 10, -65, -34, -80, -112, 99, 121, 79, 79, -98, -34, -109, 63, -64, -26, -110, -31, -98, 12, -122, -68, -21, 29, -99, 107, 48, -29, -28, 117, -69, -44, 82, 103, 34, 21, -49, 1, -56, -124, 40, 89, 11, 76, -5, -112, 41, -71, 17, 17, 33, 88, 114, -17, 8, -80, 10, 49, -117, 45, -26, -110, 37, 80, 72, -104, -119, 78, 10, 112, 101, -72, -119, 60, -10, -51, 3, -40, -83, -95, -43, 112, -37, -41, 2, -57, 20, 106, -7, -2, 46, 26, 24, -80, -105, -31, 63, 100, -72, 48, -59, -21, 23, 61, -76, 19, 57, 55, -73, 71, -128, 23, -37, -31, -127, 10, -3, 12, -10, -29, -83, -5, 90, 109, -116, -41, -84, -93, 56, -88, -48, -10, -84, -36, -83, -26, -20, 68, -77, -119, -96, -31, 87, 4, -110, 97, -112, 44, 115, 40, 25, -20, -72, 71, -24, 113, -99, 12, 102, -2, -33, 122, -22, 21, 67, -106, -68, 50, -119, 84, -86, 38, -17, -27, 25, -19, -61, 12, -67, -121, 15, 62, -94, 89, 108, 58, -13, 83, 35, 120, 6, -5, -47, 2, -22, -32, -121, -121, 94, 75, -55, 86, -70, 95, 32, -116, 70, -70, -80, 96, 109, -38, 113, -120, 125, 3, -21, -100, 94, 104, 97, -30, 64, 74, -84, -124, -40, -104, -40, -22, -80, 109, -63, -98, 86, 58, 36, 99, 119, -44, 53, 110, -77, 68, -116, -81, 108, -2, 125, 91, 23, -51, -26, 47, -8, -118, 21, 39, -34, 78, -71, -95, 93, 31, -46, -98, 1, 41, 18, 20, -61, -42, -108, -115, -85, 40, -16, -15, -43, -58, 82, 93, -93, 42, -95, 96, 82, 103, 92, -111, 98, -115, -63, 40, -75, 10, -69, 116, 26, -66, -82, 1, -35, -4, 75, 109, 24, -128, -126, 49, 52, 80, -74, -23, -109, 113, -32, -97, -96, 84, -100, -115, 64, 9, -128, 61, -86, 103, -5, -61, -86, -93, 20, -47, 20, -124, -3, 37, 71, -84, -31, -60, -110, -109, -66, 68, 108, 121, 24, -17, -5, -73, 75, -66, 121, -98, 21, -103, 13, -95, -107, 13, 121, -72, 106, -5, 73, -54, 32, 62, 75, -127, -3, 18, 74, 60, 73, 118, 118, 119, 92, 111, -27, 117, 40, -93, -10, 117, 99, 44, 55, -70, -113, 45, -49, -43, 26, 25, -113, 40, -51, 18, 50, 73, -55, 57, -18, -113, -104, -77, -31, -61, 19, 73, -93, 95, 125, 120, -89, -66, -76, -118, -28, -24, 56, -73, 70, -78, 124, 90, 88, -119, -2, 3, 52, 122, 3, -95, 7, -19, 9, -61, -86, -48, 68, -113, 30, 59, -98, -79, -95, 14, 90, 14, 2, 76, 43, 79, 80, -90, -86, 26, 50, 96, 38, 114, -85, -43, -51, -24, -59, 106, 116, -42, 87, 60, 49, 103, 34, 96, -29, -96, 81, 36, -2, 109, -57, 22, 46, 65, 44, -42, -2, 61, -62, 112, -50, -11, 17, -86, 84, 13, -49, -70, -53, -44, 30, -61, -109, 32, 25, 61, -17, 102, -119, -90, -73, 55, 48, 20, -64, 107, 36, 55, -90, 50, -44, -42, 81, 3, -44, -120, 7, 27, 64, -107, -122, -47, 124, 45, -92, -49, 59, -77, 74, 3, 106, -120, -17, 106, 82, -52, 58, -15, -11, -54, 106, 67, 57, -43, 71, -108, 24, -45, 46, -71, -32, 64, 64, 3, -111, 55, 76, -100, 22, -1, -28, -49, -93, -82, 90, -74, -52, 73, 1, 28, -8, 48, -3, -123, -39, -73, 97, -52, -41, 103, 72, -9, -118, -41, 72, -17, -90, 126, -71, 70, 9, 126, -12, 60, -6, 65, -64, -108, -40, -7, 10, 70, 6, -65, 122, 81, 45, -122, -82, -2, 45, 116, -96, -112, -81, -37, 71, 89, 105, 59, 10, -83, 81, -13, -62, -39, 29, 67, -122, 8, 75, 100, 124, -66, 73, 81, 54, 96, -107, -1, -65, 34, -113, -27, -20, -48, -15, -86, -17, 69, -32, -114, 122, 12, -5, 114, 75, 38, -57, 2, -97, 29, 127, 65, 41, 8, 116, -107, -44, 42, -35, -2, -97, 38, -98, 123, 68, 8, -28, -121, -44, -65, 90, -70, -50, -5, -36, 78, 38, 33, 38, -16, -21, -7, 36, -90, 103, -5, -120, -57, -52, -67, -87, 100, 64, -126, 69, 15, 115, -86, -16, 4, 29, -61, -58, 39, -75, -89, 67, 106, -92, 73, 75, -100, -11, 109, -57, 75, 126, 86, 50, -26, 72, 4, -25, 106, -72, 0, -8, -33, 37, 21, -60, 67, -36, -19, 42, 41, 28, -83, 16, -67, -104, -50, 3, 93, 35, 27, 79, -77, -8, -60, 77, 69, -62, -60, -38, -28, 120, -116, -93, -72, -40, 92, -107, 67, 57, 107, -50, 114, 23, -5, 65, -2, -18, 39, 2, 87, -49, -61, -92, 58, 104, -57, -127, 94, -84, -76, -21, 14, -105, 104, 22, -118, -79, 88, 91, 94, 77, 62, -2, -21, -75, -53, 92, 122, 7, 57, 58, -5, 31, 125, -123, 64, -32, -8, -46, -52, -37, 75, 118, -72, -97, 26, 16, 114, 16, -41, -104, 64, 85, -73, -101, -67, 55, -40, 9, 106, 69, -16, 68, -43, -69, 63, -127, 125, -52, -96, -4, 57, 92, 120, 12, -19, -62, -98, 114, 67, -21, 81, 95, -21, -28, 71, 99, 17, -92, 33, -124, -73, -122, -105, -89, -5, -67, 37, -31, 65, 102, -22, -52, -80, 118, -50, -41, -116, -6, -85, 33, 53, 14, 100, 63, 124, 59, 124, -117, -121, -48, 23, 62, -27, 41, 103, -109, 55, 126, -56, -29, 89, -109, -49, -50, 85, -25, -38, 115, -3, -125, 78, -128, -126, 90, -116, -67, 86, -28, 38, -65, 115, -63, -79, -127, 60, 33, 83, -55, -118, 42, -55, -97, -12, -6, 53, 2, -103, -76, -18, -33, 62, 28, -117, -15, -108, -33, -32, -122, -126, 77, -59, 15, 51, 53, -97, -39, 60, -40, 126, -51, -99, 72, -31, 3, -111, 124, 59, -3, 27, 23, 88, 126, -18, -83, 51, -128, -10, -63, -63, 84, 70, 32, -101, 47, -54, -68, 38, 97, -23, 94, -4, -118, 65, -21, -20, 16, 117, 62, 85, -101, -27, 126, 42, -109, -15, 45, 84, 102, 27, -125, 41, 17, -109, -123, -23, 4, 79, 7, 44, 45, 121, 57, -26, -128, 50, -49, 46, 51, 119, 70, 71, 78, -88, -66, 87, 74, -77, -100, -101, -53, -60, -71, -37, 0, -84, -4, -115, 4, -76, -80, 21, -79, -111, -78, 2, -19, -91, 105, -45, -17, 116, -17, 93, -116, 7, -110, -70, 109, -18, -63, -50, 7, 13, -19, 41, -81, 85, 38, -127, -63, -9, 5, 46, -50, -73, -43, 24, -96, 27, 119, -100, 122, -83, -7, 121, -41, -40, -67, -37, 33, 59, -67, -63, 40, 50, -19, -42, 107, -84, 19, 123, 123, 30, 104, 20, -105, 61, 62, 102, 33, -106, 65, 91, 62, -6, 3, -36, -36, 49, -95, 61, -109, -43, -98, -79, -66, 75, -88, 119, 93, 10, 91, 111, -52, -108, 100, 87, 88, -37, -13, 120, -107, 78, -99, -7, 6, -15, -117, 60, -29, 59, 81, -31, -7, -70, 102, 100, -128, -49, 37, -98, -1, -121, -123, -117, -70, -117, 95, -4, 56, 87, -45, -88, 64, -106, 83, 64, 30, -105, -106, -115, 109, 42, 70, 11, 110, -79, -83, 40, -27, 38, -81, -102, 67, -10, -82, -18, -115, 88, -45, 102, 85, 103, -63, -64, 46, 36, -21, -101, 62, 107, -84, 17, -24, 5, -14, 64, 84, -105, -122, 72, 70, -67, 86, 27, 26, 96, 127, -70, 125, 100, 54, -17, 60, 103, 109, 62, 16, -114, -5, 35, 120, -106, 21, 4, -26, -73, -92, -69, 63, -83, -44, -128, 36, 81, 12, -117, -103, 13, 86, 3, -93, -67, -109, -94, 97, -3, -66, 68, 71, 64, 120, 10, -108, 123, 50, -8, -112, 111, 46, 11, -55, -76, -35, -92, 4, -58, 112, 114, -118, -56, -13, 112, -128, 103, 119, -37, -82, -36, -122, 13, 91, 68, -74, 21, 2, 94, 14, 62, -109, -77, -91, 26, 45, 21, -13, 76, 118, 42, -101, 80, 13, 53, 56, -103, -66, -103, 121, 86, -3, -54, -31, 42, -66, -126, -31, -109, 14, 14, -63, 58, -42, -45, 31, -1, 119, 124, 75, 16, -56, 7, 58, 3, 27, 29, 114, -64, 72, -102, -82, -51, -68, 77, -78, -57, 38, -101, 111, -18, 76, 127, 110, -2, 36, 95, 65, -23, 126, 106, -127, -78, 42, -121, -47, 44, 78, -6, -62, -109, 23, -77, 125, -95, 124, 100, -112, 86, 127, 33, -126, 101, 90, -40, 54, 44, -81, -101, 1, -26, 47, -71, -126, 108, 77, 74, 83, 71, 124, -98, 80, -38, -125, -36, -110, 65, -11, -79, -117, 69, -95, -57, -69, 64, 4, -27, -19, -4, 85, 107, 12, -56, 21, -106, 102, -7, -62, 21, -89, -112, 14, 52, 118, 8, -80, -111, -8, -36, -39, -47, -53, -36, -28, -11, 112, -46, 17, 38, 36, -33, 74, 51, -28, 2, 126, 95, -37, 115, -31, -107, -121, 97, 103, 70, -32, -61, 67, 14, 60, 30, -79, 53, -70, 54, -118, 107, -3, 121, -104, -108, 69, -54, 51, -66, 92, -97, -15, -22, -20, -62, 72, -122, -105, 125, 77, -28, 45, -82, 11, -82, 93, -27, -55, -48, -81, -81, 81, 115, 16, -128, -106, 21, 15, 109, 76, -121, -14, 73, 100, -122, 1, 84, 96, -73, -119, 20, -57, 49, 83, 34, 122, -113, 56, -7, 8, -35, -60, 67, -125, 107, -121, 115, 42, 101, 9, 27, -106, -89, -1, 83, -128, 126, -95, -85, 58, 17, 15, -114, 64, 103, -48, -64, -85, -95, -2, -12, -86, 65, 61, -19, 11, -128, -3, -95, -22, 110, 66, 6, -30, 2, -109, -103, 44, 126, 103, -117, -64, 118, -114, -43, 37, -56, 100, -34, -55, -115, -26, -23, -26, -74, -7, 108, 52, 63, -115, -99, 9, 97, 37, -65, -2, -41, 10, 23, -49, -31, 80, -24, -111, 116, -126, 57, -46, 32, -43, -102, -26, 26, -6, 32, 64, -101, 92, 80, -123, 84, -117, -122, 77, 43, -110, -103, -95, -8, -13, 12, -5, -104, -98, -45, -74, -66, -7, 61, 12, -58, -96, -8, 103, 28, -107, -30, -37, 12, 82, 39, -46, -74, -77, -64, 124, 53, 4, -24, -26, 31, 119, -36, -112, 123, 83, -5, -118, -123, -27, 89, -28, -31, -101, 27, -123, 35, 125, 45, -120, 95, -20, -8, -78, -25, 9, 12, 52, 11, -64, 111, 25, 25, -49, -7, 66, 82, 68, -87, -30, 76, 69, -8, 53, 91, 35, 125, -75, 99, -41, -75, -2, 110, -2, 73, 51, -43, 0, -110, -120, -21, -79, 71, 91, -18, -57, -61, -48, 121, -123, -27, -19, -21, -42, 7, -24, -33, -116, 101, 69, 10, -59, 81, 127, -45, -101, -16, -29, -122, 4, 37, -5, 55, -103, -10, -20, 82, -76, 83, 126, -85, 92, -126, -90, 116, 106, -58, -77, -60, 79, 82, 55, 115, -65, -59, 38, -70, 34, -24, -27, 88, -50, 5, 47, 25, -26, 25, 119, 15, 108, 120, -54, -63, 6, -60, 89, -31, 76, -15, -37, 12, 124, 81, 115, 109, 82, -110, 61, -94, 56, 117, -8, -79, 6, -38, -76, -5, -30, -14, -112, -122, -81, -1, -125, -11, -81, -74, -28, 91, -81, -112, 20, 65, -32, 92, 109, 52, 5, -109, 107, -118, 66, -41, 94, 11, -112, 20, 58, -9, -43, 88, -20, 106, -100, 71, -70, -26, -27, 113, -54, -49, -27, 111, 75, 21, 5, -87, 45, 33, -68, -31, -111, -84, 63, -5, -78, 31, 89, 15, -52, -63, 67, 92, -69, -71, -60, 70, -95, -124, -82, 47, 20, -119, 30, -103, -93, 13, -23, -16, -66, 83, -113, -89, 11, -53, 8, -77, -22, 12, 24, 63, 101, -109, -75, 42, -86, 33, -25, -13, 77, -58, 95, 21, -90, -68, -41, 65, -44, 32, 39, 16, -73, -103, -14, -46, 109, -102, 117, -123, -77, 73, 57, -9, 43, -99, -66, -116, 127, -96, -14, 30, 21, 44, -35, -62, 53, -35, -3, -58, 2, -122, -31, -64, -69, 56, -64, 91, 85, -107, -79, 64, 76, -67, -92, -31, 51, 39, 94, -17, 73, 24, 82, 76, 115, -57, 41, 19, 70, 10, 44, 52, -56, -59, -114, 40, -60, 76, -31, 74, 95, -100, -94, 102, 38, 83, 21, -100, -113, 25, 96, -70, -28, 24, 61, -27, 43, 38, 112, -7, -31, -41, -20, -40, -101, -27, 33, 59, 48, 22, -34, -71, -5, -15, -44, -6, 10, 56, -108, 14, 9, -53, -125, 73, 103, 67, 7, 96, -76, 8, -45, 103, 103, -62, 95, 37, 118, 1, -104, 71, -69, -109, 59, 50, 32, -49, 87, -13, -20, -125, -118, 106, 60, 103, 89, 84, 115, -17, 85, -125, -51, 85, -128, 79, 25, -50, 21, -107, -18, -58, 49, 102, -83, 60, 11, -93, 101, -21, -94, 44, 38, 42, 26, 123, -121, -70, 75, -123, -4, 120, 32, -83, -114, -55, 17, -121, 54, -77, -79, 80, 18, -83, -28, -105, 121, -122, 55, 65, -18, 64, 47, -72, 64, -117, 79, 127, 87, -69, -76, 7, -35, -10, -103, -75, -63, -27, 41, -13, -53, -33, -114, 97, 12, -24, -37, -6, 68, -23, -66, 90, 30, -43, -8, -64, -25, 50, 121, -10, -75, -126, -91, 17, -81, 77, -66, -49, 42, -34, 110, -27, 83, -25, 24, 22, -54, -52, -111, 3, -97, -82, -47, 75, 94, 118, 23, 116, -103, -127, -4, -100, 50, 96, -75, -30, -69, -46, 69, 8, 82, 63, -57, -52, -124, -106, -31, -120, 10, 74, 48, 112, -108, 86, 1, 53, -73, 38, -78, 97, 43, 43, 110, 94, -99, -70, -96, -84, 34, 16, 78, 4, -65, 84, 122, 82, -35, 60, -127, 40, 10, 14, -124, 35, -20, -90, 56, 110, -49, -121, 78, -44, 125, 104, -118, 59, 61, 126, -85, 0, -5, -59, 75, 124, -2, 35, -98, -64, -37, 63, 106, 0, -85, 123, -71, -54, 6, -85, 50, -124, -41, 108, -54, -84, -62, -70, 61, -11, 96, 85, 123, -104, -76, 20, 45, -15, -13, -117, -100, -126, 43, -104, -41, -49, -62, 73, 94, 103, 92, 19, 64, -73, 7, 100, 87, 8, -111, 54, -33, -48, -71, 83, -88, 68, -36, 101, 4, 34, 69, -123, 103, -15, 40, -2, 50, -36, 45, 96, 89, -29, 31, 48, 2, -78, -18, -115, 35, 109, 24, 30, -29, -2, 107, -77, -45, 115, 4, -65, -33, -125, 110, 10, -116, 110, 76, -76, 22, 68, 77, -23, -86, -120, 97, -110, -51, 70, -34, 117, 119, -95, 24, 90, 69, 47, -64, -103, -6, 125, -84, -62, 47, -49, 8, 8, -102, -72, -49, -72, 6, 60, 50, 6, 39, -103, -112, -77, -72, -123, 34, -58, -88, 58, -39, 19, -124, 108, 73, 126, -106, 81, -48, 60, 53, -33, -91, 41, 59, -60, -21, 108, 86, -75, 67, -93, 20, -124, 46, -24, -27, -48, 109, 3, 54, 116, 104, 37, 65, -108, -104, 40, -56, 114, -55, -5, -10, -6, 77, -36, -89, 8, -58, -2, 98, -127, 56, -9, -87, 24, 12, 82, -61, -41, -97, 16, 83, -72, 38, 5, 93, 75, 120, 38, 29, 33, 57, 62, -81, -118, -80, -96, -84, 22, -112, 10, 28, -8, 40, 121, -29, 5, -78, 71, 65, 66, -77, 113, -85, -118, -113, -35, -100, 22, -108, 0, 9, 97, 50, 7, 97, 56, -17, 84, 83, 88, 60, 94, 25, 1, -30, -25, -51, -71, 88, 15, -67, 41, 63, 113, -111, 98, 32, -14, -115, 50, 65, 112, 56, -35, 112, 9, -80, -43, 80, -34, 17, 2, 111, -53, 24, -126, -2, 10, -48, 13, 17, -70, -31, 116, 10, -124, 80, 76, -82, 45, -89, 58, 84, -79, 42, -23, 103, 108, 104, -34, 36, 65, -11, 51, 90, 63, 98, -119, -81, -104, -23, 107, 84, -6, -115, -34, -50, -86, 79, -14, 18, 69, -110, -1, 30, 124, -99, -53, 81, 44, 69, 32, -60, -53, 102, -38, -52, -103, 92, 34, 116, -79, 82, 8, -5, 98, 114, -32, 97, -19, -47, 17, 38, -69, -19, -71, -74, -113, 95, -1, 60, 15, -11, -75, -24, -69, 92, 75, -109, -73, -72, 9, 8, 17, -124, -84, -77, 3, -118, -8, -120, -1, -125, -81, -26, -87, -69, 84, 75, 10, -48, -116, 117, -122, 34, -91, -35, 97, 125, -24, 9, -20, -65, -86, 31, -54, 3, 1, 91, 0, -109, 69, -107, 90, 11, -17, -73, 123, -22, -124, 94, 86, 6, -125, -118, -36, -63, -121, 121, -101, -3, -25, -112, -58, 20, -13, -46, 29, -20, -127, 93, -36, 73, -78, 51, -83, -22, -1, 3, 75, -15, 7, -44, -126, -126, 125, 19, -49, 29, 6, -117, 107, 18, 4, -52, -40, 109, -37, -50, 66, -95, 24, -35, 119, 31, -91, 113, 118, -13, 9, -80, 93, -99, 43, 18, -106, 54, -35, -34, -95, -96, -43, -126, -16, 126, -43, -57, 20, 127, -108, -40, 116, -115, 113, -38, -38, -49, 5, -2, -20, 123, 31, -101, -69, -29, 92, -7, 53, -124, -94, 121, 105, -126, 103, -39, 13, -25, 113, 42, -89, 74, 19, 60, -3, -114, 100, -70, 26, -40, 6, 102, 83, 28, -16, -91, 65, -109, 79, 26, -26, 21, -42, 33, 63, -44, 18, 7, -107, 44, -3, 54, -119, 79, 54, -68, 110, -94, -10, -28, 86, 47, -101, 49, 123, 114, 97, -66, 58, -100, -66, -70, -20, 99, 122, 56, 125, 64, 67, 4, -53, -34, 93, -54, -40, 104, 49, 92, -30, -4, 67, 12, 73, -71, 4, 51, -46, -95, -63, 4, -40, 77, 42, 51, 31, 86, -125, -61, 70, 47, 32, 116, 86, 122, -125, -58, 56, 16, 22, -35, 5, -50, -115, 75, 50, -26, 112, 45, -5, -40, 113, -64, 16, -82, -87, 3, 68, 117, -112, 100, 48, 121, -61, -1, -46, 10, 73, 6, 86, -3, -54, 50, -47, 61, 93, 83, -61, 107, 31, 13, -46, -37, -108, -64, -45, 20, 70, -12, -5, -124, 49, 45, -113, 59, -77, -81, -62, 86, 80, -123, 73, 70, 114, -3, 73, -52, 38, -110, 92, -97, -97, 87, 119, -19, 73, -104, -3, 21, 0, -77, 11, 55, -58, -38, 118, -123, 27, 114, 83, 30, -45, -121, -124, -120, -66, -43, -93, -4, -3, 94, 45, -36, 110, 89, 77, -9, -26, 116, -81, 88, 8, -77, -56, -122, 66, 88, -79, -91, 87, -15, -63, 78, -125, -67, 86, 126, -40, 94, -70, 65, 51, -36, 7, 21, -42, 101, 11, -13, 64, -82, 77, -84, 120, 42, 22, 75, 41, 81, -98, 113, -82, -49, -98, 34, -103, 92, -124, -78, 79, -55, -5, -63, 14, 120, -87, 108, -18, 35, -80, 119, -112, 16, -61, 61, -37, -78, -94, 34, -30, 120, 17, 24, -47, -59, 33, 8, -29, 81, 32, 125, -81, -114, 68, -91, -57, 96, -45, -85, 59, 113, 45, 107, 53, -68, 19, 121, 62, 25, 100, -8, 113, -92, -86, 2, -123, -8, -53, -13, -13, -2, 74, -89, 22, -119, -70, 33, 61, 69, 104, 97, -29, -101, 66, 18, 12, -12, -73, 113, 117, -27, 115, -82, 90, -81, 86, 92, 123, -88, -24, 26, -57, -105, -17, -21, 2, 34, 74, 30, -51, -73, -102, -52, 26, 44, -18, 79, 98, -69, 53, -36, 62, -108, -23, 60, 110, 102, -81, -16, 15, 74, 125, 114, -120, 39, 115, -98, -14, 19, -100, 80, -44, 83, 123, 41, -53, 75, -62, -97, 6, -91, -63, 96, 3, 96, -109, -93, 89, -103, 10, 61, -96, -12, -110, -127, -2, -87, 123, 7, -19, 49, -123, 108, 35, -38, -89, 19, -107, 82, 22, 18, -35, -95, -7, 114, -90, -14, -48, -54, -77, -19, 34, 63, -35, 110, 111, -57, 95, 50, 73, -75, -100, -80, -51, -19, -60, -107, 77, -44, 115, 53, 119, 88, 12, 63, 45, -112, 4, -14, 48, 43, -118, 125, -59, 94, -62, -26, 88, 98, 57, -35, -37, 20, 101, -113, -6, 72, 90, -48, 94, 65, -13, 68, 53, 18, -106, 110, -107, -65, -45, 88, 108, 11, 79, -29, -12, 54, 25, -119, 122, 124, 83, 10, 29, -6, 12, -116, 59, -52, 4, 23, -111, 56, -118, 57, -66, 74, 55, -71, -118, 72, -6, -92, 87, 65, 20, 17, 90, -61, -36, -86, -44, -38, -31, -36, -65, 5, 31, -13, 113, -54, -70, 46, -14, 72, 17, -86, 18, 84, 118, 66, -3, 22, 90, -74, -6, 34, 74, -22, 119, 101, -74, 12, -1, 62, 90, -92, 73, -47, 104, 127, 54, -29, -28, 95, 17, 9, -84, -117, -20, 46, 72, -109, -38, -69, -82, 43, 68, 101, -19, -24, 111, 64, 10, -25, 21, 115, 75, 72, 34, 106, 127, -11, -40, -36, 45, -24, -52, -40, 26, -75, 67, 86, 0, -106, 98, 62, -91, 38, -62, -32, 82, 40, -66, 119, -96, -11, 34, 39, -100, -92, 20, 29, -70, 4, 84, -18, -66, -70, -42, -65, -99, -63, 125, 3, -116, 84, -92, 11, 12, -25, -93, -101, -64, 67, -22, -2, 109, -45, -57, 17, 26, -16, 62, -52, -62, -8, -47, -27, 71, -7, -18, 58, 124, -57, -121, 32, 98, -96, 59, 83, 116, 37, -84, -118, -48, 124, 113, 1, -105, -59, -48, -74, -32, -121, -43, 86, 15, -75, 60, 114, -16, 26, 29, -56, -7, 57, -33, -89, 16, -102, -128, -56, 44, -68, -49, -104, 18, 60, 35, 104, -63, -31, -44, -80, 37, 83, 2, 90, 56, 85, 116, -28, -24, 63, -95, -116, -59, -105, -37, -120, -2, 64, 10, 116, 79, -72, 20, 4, 41, 54, 78, 101, 105, -114, -9, -70, 112, 85, -115, -54, -64, 67, 73, 62, 43, 100, 112, 96, -63, -76, 18, -100, 43, -23, -41, -1, -121, -32, 116, 82, 11, 91, 68, 6, -115, 89, 110, -66, -33, -39, 37, 6, -26, 123, 73, -49, 88, 111, -45, -88, 58, -79, 47, 10, -68, -120, 2, -3, 30, 63, -62, 44, 58, 16, 106, -7, 99, 3, -118, -100, 32, 87, 3, 25, -92, -38, -102, 95, 62, 5, 54, 62, -103, 55, -75, 126, 99, -17, -56, -89, 103, -8, -110, -61, 125, 69, 116, 39, -10, -90, 64, -31, 30, 33, 82, -16, 29, -105, -104, 47, 109, 29, -33, 59, 30, -109, 46, -25, -37, -123, 84, -3, 15, 57, -74, -41, -67, 10, 124, 92, -12, -53, 48, -90, -21, 27, 6, 61, -36, 71, 123, 104, 47, -91, -4, -106, 26, -54, -113, 118, 74, 50, -71, 110, -14, -20, -70, 49, -73, 101, 10, 14, 98, 126, 8, -65, -9, -64, 99, -21, 103, 25, 83, 40, 101, 84, 72, -108, -108, -47, -3, 98, -4, -2, -92, 36, -26, 110, -8, -66, 65, -93, 79, 115, 126, 99, 13, 32, -40, -101, -88, -5, 81, 122, -125, 46, -91, -54, 14, -103, 70, 120, 34, -30, -66, -128, 57, -113, 107, 75, 16, -23, 118, 2, 43, -68, 91, 10, 125, 126, 5, 42, -48, 97, 93, -101, -75, 44, -82, -115, 63, -96, 25, 115, 45, 75, 85, -41, 47, 30, -56, -6, -56, -1, -28, -117, 90, 74, -122, -43, -2, 18, 101, 82, -64, 33, 112, 57, 86, 86, -10, 126, 91, -22, 65, 68, -48, -96, 72, 34, 55, -108, -5, 3, -80, 53, 118, 83, 61, -68, -120, 50, -95, -56, -7, 60, -124, 95, 58, -33, 64, -23, 52, -29, 72, -119, -2, -123, -84, 38, 17, 2, 14, 113, -66, 98, 24, -73, -28, -93, 19, -3, -121, 21, 53, -99, -44, 63, 8, -12, -116, 19, -41, 17, -41, -73, -107, 44, -23, 29, 125, 66, 80, 74, -42, -15, 105, 4, -10, 9, 50, -104, -71, -116, 106, 29, 65, 118, -43, 86, 95, -35, -124, -28, -108, -22, 119, 95, -11, -124, 70, 58, -87, 80, -91, -80, 98, 28, -84, 87, 85, 27, -66, 39, 108, -31, 84, 51, 18, -32, -128, -75, 89, -84, 56, 123, 49, 115, 66, -66, 77, 47, -127, 66, -32, 64, 66, -69, 19, 70, 116, 61, -118, 65, 72, -24, -108, 33, -54, 122, 123, 122, -49, 11, -73, -25, 92, -103, -98, 52, 90, -32, -53, -22, -101, 73, 1, 114, 123, -56, -93, -40, -124, -32, -29, -52, 69, 73, 65, 101, 29, 38, 80, 76, 53, -128, 42, -26, -45, -109, -94, -71, 78, 24, -14, -41, 87, 124, -51, 56, -95, -125, -75, -84, -63, 33, 87, -64, -3, -16, 77, 73, 112, 78, 58, 67, -39, 10, -79, 31, 109, 4, -67, -9, 109, 95, 79, 65, 21, 19, 19, -75, -107, -99, 61, -62, -57, 59, 69, 98, 1, -113, -71, -53, -49, -85, -15, -36, 87, 29, -110, 62, -77, -54, -123, 14, -65, 52, 63, 2, -116, 14, 99, -98, -111, 88, 123, 124, 94, 69, -126, 4, -67, -125, 80, -82, -39, 126, 64, -20, 107, -8, 26, 31, -105, 67, -51, -30, 41, -3, 80, -44, -37, -83, 93, 49, -82, -30, 60, -101, 39, -123, 58, 60, -1, -24, 100, 60, 120, 63, 5, 88, 100, -27, -31, -63, -55, -82, 58, 2, 84, 8, 10, 81, 88, -70, -71, -76, -21, 29, -72, -31, -73, 54, -49, -113, 91, 62, -60, -91, -8, -60, 73, -126, 40, -30, -46, -73, 67, -2, 113, -113, -56, -32, 33, -113, -85, -12, -11, 115, 59, -81, 103, -128, 102, 78, 25, 27, -31, 110, 91, 114, -61, -91, -96, -3, 115, -37, 118, -46, 40, 6, 43, -106, 106, 89, 46, -7, 53, 35, -103, -60, -35, 75, 118, 15, -116, 85, 110, -28, 5, 21, -92, 31, -69, 8, -95, -85, 90, -7, 0, 49, -9, -124, 51, 69, 9, 37, -118, -5, 18, -73, -85, 57, 35, 82, 52, 84, 22, -15, -127, -60, 58, 50, 54, 86, -44, 116, 6, -92, -61, -128, -55, -31, 38, -14, 2, -26, 62, 42, 17, 68, -68, 8, -76, -63, -9, 71, -30, 74, 87, 126, 99, 11, -66, -30, -121, -108, -89, 22, -76, 127, 31, 10, 100, 8, -33, -40, 55, 39, 32, 66, -72, 89, -27, -37, 22, -42, -3, -3, 115, 40, 88, -8, 39, 29, 38, -83, -78, -77, -101, 117, 70, -52, 4, -24, 54, -127, 126, -9, 68, 58, 86, -81, -82, 44, -57, -18, 10, -127, 74, 33, 121, -114, -30, -74, 11, -61, 63, 16, -106, -119, 52, -37, -38, 15, 121, -69, -124, -68, -23, 45, -29, -73, 66, 38, 115, 2, -60, 87, -32, -12, -85, -11, 107, 8, 91, -108, 90, 70, -100, 22, 13, -109, 74, 93, -105, 93, -118, 9, 23, -19, -124, 39, 89, -19, -9, 6, -58, -93, -91, -14, -94, 90, -98, -59, 44, 0, 117, 57, -22, -100, 7, 62, 9, 95, 95, -84, 45, 65, 66, 70, -57, -72, -40, -96, -98, -125, -37, -99, 57, 69, -42, -61, -78, -18, -97, 113, -2, 105, -87, -104, -27, 41, -91, -49, -19, 17, 83, -23, 93, 108, -56, 94, 20, 116, 96, 69, -37, 48, 53, 86, 77, 20, -116, 113, -41, 96, -110, -83, -53, -92, -85, -62, -103, -9, -101, 61, -13, 76, -20, -89, -96, -83, 64, 118, 103, 36, 98, -30, -20, -94, -18, -62, 114, -46, 3, 32, 73, 62, -128, -64, 58, -24, 120, 49, -64, -99, -83, -12, -52, -70, -117, -48, -44, 60, 51, -94, 104, 34, -32, 19, -116, -98, -17, -69, 125, -66, -50, 77, -87, 52, -3, 7, 115, 119, 17, -49, 77, -10, 119, 37, -83, 59, -83, -108, 126, -12, 125, -113, -125, -66, 57, 88, 103, -47, 21, -77, -106, -53, -18, -5, -107, 111, 3, -100, 72, 100, -31, -87, -37, -109, -109, 14, 87, -58, -53, 63, 126, 53, 6, -65, -79, -17, -57, -125, -94, -69, 66, -115, -105, 55, -123, -35, -85, -80, -13, -55, 118, -73, 97, -102, 95, -115, -116, -23, 115, -99, 26, 109, -23, -48, 17, -13, 59, -56, 28, -28, 61, 126, -46, -14, -39, -74, 29, 82, -11, 95, 29, 93, 118, 126, 110, -34, -5, 62, 21, -111, 57, -108, 28, 112, 83, 70, -2, 39, -122, 40, -99, 48, 39, -117, -105, -21, -128, -50, -122, 58, 109, 77, 18, -74, -94, -93, -114, 3, 67, -80, -65, 72, 127, -36, 23, -44, -11, 11, -21, 68, -13, 31, -87, 122, -102, 74, 104, -83, 11, 74, 75, -70, -79, 93, 51, -45, 12, 29, 48, 70, 1, -94, -111, -98, 101, 123, -24, 82, 46, -60, -38, -96, 127, -15, -16, -85, -13, 9, 21, -4, 90, 67, 108, 58, -62, 107, 101, 65, 1, 76, -8, -26, -14, -106, 65, -78, -38, -121, 26, -50, 85, 106, -24, 74, 33, -86, 60, 75, 76, 2, 94, 81, -78, 50, 27, -103, -56, -35, -5, 6, 100, 110, -120, -123, -37, -32, -43, 1, 40, 81, 53, 34, -98, 21, -46, -47, 72, 79, -37, -83, -32, -6, 79, 122, 79, 100, -87, 60, 16, -48, -88, -24, -6, 112, -98, 32, -42, -51, 120, 91, -48, -109, -68, 84, 24, -102, 80, 109, -78, -69, 120, 10, 76, -57, 88, -38, -68, 58, -10, -109, -127, 83, 121, -33, 54, -35, 54, -43, 73, 109, 112, -95, 105, -62, -4, 125, -71, 65, 103, 98, 58, 99, -80, -38, 125, -6, 44, -5, -8, 118, -21, 67, -9, 69, -102, 19, 72, 58, 4, -63, 41, -46, 50, -116, -101, 104, -80, -18, 4, -38, 110, -113, 16, -109, -110, 53, 34, 114, -25, -95, -87, 9, 84, 72, 94, 122, -51, 29, 64, -117, -108, -15, 125, -79, 69, -6, 45, 95, -14, -51, 121, 25, 83, 17, 12, 65, 77, 105, 118, -6, -85, 78, -111, 85, -111, 46, -73, -17, 95, 10, 90, -86, -14, -66, -1, 11, 37, -64, 25, 0, 47, 9, -34, -15, -128, 6, 79, 82, 29, -123, -88, 52, -128, 87, -102, 13, -97, -62, 47, 50, -111, -52, 5, 104, 58, 36, 81, 64, -121, 99, -99, -65, -37, 83, -128, 41, 51, -41, -23, -30, 127, -43, -15, 65, -49, 80, 44, 101, -84, 92, -50, 47, -91, 49, -63, -38, -55, 92, 26, -83, -29, -104, 85, 40, -69, -84, 42, 112, -101, 3, -80, 6, 84, 64, -61, -73, 4, 96, -22, 38, 76, 100, 55, -56, 111, -87, -89, -111, 24, 19, 39, 126, -110, -64, -77, 117, 26, 49, -98, -69, 13, 72, -15, -55, -98, -102, 82, -26, 125, -124, -60, -121, 10, -18, 51, 32, 93, -54, 123, -78, 64, -112, -30, -58, 41, -46, -16, -95, -96, -99, 1, -95, 81, 95, -38, -75, -106, 68, -103, -83, -21, -1, -41, 62, 32, -76, -62, 12, 121, -39, -31, 3, 61, -30, 103, 106, 4, -66, 68, -44, -9, 11, 121, -69, 13, 48, 102, 76, 109, -25, -118, -86, -5, -107, -43, 101, 79, -78, -73, -41, 7, -123, -109, -48, -23, 44, 103, 40, 103, 111, 87, 6, 31, -40, -60, -57, -88, 99, 108, 51, -103, 51, 61, -86, 105, -88, 16, 64, 92, 96, -101, -56, -87, 32, 76, 42, -123, -118, -122, 25, -52, -61, -30, -121, -27, 69, 65, -86, 105, -36, -65, -78, 86, -54, -34, 5, 52, -37, 26, -88, 107, -125, -41, -126, -105, -56, 43, 72, -59, 25, 108, 105, 35, -19, 119, 50, -45, -9, -32, -30, -31, 26, -84, -27, 47, 73, 101, 91, -102, -29, 64, 21, 112, 82, 79, -46, -93, -58, 40, -103, -11, 42, -21, -62, 51, 114, -83, -34, 26, 13, -106, -15, -123, -81, 92, 59, 65, -16, 35, -92, -128, -67, -110, -44, -88, -96, 67, -41, 97, 2, -48, -57, -111, -36, -40, -60, -77, 104, -9, 1, 18, -44, 2, -36, -81, -94, 5, -98, -3, 40, 5, 109, 69, 22, -63, -41, 110, 3, -6, -86, -23, 59, -111, -114, -66, 47, 88, -6, 10, -105, -18, 6, 36, 0, 123, 63, 55, 37, -106, 52, 35, 66, -111, -79, 8, 118, 68, -121, -75, 106, 22, 122, 84, -84, 67, 12, 26, 126, -87, 124, -89, 67, -31, -20, -15, -83, -79, -36, -116, 88, 121, 104, 78, -60, -100, 40, -82, -28, -105, 80, -125, -119, 117, -82, -17, -70, 42, 122, 31, 62, 30, 14, -2, -76, 29, -72, 89, 36, -4, -79, 24, 35, -56, -92, -63, -98, -95, -109, 76, 95, -67, -24, 10, 4, 117, 92, -3, -4, -32, -5, -107, 8, 53, -128, -120, -108, 98, -117, 84, -48, -73, 109, 62, 26, 68, -53, -85, 68, -95, 1, 20, -12, -116, 98, -91, 15, 14, 70, 9, -77, -55, -43, 44, -67, 10, -2, 99, -56, 37, 43, 52, -31, -79, -48, 120, -124, -99, -93, -88, -23, 99, -55, 69, 3, 92, -89, 114, 14, -58, -40, 77, -74, -25, -45, -25, -111, -118, -97, -110, 107, -29, -44, 96, -105, -6, 61, -45, 72, -125, -24, 107, -42, -95, 39, -121, -87, 32, 47, -25, -88, 10, 68, -8, -75, 36, -115, -65, -126, 17, 95, 93, -55, -121, 28, -21, -22, -51, 127, 42, -128, 126, -106, -109, 39, -38, 57, 126, -120, 42, -5, -89, -117, 15, 72, -86, -2, 109, -25, -16, -24, 60, 96, 100, -124, 90, 108, 6, -84, -56, 96, 40, 74, 33, -66, -27, -39, 31, -23, 45, 2, -42, 17, 121, 28, -9, 18, -122, 113, -81, -37, 32, 117, -111, 90, -70, -57, -116, -33, 63, -127, -51, 84, -66, 69, -106, -10, -63, 74, 119, 81, -26, 46, 65, 67, -62, 127, -59, 18, -81, -105, -59, -110, -91, -119, 120, 43, -128, -4, 69, -22, -63, 19, -90, 100, 35, -20, 96, 24, 0, -127, -52, 0, 40, 44, -118, -95, -69, -70, 102, 37, 80, 39, 73, 48, 16, 40, 118, 64, -115, 121, 70, 23, 72, 66, 25, 116, -50, -63, 66, -84, -83, -107, 25, -92, 0, -120, 26, 59, 43, 66, -109, 5, 85, -53, 94, -88, -108, -71, -101, -76, -81, -118, -41, -125, -104, -5, -77, -74, 18, -28, -63, -127, -33, -49, -101, 35, -106, 91, 78, 38, 46, 46, 104, 2, 37, 92, 111, 50, 47, 8, 13, 16, 106, -66, -8, 103, 49, 124, 50, -55, -76, 92, -88, 0, 15, -84, 63, -18, 98, -77, 88, 67, -38, 112, 46, 85, 105, 65, -76, 113, -53, 57, 91, 34, 16, 67, -7, 124, -64, -83, 108, -10, 39, -100, -34, 118, 125, -41, -38, 9, 3, 3, 63, -128, 123, 61, 53, 117, 99, -41, 54, -106, 96, 24, -90, -119, 52, 74, -30, 78, 107, 101, 62, -13, 8, 109, 67, 106, 53, -47, -100, 91, 29, 69, 32, -114, 79, -2, -103, 14, 36, -26, -66, 81, 97, -84, -54, -115, 37, -11, 70, -78, -37, 0, -77, 72, 73, -46, -105, -14, 4, 36, 62, 99, 97, 43, -119, 55, -6, -117, 73, 90, -65, -120, -85, 80, -32, -58, 59, 97, -12, 45, 84, -60, -117, 17, -100, -107, 64, -36, 42, 45, 122, 14, -51, 126, 11, -40, 4, -49, -45, 33, 90, 121, 98, -43, -45, -122, -108, -26, 9, 84, -75, 8, 127, -41, 109, -87, -12, -58, 30, 113, 91, -64, -76, -31, 95, -23, 102, -83, 76, 43, 91, 26, 71, 116, -117, -76, -115, -121, -119, 10, -127, 15, -38, -8, 82, 33, 41, -72, 13, 101, -55, 114, -60, 47, 73, -89, -59, 2, -51, -52, -8, -99, 0, -123, 55, 22, 36, -110, -107, 107, -117, -94, -90, 109, -57, 91, -122, 117, -32, -29, -4, 110, -6, 70, 90, -18, 29, -93, 70, -51, -108, 71, 10, -111, 110, -74, 48, 92, 77, -91, -92, -49, -77, -127, -72, 12, -99, 13, -30, -39, -6, 116, 100, 46, -123, 38, 65, 54, -93, 89, 102, -67, 79, -86, 84, 41, 8, 111, -16, 78, 18, 78, 51, -28, -106, 111, -74, -13, 107, -33, 45, 68, 63, -55, -55, -127, 10, -86, 101, -28, -82, -97, 66, 112, -121, 106, 50, 5, -33, 105, -58, -121, 75, -95, -26, 102, 51, -96, -88, 79, -121, 95, 8, -87, 73, 25, 109, 31, 79, 8, 110, 22, 43, -102, -3, 61, 44, -45, -55, -20, 113, 63, -91, 87, -53, 44, -117, -19, 3, -81, 22, -52, 108, -69, 63, -85, -20, 44, -31, -96, -95, 21, 94, -64, -10, -30, 11, -92, 126, -55, 24, -106, 102, -83, -51, -11, 117, 15, -122, 86, 71, -91, 92, 100, -128, -42, 117, -17, 125, 14, 82, -46, -80, -88, -41, 123, 1, 93, -38, -86, 41, 106, 112, 13, -19, 24, -64, 46, 102, -25, 25, -33, -48, -95, 91, 9, 101, 19, -78, -51, 46, 12, -83, -35, 125, -105, -50, 77, 41, -110, 3, 13, -24, 126, -76, -109, 62, -62, 66, 5, 53, 74, 68, -48, 100, -101, -95, 11, -90, 13, 29, 22, 84, 56, 117, -105, 64, -85, 87, -41, 16, -96, -50, -77, -101, -127, 106, 119, -57, -7, 65, -66, -112, -128, -26, -29, -4, -33, 64, 117, 89, 127, -107, 46, 116, -72, 30, 52, 126, 58, 109, 116, -107, -15, -99, 105, -19, -48, 54, -74, 3, -6, 88, -65, -89, -112, -118, -23, 51 );
    signal scenario_output : scenario_type :=( 127, 127, 127, -128, -128, 127, -17, -128, -128, 127, 127, -128, 127, 42, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 113, -128, 127, 22, -128, 54, -128, -128, 127, -128, 71, -101, 127, -123, 127, 127, -57, 127, 127, 127, 107, -128, -128, 127, 127, -128, 127, -87, -128, 127, 127, 127, 127, 127, -36, -128, -128, -128, 127, -101, -128, 127, -64, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 66, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 114, 92, 127, -128, -128, 127, -100, 127, 127, -21, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -42, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -26, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 47, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -113, -128, 127, -91, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -64, -128, -128, -59, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -38, -48, 127, -128, 90, 127, -128, 127, 127, -128, -128, 127, -128, 127, 106, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, 127, 27, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 112, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -28, 127, 127, 127, 127, 127, 127, 127, -128, -128, -55, 127, 127, 127, 127, 127, 127, 127, -111, 127, 127, -128, 127, 127, -128, -128, 17, -128, 127, 79, -128, 74, -128, -128, -33, -128, 127, 127, 127, -128, 127, 127, 127, -55, 127, -128, 127, 127, 127, 121, 80, 127, -128, -128, 127, 127, 127, 127, 127, 127, 122, 127, 127, 127, 127, -128, 127, 127, -128, 127, 33, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 114, -128, -128, 27, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -95, 127, 127, 127, -128, -128, -128, 63, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 101, 127, -128, -128, -128, -128, -17, 127, 127, 127, 127, 113, -128, -128, -128, -128, -128, -128, -10, 127, -128, 127, 127, 127, 127, 127, -32, 127, 127, -128, -18, -53, -128, -128, -28, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 91, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -17, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 102, 127, 127, 127, 127, -128, -128, 127, 127, -128, -107, 127, -128, 12, 127, -128, -128, -128, -128, -128, -128, -101, -128, 127, -128, 127, -128, -3, 127, -128, -128, 127, 127, 127, 127, -122, 119, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -109, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 87, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 116, -128, 127, -47, -128, 127, -128, -128, -128, -128, -128, -128, -128, 13, 127, 127, -128, 70, 127, 127, 127, -128, 127, -108, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 10, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, -36, 127, 127, -128, 127, -128, -128, -6, -128, -16, 127, -128, 5, 127, 127, -128, 127, -128, -128, 127, -95, 127, 127, -128, -128, 127, -128, -6, 24, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, 87, 127, -121, -128, 127, -23, -128, 127, -128, -128, 70, -128, -128, -128, -128, 127, 91, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 86, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 75, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 81, 127, 127, 127, -128, 127, -5, -128, 11, 127, -16, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 23, -54, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -58, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, 60, -128, 97, 127, 26, 127, -128, -128, 73, -128, -88, 127, -128, -128, -128, 127, -128, -128, 101, 127, 127, -128, -128, 92, 127, -1, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 29, 28, 127, 127, 127, -66, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -10, -128, 127, -128, -128, -128, 108, 127, -128, -128, -128, 127, -128, -128, -44, -128, -128, 127, 127, 121, 127, 127, -128, -128, 127, 127, -128, -128, 3, 127, 122, -128, 127, 127, 127, -106, -128, -128, -128, 127, 102, -128, 127, 127, -128, -27, -108, -128, -128, -128, 98, 127, 127, 127, 127, 127, 127, 127, 127, -79, -128, -128, -128, 127, 127, 127, 127, -128, 31, 127, -128, -128, 127, -23, 127, -128, -128, -103, 127, 127, -74, -26, 127, -128, 127, 127, -128, -128, -128, 36, 127, -128, -128, 127, 127, 127, 127, -117, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 49, -128, 11, 127, -128, -8, -128, -128, -128, -128, 6, 127, 127, 127, -128, -128, -128, 127, 54, 127, 127, 127, 127, -128, -23, -128, -128, -52, -128, -128, 68, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -107, 127, -128, -128, 127, -128, 127, -21, -128, 127, -128, -128, 127, -2, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 10, -128, 127, -128, -128, -81, -128, -128, 10, -128, -128, -44, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 48, -128, 127, 127, -128, 127, -42, -128, 127, -128, -128, 127, 127, 127, -33, -128, -128, 127, -128, 96, 127, 123, 127, 127, -128, -128, -111, -128, -128, -128, -128, -128, -128, 127, 127, -128, -65, -128, -128, 127, -128, 127, 127, -68, -128, -128, -119, -128, -128, 127, -109, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -26, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -76, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -102, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -114, 127, -80, -128, 127, -6, -128, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 29, -128, -128, 127, 127, -111, 127, 127, 127, -128, 127, -128, -128, -29, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 106, 127, 127, 127, 2, -128, 109, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -65, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -5, 1, -5, 127, -128, -128, 127, 127, 127, 127, 10, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -97, 127, 127, 127, -128, -128, -128, 127, 127, -128, 81, 127, 127, 127, 127, 127, 127, 127, -32, 127, -128, 127, 127, -128, 111, 127, 127, 127, -121, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 118, -128, -128, 127, 127, 127, 127, -91, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -53, 127, 127, -128, -128, 127, -96, -128, 127, 111, -81, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -5, -128, 127, 127, -128, 127, 123, -128, 70, -128, 127, -128, -121, -128, -128, 127, 127, 127, 127, 16, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -102, 127, 127, 127, 127, -128, -128, 127, -128, 127, -111, -119, 127, -128, 127, -90, -128, 127, 127, 103, -128, -128, -124, 127, -128, 127, 96, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -124, -31, 127, 127, 127, 6, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 6, -128, -128, 127, 78, -128, 127, 127, -95, 127, 127, 127, 127, 127, 127, 127, -128, -128, 119, 127, -38, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -95, 127, -128, -128, 127, -109, 127, 127, -128, -128, 5, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 0, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -65, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 24, -128, -128, 127, 127, -128, -128, 127, 127, 121, 127, 127, 127, 127, -128, -128, 64, 127, -128, -128, 127, 127, -128, 127, 127, 127, 7, 31, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, 127, -128, -21, 127, -113, 80, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 87, -128, 127, 127, 127, 127, 118, -128, 6, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -17, 127, 127, 127, -128, 88, 127, 127, 127, 127, 127, 127, 127, 38, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 114, 127, 127, 127, -128, -128, -103, 127, 127, 127, -128, -16, 127, 127, -128, -128, -128, -128, -128, -128, 127, -112, 127, 127, 127, 127, -128, -47, 127, 127, 127, 127, 127, 127, 127, 127, -128, -52, -128, 127, 106, 127, -128, -128, 127, -128, 124, 127, -79, 127, 127, -37, -128, 127, -128, 127, 127, 29, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 18, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -75, -128, -128, -128, -128, -128, -128, -128, -128, 127, -52, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -102, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -1, -128, -128, 0, -128, 127, 127, -128, 127, -128, -93, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 71, -128, -128, 127, 127, -128, -128, 45, -128, -128, 127, -90, -128, 127, 127, 127, -44, -128, -128, -128, -128, -128, -128, -128, 127, 38, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 113, 127, 127, -47, -128, -128, 127, 127, -96, -128, -128, 127, 127, 127, -118, -128, -128, -128, 127, 127, -128, 127, 121, 26, 127, -128, 127, -128, -128, 127, 127, 117, 127, -128, 127, -128, 34, 13, -128, -73, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 5, -128, -128, -128, -128, -128, -128, -128, 86, 127, 74, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 74, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 54, 127, 127, -128, 127, 127, 127, 127, 127, -42, -128, -128, -128, -128, 127, -128, -128, -128, -22, -128, 127, -128, -128, -128, 71, 127, 127, -128, -22, 78, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 10, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 121, -128, -97, -128, -128, 127, 108, 127, 127, -128, -128, -128, 127, -128, -128, 127, 114, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 22, 127, -16, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -16, 127, -128, 127, 127, 127, -71, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -108, -128, -128, -128, 127, 0, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 114, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 92, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -74, -128, 127, -128, 127, 127, -128, -6, 78, 127, 103, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 100, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 37, 127, -86, 127, 127, 73, 127, 34, -54, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 103, -128, 127, -96, -128, 127, 127, 127, 127, 127, 127, -113, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -108, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -63, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, 90, 22, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 59, -128, -128, -38, -128, -128, 127, -128, 127, -18, -128, 127, 127, 127, -128, -128, 127, 127, -13, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 68, 127, -98, -128, 127, -128, 98, -128, 95, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -26, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -43, -128, 118, 127, 127, 63, 127, -128, -128, 127, -128, 127, -68, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 33, 38, -128, 66, -128, -128, -128, 127, -128, 123, -128, -128, -128, -128, -128, -128, 127, 16, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 98, -128, -128, -128, -128, -123, -128, -128, -128, 127, -128, -128, -128, -128, 123, 127, 127, 127, 127, 127, 127, -128, -6, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -92, 127, -65, -128, 127, -128, -128, -128, -128, -128, -128, 127, -18, -128, 127, -128, 8, 127, 127, 127, 127, 1, -128, -24, -128, -128, -112, 127, 13, 127, 127, 127, 87, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -48, 127, -18, -128, 127, 8, 118, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -8, 127, 127, 116, -128, 127, -128, 127, -111, -128, -128, -128, -128, -127, 127, -128, 127, 127, 59, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -3, -128, -128, 2, -128, 127, 127, -128, 127, 127, 3, 127, 127, -128, 68, 127, 127, 127, -128, 109, -128, -73, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 10, 54, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -63, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -114, 69, -128, 127, 127, -128, -39, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 57, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 106, 127, 127, 127, 127, 127, 127, 127, 127, -128, 1, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 27, -128, -128, 127, 48, -128, -128, -128, -58, 127, 127, 127, -128, 127, 127, -114, 127, -128, 127, -128, -116, 127, -128, -128, -13, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 22, -128, 127, -128, 127, 127, 127, 127, 127, -78, -128, 16, 127, -128, -128, 127, -127, -128, -128, 127, -128, 127, 127, -128, -47, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -55, -128, 127, 127, -124, -128, -128, -128, -8, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 43, -128, 127, -80, -128, -124, -10, -128, 81, 127, -128, -128, -128, -128, -128, 127, 2, 127, 127, 127, 127, 127, 127, 71, 26, 80, -128, -31, 127, -128, 0, 127, 91, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 122, -128, -128, 86, -7, -128, -128, -128, -119, -128, -128, 127, 127, 119, 127, 127, -78, -128, -128, -128, -128, -128, 13, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -106, -128, 127, 127, -70, -128, -128, -128, -128, -11, 127, 127, 127, 127, 127, -36, -128, -128, 44, -128, -128, -12, 127, 127, -128, -85, -112, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 90, -128, -128, -128, -10, -128, -117, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 7, -8, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -47, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 98, 127, -128, -128, 127, 127, 15, -128, -128, -128, 127, -49, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 80, -128, -128, 127, -128, -128, -128, 101, 59, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 96, 127, -44, -128, 36, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -79, 127, 127, 127, -128, 59, -128, -128, 127, 127, 127, 127, -128, -128, -79, 127, 127, 127, -128, 127, 127, -128, 127, -44, -128, -128, -128, 127, 127, 127, 80, -128, -128, 127, 127, -128, -21, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 93, 127, -128, 127, -122, 127, 127, 127, 127, -128, -100, 102, -128, 127, -128, -128, -128, 127, 127, 127, -58, -128, -128, 127, 127, 55, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -122, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, -97, -128, 127, -128, 7, 127, -128, -128, 60, 127, -128, 127, 127, -128, -128, -128, -128, -8, 127, -128, -103, -128, -128, 127, -128, 127, 127, -128, 127, 127, -8, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -26, -52, 127, -128, -128, -88, 127, 127, 127, 127, 116, 127, 127, 127, 90, 127, -128, -128, -128, 113, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 5, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 109, 127, -128, -128, -128, -128, 127, -128, -128, 127, -18, 8, -128, -128, -128, 127, 127, 42, 127, 127, 127, 127, 127, 127, -128, -128, 127, -118, -128, 127, -128, -128, -128, 127, -91, 63, -66, -128, -128, -128, 76, 127, 127, 127, 90, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -64, 127, 127, 127, -128, -128, -128, -3, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 42, 127, -128, -128, -128, -128, -128, -128, 2, 127, 127, 127, -128, -128, 127, 127, 127, -114, -128, -128, -128, -128, 127, 127, 127, -128, -128, 111, -128, 118, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 81, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -28, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 28, 127, 127, 68, -128, 54, -128, -128, -128, 127, 127, -128, 127, 127, -87, 127, -114, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, -79, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -79, -128, 127, 53, -80, 127, -128, -128, 60, -128, 127, 127, 127, 127, 127, 127, 127, -128, 74, 32, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -47, 127, -128, -128, -36, 127, -128, -128, -15, -128, -128, 127, 75, -128, 98, -128, 34, 127, -128, -128, 101, -128, 127, 127, 127, 127, 57, -128, 127, 73, -128, -128, 127, 127, -128, -128, 127, 29, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -8, 127, 127, -128, -128, -128, -128, 127, -13, 127, -22, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 29, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 90, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -45, -128, -128, -128, 127, 127, -128, 127, 127, 97, 127, 127, 76, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 3, -128, 127, -128, 127, 127, -128, 11, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -32, 127, -128, -128, -128, 127, -116, 127, 127, 127, -128, -128, 12, -128, -128, -128, -128, 127, 127, 81, 127, -15, -128, -42, -128, 127, 127, 73, 68, 45, 127, -128, -128, -128, -128, 90, -91, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 65, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -75, 127, 127, -128, 127, 127, -128, 127, 12, -128, 127, 127, -128, -128, -128, -24, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -48, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 60, 127, 127, 127, 127, -128, -128, -112, 127, -69, -32, 127, -128, 127, 127, -128, 127, 127, -128, -128, -101, 127, 127, -128, 127, 127, -128, -68, -128, -128, 127, -128, 12, 127, 127, 127, 28, 127, 127, 127, 127, 127, 127, -128, 127, -87, -128, 127, -128, -43, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 37, -128, 127, 127, 2, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 71, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 58, -128, -128, 59, 127, 127, 127, 127, 111, 13, -128, 3, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -78, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -22, 127, -128, -128, -128, -128, -50, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -88, 127, 127, 127, 7, -128, 55, 127, 127, 127, 127, 127, 127, -128, -21, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -114, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -96, 127, 127, 127, 127, 127, 127, 127, -23, 127, 127, -128, 127, 127, -128, -128, -128, -128, 70, 127, 127, 21, 127, -128, -128, 127, 127, 127, 127, 127, 127, -108, -128, -128, -128, -128, -76, 127, 127, 127, 127, 127, 127, 0, 127, -128, -128, 127, -128, -128, -128, -128, 44, 127, 47, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 59, -128, -128, 101, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -49, -128, 127, -128, 127, -128, 58, 127, -128, -128, -128, 127, 127, -80, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -43, 127, 65, -128, 127, -124, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 87, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -58, -128, -128, -128, -128, -128, -128, -128, -128, -50, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, 17, -128, -128, 127, 6, 127, 127, -128, -128, 127, -128, -52, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -12, -128, -128, -128, -128, 127, 5, 6, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 108, -128, -128, -128, -128, 127, 127, 23, 127, 127, 127, -128, -128, -10, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 121, 127, -128, 127, -128, -128, 127, -106, -128, 127, -39, -128, -38, 127, 127, 127, 127, -128, 127, 127, 127, -33, -70, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 36, -128, -128, 127, 47, -127, 127, 96, -128, -128, 127, 127, 127, 127, -128, 57, -128, -128, -128, 127, 1, -128, 127, 127, -10, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 112, 127, 127, -128, -128, -11, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -85, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, 15, -128, -128, -128, -128, 127, -93, -128, 85, -128, -128, -128, 127, 127, 127, 127, -69, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 75, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 48, -128, -128, 7, -45, -128, 38, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 59, 127, -128, 127, 127, -128, -128, 127, 42, 127, 127, -128, 127, 127, 127, 39, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -23, 127, -128, -128, 116, -128, 127, 127, -128, -34, 127, 127, 0, -128, -73, -128, 127, 127, -128, 127, 127, 127, 3, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -81, -128, -128, -128, 15, -128, 127, 127, -128, -128, 127, -128, -128, 124, -128, 127, 127, 49, -128, -128, -33, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -54, -58, 93, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 55, -128, -128, -128, -124, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -107, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 37, 127, 127, 127, -92, -128, 37, 12, 127, 113, -128, 127, -45, -128, -128, -128, 127, -128, 127, 127, -128, -87, 127, 127, 127, 80, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -43, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -75, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -107, -128, -128, 127, 127, 127, 127, 127, -128, 32, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -32, -128, 66, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 92, 127, -128, 85, 58, 127, 127, 127, 127, -128, 113, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -76, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 122, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 114, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -18, -128, -128, -128, 127, 127, -128, 119, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 118, -128, -128, 127, -128, -107, 127, 127, 127, 103, -128, 121, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 60, -128, -66, 127, 127, 127, -128, 127, 127, 13, 127, -128, -128, 127, 123, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -15, -128, -128, 127, 127, -128, -59, 127, 127, 127, -128, -128, -128, -42, -128, 127, -128, 127, 127, 127, 127, 127, -128, 21, 127, 127, 127, 127, 127, -128, -128, 113, -128, 127, 127, 127, 127, 127, 127, 127, -107, -93, -128, -128, -128, -128, -128, 127, 113, 49, 127, -128, -128, -102, 127, -12, 127, -128, 127, 127, 127, -55, 98, -28, -128, 127, -128, 73, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -102, 127, 127, 127, 16, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -34, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -74, 13, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -37, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 23, -128, 22, -128, -128, -128, 127, 127, 127, 127, 127, -128, 69, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 86, -128, -128, -128, 127, 17, 127, 127, -128, -128, -57, 127, 127, -22, 127, -128, -128, 127, 50, -128, 127, -128, -128, 55, -85, 127, 127, 127, 127, 127, 127, 127, -97, 127, 127, -128, 90, 127, -128, 116, 127, 127, 127, 127, 127, -128, -49, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -103, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, -93, -128, -128, 42, -128, -128, -128, -128, 127, -128, -128, 36, 127, -128, 127, 127, -127, 6, -128, 127, -92, 127, 39, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 28, -128, 127, 127, 127, -52, 63, 127, 127, 127, 86, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 2, 127, 127, -128, -128, -128, -128, 127, 29, 127, 117, -128, -128, 127, -128, -128, 127, -128, -128, 127, 116, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, -95, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 38, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 54, -128, 127, -128, -128, 127, -128, 127, 127, -128, -108, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -6, 127, 127, 127, 39, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -18, -128, -3, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -60, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 70, 86, 127, -128, 21, 127, 127, 127, 127, -128, -79, 127, 127, -128, -128, 127, -128, -128, -128, -21, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -123, -128, -128, -128, -128, 127, -128, -128, 118, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 0, -128, -128, 127, -78, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 108, 127, 127, -128, -128, 80, -128, -128, -128, 33, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -111, -128, 22, -128, 127, -128, -7, 127, -128, 28, 127, 127, 127, -128, 127, 16, -55, 127, 127, 3, 127, 127, 127, 16, -39, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 112, 127, 127, 127, -128, -128, -128, -128, -128, -128, -127, 127, 127, 127, -128, -128, 127, 127, -7, -128, -128, 127, 127, 127, 59, -128, -128, -128, -128, 127, 112, -128, 123, 127, -128, -128, 127, 127, -128, -36, -128, -128, -128, 127, -128, -128, 127, 127, -128, -80, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -112, 127, 127, -128, 127, -128, -128, -23, 127, -128, -59, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -37, 127, 127, 127, -59, -128, -69, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 53, 127, 127, -128, -73, 127, 22, 127, -128, 127, 127, -91, 127, 127, 127, 66, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 55, 127, 109, 127, 127, 127, 127, 127, 127, 127, 127, -128, -53, -128, -128, 127, -128, -128, 127, 127, 13, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 47, -128, 127, -128, 127, -128, 127, 127, -128, -109, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 54, -128, 127, 127, -128, 127, 127, 127, 49, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 31, 127, -128, -128, 127, -128, -128, 127, 29, 127, 86, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -103, 97, -128, 127, 127, 127, 127, 127, 127, -57, 127, -128, -128, -38, 127, 127, 127, 127, -128, -128, 127, 127, 106, -128, 127, 127, -128, 127, -128, -76, 52, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -24, -128, -128, -39, 127, 127, 127, 127, 127, -96, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -38, -50, -128, -128, 127, 127, -128, -128, 127, -128, -112, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 6, 127, 127, -128, -128, 127, -15, -128, -128, -128, -128, -128, -128, -128, 118, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -121, -128, 127, 127, 127, 127, -49, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 65, -15, 127, 127, 127, 127, -128, 127, -128, 127, -11, -128, 127, 127, 127, 127, 127, -128, 127, 127, 95, -128, 127, 127, 127, 73, 127, 127, -128, 55, -128, -128, -122, 127, 127, 127, 127, 127, 127, 114, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 38, 127, 127, -97, -128, 127, 127, -128, 127, -128, -128, -128, 32, -128, 55, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -118, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 6, 127, -128, 80, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 24, -128, 127, 127, 127, 127, 127, 66, -113, -47, -128, -128, 127, 127, 127, 127, -28, 127, 127, -128, -128, -128, -128, -80, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -52, -128, 127, 60, 127, 127, 127, 127, 127, -92, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -102, -128, -65, -128, -128, -54, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -69, 6, -128, -50, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 73, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -44, -128, 31, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -109, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, 26, 127, -128, -128, -128, -128, 127, -127, -128, 127, 127, -86, -128, -128, -87, 127, -128, 127, 127, -128, 79, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -114, 127, -128, 106, 127, 127, 127, -98, -128, -128, -128, 127, 127, 127, -128, -128, -128, -17, 127, -128, -128, 65, -128, 127, -128, -128, -74, 127, -121, -128, -128, 127, 23, 127, -60, -128, -128, -128, -128, 76, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, -70, -128, 127, 127, 127, -128, -128, 127, -108, 127, 127, -127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -87, 127, 127, 127, 127, 43, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 18, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 43, -128, -42, -128, -128, 127, 2, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, 0, 127, -128, -49, 127, -128, -128, -128, -128, -24, -128, 127, 127, 127, 127, -97, -43, 127, -128, -128, -128, -128, 124, 127, -128, -128, 127, 127, -128, 127, 127, -128, 101, -128, -128, 127, 92, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -64, -128, 127, -128, -128, 127, 127, 127, 1, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -60, 23, -128, -128, 59, -128, 127, 127, 127, 112, -128, -128, -128, -128, 127, 127, 127, 127, 54, -128, 96, 127, -65, -128, 127, 127, -128, -128, -128, -128, -55, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -60, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 53, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 13, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -116, -128, 47, -43, -128, -128, -128, -128, -128, -128, -128, 127, 127, 76, 127, 127, 127, 127, -88, 81, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 60, -128, -128, 127, -128, -42, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -92, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, 117, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -28, -128, -74, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 108, -128, -106, 102, -128, -128, 127, 127, 127, -128, 50, 45, 127, -128, 127, -128, -128, -128, 127, -65, -128, -18, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 59, -29, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, 12, 127, -128, 127, 127, 28, 127, 127, 127, 127, -128, -128, 65, -128, -128, -128, 11, -128, -128, -128, -128, 127, -128, -128, -128, -128, -95, -128, 98, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, 43, -128, -128, 34, 127, 127, -128, -128, -128, -128, -128, 106, -128, 127, -128, -128, 103, -128, -128, 18, -74, -128, -128, -128, -128, -128, -128, 127, 91, 127, 127, -128, 27, 57, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, -22, 34, -128, -128, 44, -128, -128, -128, -128, 127, -128, 38, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 7, 127, -27, -128, 127, 100, -121, 127, 127, -48, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 32, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 36, -1, 5, 71, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 42, -128, -16, 127, -128, -128, 127, -106, -128, 127, 127, -128, 127, -128, -75, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 88, -128, 127, -81, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -116, 127, 127, -128, 21, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -64, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -23, -5, 127, -128, -128, -128, -128, -128, -128, 127, 127, 96, 127, -128, 87, -128, -128, -128, -128, 127, 127, 127, -128, -48, 69, -128, -86, 127, -128, -128, 127, -128, -128, 69, 127, 127, 127, -128, -128, -128, 127, -128, -128, -2, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 24, -128, -128, -128, -87, 127, -128, 127, 123, 127, 127, -128, -128, -128, -128, -128, 88, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -45, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -103, 0, -128, -2, 127, 127, -128, -128, 127, -128, -128, 127, 0, 127, 127, -128, 28, 127, 38, 127, -128, -128, 6, -128, -128, 127, 127, -128, 57, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -29, 74, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -32, -119, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 85, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 42, 127, 127, 127, 127, -32, 103, 127, 112, -128, -128, -128, -128, 127, 127, 127, -128, -123, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -50, 127, 127, 127, -128, 127, -128, -128, 127, -43, -128, -79, -128, -128, -128, -128, -128, -128, -128, -128, 36, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 17, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -78, 127, -95, -128, -54, 127, -128, 7, -128, -128, -128, -124, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 11, 127, -128, -128, 127, -42, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -8, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 0, 127, 127, 127, -128, 127, 127, 127, 127, 127, -6, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -27, 127, 127, -32, 127, -128, 127, -128, -90, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -78, 127, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 8, -71, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -114, -128, -128, -128, -128, 93, -128, 127, 127, -128, -81, 127, 127, -128, 127, 127, 74, 127, 127, -128, 127, -128, 127, 127, -128, -91, 127, -128, -128, -128, -128, -15, 127, 127, -128, -128, -128, -128, -103, -21, 127, 127, 127, -128, 127, 127, -128, 127, 127, 65, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -52, 127, -128, -128, 127, -128, -128, 127, -128, -128, 11, -128, -128, 127, 127, -39, 127, 127, -128, -128, 127, -128, -128, -128, -128, 31, 127, 127, -106, 127, -36, 127, 127, -128, -128, -128, -128, 127, -16, 70, 127, 127, 127, 127, 92, -128, 127, -64, -128, 127, -119, 127, -107, 97, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 33, 127, -128, -128, -128, 50, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 86, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -90, 127, 127, 127, -128, -128, -128, -128, -128, 38, 127, -128, 127, 127, 127, 127, -128, -47, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -6, -37, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -13, 107, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 101, -128, -128, -128, -128, 127, -128, 127, 55, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 21, -128, 127, 127, 127, 127, 127, 127, 127, -78, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -23, 127, -128, 127, 127, 127, -128, 74, 127, -128, 90, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 28, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 5, -128, -128, -128, -128, 127, -128, -128, 53, -128, 127, 127, 10, -70, -128, -128, 127, 127, -103, 127, -128, -52, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -76, 127, 127, -128, -128, 127, -128, 68, 127, -128, 127, 127, 127, 109, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 7, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -108, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 3, 127, 127, -128, 127, 127, 127, -128, 31, -128, 127, 127, 127, 127, 55, 127, -128, 127, 127, 127, -118, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 10, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 6, -128, 127, 127, 127, -128, -128, -111, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 10, 127, 127, -128, 127, 127, -78, -128, 127, -128, -128, 127, -128, 0, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, -21, 127, -128, 127, 127, 127, 127, 127, 127, -6, -128, -128, 47, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -100, -128, -128, -128, -57, -128, -128, -86, -128, 127, -15, -128, 127, -128, -28, 127, -128, 127, 127, -128, 116, 127, -128, -128, 95, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -45, -128, 127, 127, -1, -128, -128, -128, -128, -128, -128, -91, 127, 127, 127, 127, 127, -116, 127, 45, -128, -128, 127, -28, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, 65, 127, 124, 127, 127, 123, -128, 127, 127, -128, 127, -128, -52, -44, -128, 127, 127, -128, 92, -128, -128, 127, -34, 127, 127, 127, 127, 127, 127, -128, -103, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -11, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 78, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 2, 1, 127, 127, -128, -128, -128, 127, -128, -5, -28, -128, 127, 127, 127, 127, -81, 127, 127, -128, 127, -65, -128, -128, -128, -128, -128, -128, 127, -128, 27, -128, -128, 127, -128, 118, -85, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -44, 127, 127, -128, 127, 127, -128, 2, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 23, 127, -128, -128, 127, -128, -128, 50, -128, -128, -128, -128, -128, 78, 127, 127, 127, 127, -128, -64, -128, -128, -5, -128, -128, -128, -128, -128, 127, 127, 127, 127, 18, -128, -128, 127, -75, -128, 69, -128, -128, -73, 79, 127, 127, 127, 127, 127, 106, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 116, -128, -128, -128, 127, 127, 92, -128, 39, -121, -128, -128, -128, 127, -128, 101, 97, -128, 127, 127, 127, -128, 70, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 18, -128, -128, -128, 91, -128, -128, 127, 127, 127, 33, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, -88, -128, -128, -128, -128, -128, -128, -128, -128, 5, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 121, -128, -128, 127, 127, 127, 127, -128, 127, 127, -18, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 112, 50, -128, -128, -128, -128, -128, -128, 127, 127, -63, -128, 63, -128, -128, 1, -128, -128, -38, -128, -128, 127, 127, 107, 38, -128, 127, 127, -128, 127, 127, -100, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 75, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -39, 127, 127, 127, -128, 24, 127, 100, 93, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -92, -128, 127, -55, 127, 127, -128, 127, 127, -128, -128, -18, -128, -128, 127, 127, 127, -128, -128, -34, 127, 127, 127, -26, 127, 127, 127, 127, 23, 127, -128, 127, 127, 127, 127, -103, -128, -128, -128, 127, 127, -128, -54, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, 88, 102, -128, -128, 127, -128, 79, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 108, 42, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -60, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 36, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -48, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -107, -128, 127, 127, -128, 10, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -44, 65, -128, 127, -128, -128, -128, -112, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 48, 127, 127, 127, -57, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 64, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 96, 127, -7, 127, -128, -128, -80, 127, 127, 127, 127, 127, -128, 127, -128, -128, 15, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 39, -128, -128, 58, 127, -128, 127, -128, 119, 127, -128, -128, 127, 54, -128, -1, 127, 127, 127, -55, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -98, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -74, 127, 127, 127, 127, -128, 127, -128, 95, -16, -128, 127, 127, -128, 127, 88, 127, 127, 127, 127, 127, 127, 127, 101, -128, -128, -128, -128, -128, -21, -128, -128, 127, -55, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -57, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -28, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 73, 127, -18, -128, -128, -128, -117, 127, 127, 127, 108, 127, 127, -128, 127, 127, -128, -128, -128, 26, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 68, -128, 127, 127, 127, 127, 10, -63, 127, 101, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 79, -128, 127, -128, -128, 13, 103, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 64, 127, 127, -64, -128, 45, -128, 88, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -10, -128, 127, 117, -128, 127, -128, -128, -28, 127, 127, -109, -128, 45, 127, -128, -6, 127, -128, 127, -128, -128, -128, -128, -86, -3, -128, -128, 119, 127, 78, 127, -128, 127, 127, 70, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -78, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -48, -128, -103, 98, -128, 127, -128, -128, 127, 127, 29, 127, 127, -128, -128, -128, 127, -128, -81, -71, -128, 127, -128, 127, 127, 127, 127, 127, 15, 127, 127, -128, 119, 127, 127, 127, 127, 44, -128, -128, -128, -128, -128, -128, -128, 127, -128, -122, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 0, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 2, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 55, 127, 127, -128, 69, 127, -128, -128, -128, -128, -128, -128, -128, -59, -128, -128, 53, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -18, -128, -128, 127, 127, -128, -128, -90, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -27, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 109, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -54, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -26, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 87, -70, -128, -66, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -54, 127, 54, 127, -128, -128, -128, -128, -128, -128, -73, -128, 127, 118, -128, 127, 127, -128, 127, -81, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -111, 127, -128, 127, -128, -128, 127, 127, 127, 24, 127, 127, 86, 127, -128, -128, -31, 127, 127, 127, 127, 127, -128, -128, 127, -128, 117, -128, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 33, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 80, 127, 92, -128, -128, -128, -128, 127, -128, 90, 127, -128, 127, 81, 127, -96, -109, -128, -128, 127, -128, 27, -128, -128, -128, -128, -111, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -78, 127, 127, 127, -60, 127, -95, 127, 127, 127, 127, -128, -128, -128, 127, -128, 80, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 17, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 28, -128, 127, -128, -128, 97, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 96, -128, -128, -128, 127, 127, -128, 127, 127, 57, 127, 127, -128, 127, -128, -47, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -93, -28, -128, 127, 127, -128, -24, 127, -128, 127, 127, -80, 127, 127, -128, 52, 127, -128, -128, -128, 127, -119, 122, -128, -128, 127, -128, -128, -128, -128, 127, 22, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 23, -128, 127, -128, 127, 127, 71, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -106, -128, -128, -128, -128, 127, 112, 127, 127, 127, 127, 127, -39, 127, 127, 127, -128, 2, 127, -128, 109, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 1, -22, 127, 127, 127, 127, 127, 127, 106, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -107, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -117, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -86, -128, -128, -128, -128, -128, -128, -95, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 59, -128, -36, -128, -128, -128, 127, -108, -128, -128, -128, 121, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 75, -128, -128, -128, -128, -1, 127, 127, -96, 39, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -2, -128, -128, -128, 127, -128, -128, 127, 106, 127, 127, -128, 127, 127, -128, -128, 127, -128, -70, 127, -128, -128, -10, -128, 29, 127, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 54, 127, 127, -128, -44, -128, 127, 127, 127, -128, -128, -33, -128, -128, -128, -128, -128, -50, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 71, -31, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -69, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -34, 127, 127, -27, -128, -128, 127, -128, 39, 127, -128, -128, -118, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 102, 127, 127, 127, 127, -15, -128, 127, -128, 127, -128, 95, 127, -128, 49, 127, 100, -128, 127, 127, 127, -128, -128, 127, 127, -54, -128, -128, 127, 127, -114, -128, 127, -128, -128, 127, 127, 127, 127, -44, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 49, -128, 127, 127, -96, 127, 127, 127, 127, 127, -128, -78, 127, 123, 28, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -79, 127, -128, 127, 127, -114, 127, 127, -21, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -116, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -103, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -114, -65, -128, -128, -88, 127, 127, 127, 127, 127, 127, -6, -38, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -63, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -23, -128, -128, -128, 127, -128, 58, 127, 127, -128, 127, 127, -88, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 88, 127, -85, 55, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 116, 127, 127, 93, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 70, -128, -128, -128, -128, -128, 100, 127, -39, 127, 127, -128, -128, 127, 127, 76, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 32, 127, 127, 127, -128, -128, 31, 69, -128, -128, -128, 127, 127, 75, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -38, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 117, 127, -128, -128, -128, 5, 93, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 26, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 97, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -108, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -16, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 63, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 10, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 85, -128, -128, 127, 31, -128, 127, -128, -128, -128, -128, -128, -128, -128, 91, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -37, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -69, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 28, 127, -128, -128, 127, 127, 127, -29, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -116, 127, -128, -128, 16, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -98, -128, 127, 127, -128, -63, -128, -128, 127, 66, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -53, 127, 112, -128, 127, 2, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -80, 127, 127, -128, -55, 75, 127, -128, 100, -128, -128, -128, -128, -128, -128, -128, 127, -36, -128, -128, 7, 127, -128, 24, 127, -128, -128, -52, 127, 127, 127, 127, 127, 127, -29, 127, -128, 95, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -49, 127, 127, 127, 127, 127, 58, 127, -112, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -100, -128, 63, 127, 127, 127, 127, 127, 127, 29, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -98, 127, -54, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 114, 91, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 10, 127, -128, -13, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -80, 127, -128, -128, 127, -128, 127, -22, -128, 127, 127, 127, 127, 57, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -23, -128, 127, 127, 117, 127, 127, 127, -18, 127, 45, -128, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -37, 127, 127, 127, 127, -128, 39, 86, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -97, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -32, -128, -128, 2, -128, -128, 66, -128, -55, 127, -128, -128, 127, 127, -128, -128, 78, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -68, -128, 127, 5, -128, 45, -128, -128, -128, 102, 127, 127, -128, 127, 127, 65, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -118, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 117, -128, -128, -128, 98, 127, 127, 127, 10, -128, 127, -128, 27, 127, -128, -73, -128, -128, 127, -128, -128, 95, -128, -128, -128, 127, 44, -128, 121, 127, -128, 127, 60, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 109, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -26, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -88, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -36, 48, -2, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 85, 127, -128, -128, 127, -128, -128, 127, -128, 64, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 18, -128, -128, -128, -128, -128, -128, -128, -128, -128, 96, -128, -128, 127, -21, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 24, 86, 127, 127, 127, -128, 23, 127, -12, 127, 127, -128, 127, -128, 90, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -12, 119, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -101, 127, 127, 127, 127, -128, -16, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -78, 127, 127, -128, 127, 127, 127, 127, -128, 7, 127, 118, 127, -128, 113, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 95, 127, 127, 127, -128, -128, -128, 127, -128, -98, 127, -128, 127, -128, -128, -128, -128, 127, -29, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 22, -128, -128, -27, -3, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -71, 13, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, 13, -91, 127, 127, 127, 127, 127, -128, -96, 127, 34, 127, -128, -128, -128, -128, 127, -128, 117, 127, -44, -29, -128, 33, 127, -128, 127, 127, 127, 127, 127, -32, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -114, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -1, 127, 127, 48, -128, 17, 127, 127, 127, 90, -128, 127, 79, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -80, 127, -22, 127, 127, -128, -128, -128, -128, -128, 127, 65, -128, -128, -128, -128, -128, -128, -128, -128, 45, -95, 127, -128, 127, 127, 127, 127, 127, 127, 78, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 38, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -107, -128, -128, 127, -128, -128, -109, 123, 127, -128, -1, -128, -128, 5, -128, -128, 127, 127, 127, 127, 127, 55, 16, -128, -128, -98, 127, 127, 127, 127, 127, 127, -128, 43, -128, -128, 127, -128, -128, 18, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -3, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, 49, -128, 127, -122, 127, -128, -128, -44, -128, -128, 127, -128, 122, 127, 127, 127, 127, 127, 127, 123, 127, 127, 114, -128, -128, -128, -80, 127, -90, 127, -128, -87, 127, 127, -128, 127, -128, 57, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -60, 127, 17, -128, 127, 127, 127, -128, -128, 127, -128, -128, 70, -128, -128, -128, -128, -128, 127, -64, -128, -128, 127, -128, 122, 127, 127, -128, -128, -128, -128, 127, 127, -88, 23, 127, 127, -128, -128, 127, -128, -128, -74, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 36, 127, 127, 127, 127, 127, 127, -128, 100, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -39, -65, 127, -128, -128, -128, -1, 127, 127, 127, 127, 127, 127, -128, -128, 127, -98, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 21, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, -68, 127, -128, 127, 112, 127, -128, 127, 127, -128, 127, 127, 127, -80, -128, -57, 12, -128, 127, -128, -128, 127, -128, -128, 127, -128, 123, -128, -128, 127, 127, -128, -88, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -111, 127, -128, 127, 127, -128, -128, 127, -87, -128, -128, -128, -128, 3, 127, 75, -128, 127, -128, 127, -128, 92, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 113, -128, 127, 127, 3, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 21, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -111, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 8, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 38, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -18, 85, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 32, -128, -103, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 102, -128, -128, 127, -128, -128, -128, -128, 127, -128, -92, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 114, 127, 127, 10, -128, -128, -128, -128, -93, 127, 127, -128, -128, -128, 127, 119, 107, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -68, 127, -127, 127, -128, -63, 127, -45, 127, 127, -128, -128, 127, -128, -128, 127, -128, 100, -128, -128, 127, -48, 127, -128, -128, -69, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 28, -128, -102, 127, -128, -128, -128, -128, -7, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 93, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -81, -128, -128, -128, -128, 127, 127, 127, -128, -128, -36, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 57, -128, -128, -128, 86, -128, -128, -128, -128, 127, 127, 127, 127, 127, 26, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, 127, 108, -128, -128, -128, -128, -128, 66, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 34, 127, 127, 65, -128, -128, -128, -128, 127, -128, -128, -128, -128, 0, -128, 127, -128, -128, -128, -128, -128, -128, 10, 127, 127, 127, 127, -128, 127, 127, -128, -128, 2, -128, -128, 93, -128, 127, 127, 127, -112, -128, -128, 127, -128, -128, 68, 127, 127, -88, -128, -128, -128, -128, 127, 127, 127, -119, 127, 127, 127, -128, 127, -17, 24, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 5, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 70, 127, 127, -128, -95, 127, -128, -45, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -74, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 59, -128, -128, 127, -37, -81, 127, 127, 127, -128, -128, -63, 127, 127, -128, 127, -128, 127, 127, 107, 127, -97, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -78, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -65, 127, 127, 60, -128, -128, -128, 127, 127, 0, -128, 127, 127, 127, 127, 127, 127, 127, 127, -97, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -21, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 127, 119, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -68, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 54, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -111, 16, -128, 127, -65, -128, 127, -128, -128, -128, -128, -123, -128, -128, 127, -44, 127, -128, -128, 127, -128, 88, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -91, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -81, 127, 127, -128, -128, -128, -128, -128, 127, 127, -69, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 45, 127, -128, -128, 127, 127, 127, 127, -128, 127, 79, -128, -15, 127, 127, 127, -102, -128, -128, 127, -128, -128, 127, -128, -128, 127, -87, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -60, 127, -128, -57, -128, -128, 127, 127, 127, -128, -128, -128, 127, -80, 127, 2, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 37, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 85, 127, 127, 127, -128, -128, -128, -128, -1, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 10, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -24, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 68, -128, -128, 127, 127, -128, -128, 127, -128, 102, -128, 117, 127, -128, -128, -128, -128, 90, 127, 127, -128, 127, 127, -128, 127, -128, 118, 127, -128, 127, 13, -128, 127, 127, -113, -128, -128, 127, -128, -128, -117, -128, -128, -128, 127, 127, 127, -128, 127, 127, 80, -128, -128, -128, -111, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 42, 127, 127, -128, -128, -111, -128, -128, 127, -97, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 119, -128, -128, 127, 127, -128, 13, 127, 127, -128, -128, -128, 127, -128, 127, 65, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 116, 52, -128, 127, -128, -128, -128, -128, -128, 64, 127, 127, -98, -68, -128, 127, 127, 21, 96, -128, 127, -128, -128, -128, -128, 27, 127, -128, -55, 127, 127, 127, 127, -124, -128, -1, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -96, -128, -128, -128, -127, 92, 127, 127, -128, 127, -128, -128, -128, 79, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -23, 81, -93, 127, 127, -128, -116, -128, -128, -128, -128, 127, -128, -128, 127, -128, 6, 127, -128, -128, -128, 127, 127, -128, -128, 118, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 121, 127, 127, 127, 127, 127, 114, -24, 127, 127, 127, 127, 118, -128, 127, 127, 127, 127, 127, 127, 48, -128, 127, -128, -1, -128, -128, 127, 127, -128, 127, 127, 127, 127, 23, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -38, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, 122, 127, 127, 127, 127, 127, -91, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -37, 127, 7, 127, 127, -128, -111, -128, -128, 127, 76, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 113, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -49, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 21, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 71, -128, -128, 102, 127, 127, 127, 109, 127, -128, 127, 127, 127, 127, 127, 127, 127, -102, -128, -128, -128, 127, 127, 86, -128, -128, -128, 127, 127, 127, 7, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, -128, -128, 32, 127, 70, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 109, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -39, -90, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 121, 127, -128, 127, -128, 127, 127, 127, 127, 28, -29, -128, 127, 127, 124, -128, -75, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 1, 127, 127, 127, 127, -128, -118, 127, -128, 127, -128, 111, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 21, 127, 127, 15, -128, -50, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 57, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -73, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 28, 127, -128, 106, 127, 127, 7, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -31, -128, -128, -128, 127, -128, -128, 127, 127, -85, -128, 68, -128, 127, 127, -128, -128, -128, -128, -128, -128, 100, 127, -128, -128, -128, 127, -128, -98, 127, 127, 127, -85, -128, -34, 127, -128, 127, 127, -128, 127, 11, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -107, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -13, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 65, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 26, -128, 127, 127, -128, 127, -27, -128, 127, 127, 127, 127, -128, -27, -65, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, 90, 127, -37, -128, -128, 127, 127, 127, -128, -15, -128, -128, -109, -128, -128, -22, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -53, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 114, 127, 127, 127, -123, -128, 48, 127, -128, -128, -90, -128, -128, -128, 127, 127, 127, -128, -128, 127, 98, -128, -16, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 27, 127, 127, 127, 127, 127, 112, -128, -128, -128, 17, -128, 127, -128, -128, 127, 18, -128, 127, 127, -128, -128, -128, -128, 127, -128, 127, 97, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 97, 127, 127, -17, -128, -128, -128, 127, -128, 127, 127, 102, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 34, 127, 127, 127, -128, -128, -128, 127, 127, -128, 122, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -71, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 39, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -64, 127, -128, 127, -128, -128, 127, -128, -128, -122, 127, -128, -128, 127, 127, -128, -75, -128, 81, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -69, -128, 127, -128, -128, -29, -128, -50, -128, -128, 127, -128, -26, 127, 70, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 54, 127, 127, -6, 127, 127, -128, 127, 124, 127, 127, 127, 7, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 47, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, -48, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 44, -128, -24, 127, 68, -128, -128, -128, -128, -128, -42, -18, 127, 127, 86, -128, 11, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 88, -128, 127, -128, -128, 100, -74, 127, 127, 127, 127, 127, -128, -86, -6, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 22, 127, -128, 97, -12, 127, -128, -128, 42, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -98, 127, -58, 127, 127, -128, -111, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 8, -91, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 18, 127, -97, 127, -128, -128, -128, 42, 127, 127, -128, -58, -128, -128, 127, -128, -128, -97, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -54, 127, 127, -128, -128, -128, -64, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 38, -128, -128, -128, -128, 127, 127, 127, -128, 100, -128, -128, -123, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -32, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 36, 127, -128, 127, 127, 127, 127, -128, -128, -128, 98, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, 34, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -87, -128, -128, 127, -128, -128, -128, -114, 127, -128, 127, -37, -128, -57, -128, -128, -128, -128, 127, -128, -128, 127, -128, -38, -128, 127, -128, -128, 127, 127, 127, 80, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 18, 127, -128, 127, -47, -128, 127, -128, -57, -128, -47, -128, -27, -128, -28, -128, 127, -128, -128, 127, -128, 127, 127, 73, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -87, 127, -128, 90, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 117, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 69, 127, -128, 127, -128, 127, 127, -128, 127, -116, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 57, 127, 127, -128, -128, -128, 127, 127, -128, 127, -55, 103, -128, -128, -128, -128, 127, 127, 127, 127, 79, 127, 91, -128, -128, -128, -54, -128, -128, 127, -128, 127, 127, -21, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 118, -128, 127, 127, 127, 127, -81, -128, -128, -128, -128, -128, -128, 127, -128, 60, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, -26, -128, -118, -128, -128, 127, -128, 48, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -66, 127, 127, 127, -128, -128, 127, -79, 127, 127, -128, -52, -128, -128, -128, 127, -98, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -124, 127, -128, -128, -128, 127, -128, -42, -128, -128, 127, -128, -29, 127, -88, 55, 127, -106, -128, 127, 127, -26, -128, -128, -7, 127, 49, 7, -128, -128, -128, -128, -128, 127, -128, -37, -31, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, -128, -1, 127, -128, -128, -128, -73, 127, 127, -103, 127, 127, -23, 127, -128, 112, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, 127, 92, 127, 127, 127, 127, 127, -47, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -12, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 88, 127, 127, 127, 127, 80, -128, 127, -88, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 108, 103, -128, -128, -123, 127, -128, -128, 127, -65, -128, -128, -128, 127, -57, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -44, -128, -128, -128, 127, -128, 127, -128, -113, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 10, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 28, 127, -128, 23, -128, -128, 127, 127, -128, -128, -128, 127, -70, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -24, 127, 119, 127, 127, 15, 127, 22, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -47, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 95, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 121, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 69, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -17, -128, -97, 127, 127, 127, 127, 49, 127, 127, 92, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 88, 127, 127, 127, 5, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 26, -128, 127, -128, -128, 74, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -112, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 17, 93, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 64, -128, -128, -59, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 45, 127, 127, 108, -128, 127, 127, -128, 127, 127, -128, -128, -21, 127, -128, -128, -128, -128, -128, -128, 127, -128, -80, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 78, 127, 127, -128, 44, 127, -128, -128, -5, -128, -128, -128, -128, -128, -128, -1, -128, -70, 11, 127, 10, -17, 127, -128, -128, 127, 127, -88, -128, -128, 127, 17, 127, 127, -128, 127, 127, 127, 127, -128, 127, -68, -15, -128, -128, 24, -128, -128, -128, -128, -128, -128, -128, 123, -128, -128, 127, 127, -128, -2, 127, 127, 127, 127, -128, -128, 127, 127, -128, -114, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 52, -128, -128, 127, -32, -128, 127, -128, 127, -128, -128, -124, 127, 127, 127, 127, 127, 127, -128, 127, 127, 48, 106, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 0, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, 127, -128, -55, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, -59, 127, 127, 127, 127, -122, -128, 127, -128, -128, 127, -128, -128, 127, 127, 111, -128, -47, 127, 127, 127, 127, -128, -52, 127, -128, -66, -112, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -43, -128, -128, -128, 127, 1, 86, 127, -128, 86, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -12, -128, 108, -128, -128, -128, 127, 127, 1, -128, -128, -128, -128, -128, -128, -28, -128, -128, -128, -128, -128, 127, 102, -128, -128, -128, 13, 127, -128, 127, -88, -128, 127, 127, 127, 127, -128, 111, 108, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, 119, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 37, -128, -73, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 79, 127, -128, 127, 127, 0, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 52, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 114, 127, 127, 127, 123, 127, -36, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 53, 127, -70, -128, -128, -128, -128, -128, -128, -128, -128, -128, -54, 127, -128, 24, -128, -128, 127, 127, 127, -55, 127, 127, -128, 127, -128, -128, -128, -2, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 8, -128, -128, -74, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -37, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 57, -121, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 106, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -117, -128, -1, 127, -128, -128, 43, -128, 127, 127, 79, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -36, -128, -7, -37, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -42, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -21, 127, 127, 127, 127, 127, -128, -128, 96, 127, 127, 127, 127, -128, -128, -128, -128, -69, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, -128, 127, -128, -113, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 27, -128, 127, -128, 127, 127, -128, -128, -128, 28, 127, -39, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 17, 127, 127, -128, -128, 127, 127, 127, 127, 127, -64, -128, 69, -128, 3, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 45, -38, -128, 127, 127, 3, 127, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 6, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -75, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, 15, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -108, 127, -128, 7, -128, 42, 127, 127, 127, 127, -128, -128, 127, -128, 28, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 59, -128, -128, 118, -128, -128, -128, 127, -128, -127, 127, -128, -128, 127, -76, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, -16, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -18, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -58, -128, -128, -128, 127, 124, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 111, -128, -128, -109, -128, -128, 127, -128, -128, 0, 127, 127, 127, 127, 127, 127, -128, -128, -6, 127, 127, 127, 127, 127, 113, 127, -97, -128, 127, -128, -48, -128, -128, -98, 127, 127, -128, -121, -111, 127, 127, 23, -128, -128, 127, -87, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 66, 127, 127, 127, 127, 13, -128, -79, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, 119, -128, -128, -128, -128, -128, -128, -128, -128, -50, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -6, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 12, -54, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, -73, 127, -128, 127, 127, -128, 127, -37, -128, 127, -128, -128, 127, 0, -88, -85, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -26, -128, -128, -128, -1, 127, -128, -128, -128, -128, -112, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -78, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -7, 127, 127, -128, -87, 127, -128, -128, 127, 123, 127, 127, -128, -45, 127, -128, -21, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -90, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -76, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -12, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 91, -128, -128, -102, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, -60, -128, -39, 127, 76, -128, 127, 116, -128, 127, 127, 127, 127, 127, -128, -113, 127, 127, 127, -128, -128, 127, 127, 127, 127, 52, -128, 127, -128, -128, -21, -128, -128, -128, -128, -91, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 16, -128, -88, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -64, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -85, 52, -128, -91, 127, -128, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 64, -128, -128, 127, -128, -128, 127, -128, -112, 103, 127, 28, -128, -128, 127, -128, 127, 127, -70, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 95, 127, 63, -128, 127, -128, -128, -128, -128, -114, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, 91, -128, 44, 127, 79, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -58, -121, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -11, 127, 127, 127, -128, 127, 127, -22, 127, -128, -128, -128, -128, 127, 127, 28, -128, 127, -88, -128, -128, -128, -128, 127, -128, 64, 127, -128, 108, -124, 127, 127, 127, 127, 100, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -68, -15, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -107, -128, 127, -128, -128, 18, 127, 127, -128, -128, -128, -128, 106, 127, -128, 127, -128, -80, 127, 127, -128, 32, 127, -128, 127, 127, -128, -128, -128, -128, -74, 100, -128, -116, 127, 127, 127, 127, 127, 127, 96, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -107, -128, 127, 127, 127, -106, 127, -128, -128, 127, -128, 127, -128, -128, -128, -2, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -65, 127, 127, 24, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -128, 114, -60, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 1, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 11, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, 121, -128, 127, -128, -128, 10, -128, 127, 127, 127, 127, -36, -128, -128, 127, -128, 78, 127, -128, 127, 127, 124, -128, -128, 127, 118, -128, -128, -128, -128, -128, -128, -128, 127, -31, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -100, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -95, -128, -39, 127, -128, -128, 127, -128, 127, 127, -128, -91, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 103, -128, -128, -128, 85, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 107, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 29, 116, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -109, -128, 127, -128, -128, -128, -107, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -112, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -50, -90, 127, 127, 127, 127, 127, -128, 127, -128, 22, 127, 85, 127, -128, -128, 127, 127, 127, 127, 127, 55, 127, 16, -128, 127, 127, -128, -60, -68, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 69, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, -96, -128, 127, -98, 127, -128, -128, 127, 49, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -73, -128, -88, 127, 75, -128, -128, 26, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -37, -128, -128, -128, -128, -128, -128, -55, -114, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -98, 119, 127, -128, -128, -128, -36, -103, -128, 127, 127, -111, -128, -128, -128, 127, -128, 92, 127, -128, 127, 127, -24, 127, -54, -128, -128, -87, 116, -128, 127, -36, 127, 127, -128, 127, 58, -128, -128, -128, -128, -128, -128, -128, -68, -128, -128, 127, -128, -128, 69, 127, -39, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 36, 127, 127, 127, 127, 127, 113, -128, -128, -128, -128, -128, 127, -128, 127, 28, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 69, 85, 127, 127, 127, -117, -91, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -109, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -85, -65, 127, -60, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -95, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 127, -128, -91, 127, -128, 127, 127, -128, -96, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 122, -128, 127, 127, -128, -128, -128, 34, -116, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -112, -128, -128, -128, -128, -128, -128, -113, 107, -128, -128, -128, -128, 127, -128, -98, -128, 127, 127, -128, 127, 127, -128, 42, -128, -128, -54, 127, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, 60, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -80, 127, 103, 100, -128, -128, -128, 127, 96, 127, 127, 127, -128, -128, -128, -128, -71, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, -49, -128, -128, 127, -128, -128, 127, 127, -128, 127, -78, -93, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, 116, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, 11, 127, 127, 127, 127, -128, -28, 127, -18, 64, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, -79, 127, -128, -128, 127, -128, -128, 127, 102, 127, -33, 127, -128, -69, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -80, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -29, -128, -128, 127, -128, 127, 127, -10, -128, 127, 127, 127, 127, -128, -128, 127, 95, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -57, -128, -128, -128, -128, -128, -128, -128, -21, -37, -128, -128, -128, 127, 127, 127, 68, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -33, 127, 127, 127, 127, 127, -128, -102, -128, 116, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 118, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 13, 127, 127, 45, -128, -128, 127, 127, -55, 127, 127, -128, -128, -128, -128, -128, -128, -128, 8, 127, 127, 127, 127, 127, 111, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 6, 127, -128, -27, 127, 127, -22, -26, 127, -75, -128, -128, 127, 127, 127, 123, 127, 127, -128, -128, 127, 63, -128, 127, 127, 127, -31, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -98, 127, -128, 118, -102, -128, 127, -128, -85, 127, 58, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, 29, -128, 127, 127, -128, -128, -128, 127, 127, 127, 38, 127, -128, 127, 127, 127, 127, 127, -128, 44, 127, -128, -128, -128, -128, -128, -128, 127, -47, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -124, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -106, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -7, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 18, 127, 127, -128, -128, -128, -128, -128, 57, 28, -128, 127, -128, -128, -128, -128, -128, -21, 127, -128, -103, 127, -87, 127, -128, 122, -128, 39, -128, 127, 127, -3, 127, -128, -128, -128, 127, -128, 127, 127, -128, -44, 127, -128, 97, -128, 127, 127, -128, 127, -128, -128, -18, 127, 127, -128, 127, 127, 127, 127, -128, 127, -22, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -63, 127, 44, -128, 127, -128, -128, 127, -128, -128, -128, -45, -128, 127, 127, -128, -128, -128, 127, 127, 127, 12, -128, 127, 127, -128, 127, 127, -128, 79, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, 96, -128, -128, 127, -128, 127, -101, -128, 127, -38, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -7, -6, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -92, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, 127, -13, -128, -128, -128, -128, -49, 127, 127, 127, 127, 27, -128, 127, 127, 109, 127, 127, 127, 127, -128, 127, 81, 112, 91, -85, -5, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 123, -128, -128, 39, 127, -128, -33, 127, 127, 127, -128, 96, -128, 127, 127, 127, 127, -128, 127, -59, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 44, -128, -128, 127, -128, 36, 127, 127, 127, 127, -128, 127, -55, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 100, -128, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -55, 127, -128, 127, 127, -128, 127, -128, 18, 8, -128, 127, -23, 127, 127, 127, -68, 127, 127, -128, -128, -128, -128, -128, 119, -128, 127, -128, -128, -128, -128, 127, -128, 127, 127, -87, -128, 127, 127, -128, 36, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -112, 127, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -70, 127, 127, 127, 127, -21, -128, 127, 127, 127, 127, 127, 127, 127, -128, 44, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 33, 127, -128, 127, -128, 85, 127, 127, 127, 127, 31, 127, -128, 127, 127, 127, -128, 127, -128, -128, -128, -128, -128, 65, 127, 127, 79, -128, -128, -128, -128, 127, -128, 127, 127, 34, 127, 127, 112, -59, -128, 127, 127, 127, 127, -128, 127, 124, 127, 127, 114, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 11, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -52, 127, -128, -128, 127, -91, -128, 96, -128, -128, -128, -128, 127, -70, 127, 127, 63, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -113, -18, 127, 127, 127, 127, 127, 127, -128, -128, 49, -128, 127, -128, 127, 127, -123, 127, -128, 127, 127, 127, 127, -128, -109, 127, -128, -128, 127, 127, 92, 127, 127, 47, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -76, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, -128, 65, -128, 127, -128, -128, -128, 127, -128, 60, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -45, 108, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, 65, -98, 127, 0, 127, -128, 93, 127, -128, 127, 127, 127, -128, 127, 127, 127, 12, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, 127, -36, 127, 127, 127, 127, 127, 127, 127, 6, -128, 78, 127, -128, -128, -26, -128, -128, 127, 127, -128, 88, 127, -128, 18, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, 16, -128, 127, -128, -128, -128, -128, -128, 26, -128, 127, 127, -128, 47, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 74, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -55, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, 0, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, -69, -128, -128, -128, -128, -128, -128, 127, -88, 127, 127, 13, -36, 127, -39, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, 116, -128, -128, 127, -128, 76, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -29, -128, -128, -128, 127, -128, 127, 127, -122, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -79, -128, 127, 106, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -93, -128, -128, -128, 127, -6, 127, 127, -128, -74, -96, -128, 127, 127, 31, -128, 52, 127, -128, -128, 127, 127, 127, 127, 127, -128, -13, 127, -128, 127, 127, 127, 127, -38, -128, -128, 127, 127, -21, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -39, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -5, 127, 127, 127, 85, -128, -128, -128, 60, -128, -24, 127, 127, 29, 127, 127, -128, -128, -70, -128, -111, 127, -128, 127, 127, 127, -107, 6, -128, 45, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 70, -128, -128, -87, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 0, 127, -124, -128, 127, -128, 97, -128, -128, 127, 127, 127, -48, -128, -128, -128, -128, 127, 127, 64, 127, 127, 127, 70, 107, 127, 127, 127, 127, 127, 127, 127, 127, -97, -128, 127, -128, -128, -29, -128, -128, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 22, -128, -128, 127, -128, -128, -49, -128, 127, 127, 103, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, -6, 127, 127, -114, -128, 127, -128, -128, 127, 127, 127, 127, -128, -111, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 107, 127, 127, -111, -128, -128, -128, -128, 12, -128, 22, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 10, -128, -128, -128, -128, 58, -128, -128, -128, -91, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, -1, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -80, -128, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -10, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 57, -128, 127, -101, -128, -128, 127, 127, -128, -28, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, -36, -128, 49, 68, 127, 127, 127, 127, 127, 127, 98, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, 127, 127, -123, -128, -128, -128, -128, -128, 106, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 6, 127, -128, 54, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -39, 127, 127, 127, 127, -5, -128, 92, -128, -128, -81, -128, 127, 127, -65, 127, 127, -54, 127, -128, -128, 127, -128, 127, -29, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 28, -128, 127, 127, 127, 127, 127, 127, 127, 127, -44, -128, -128, -128, -128, 127, 127, 127, -55, 127, 127, 127, -128, -128, -128, -21, -128, -128, -128, -128, 127, -128, -98, 127, -128, -128, -128, -128, 0, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -91, -128, 127, 127, 127, 28, 127, 127, 127, 127, -128, -128, -128, 127, 34, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -64, 127, 127, 27, 127, -128, -128, -128, -128, -128, -128, 95, 127, -128, 127, 127, -128, -128, 127, 49, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -117, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, 2, -128, -128, 117, 127, 127, 127, 127, -128, -90, -128, -128, 127, -38, 69, 127, 127, 127, 127, 55, -128, -128, -128, -128, -128, -128, -39, 127, -128, 127, 127, -113, -128, 60, 127, 127, 127, -69, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, -36, -128, -128, -128, -128, 127, -128, 57, 24, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, -112, -128, -128, 127, 127, -128, -128, -128, -128, 42, -128, 23, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, 103, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 93, -123, 127, -128, -128, -128, -128, -128, -128, 80, -128, 127, -128, 127, 127, 127, -128, -128, 127, -5, 127, 127, 7, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 127, -39, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 11, -128, -128, -128, -128, 127, 127, 127, 127, 100, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 100, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -109, -128, -128, -128, 118, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -44, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, 127, -27, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -70, 127, -128, -36, 127, 127, -128, -128, -128, -128, -128, 127, -48, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 90, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 52, -128, 124, -128, 127, 127, -128, 127, -128, -128, 127, 78, 127, 127, 127, 127, 127, 127, 127, -22, 127, 127, -128, -8, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 124, -128, -128, -128, -128, 127, -128, -128, 57, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -6, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 26, 127, -128, -128, -128, -86, -63, -92, 127, 127, 127, 127, -32, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 5, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -114, 127, 127, 127, 127, 127, -86, 8, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 47, 127, 127, 127, -128, -128, 85, -128, 107, 127, 127, -128, -128, -128, 11, 127, 127, 127, 127, -24, 127, -128, -128, -128, -128, 127, -3, -128, 127, -128, 127, 127, 127, -128, -128, -65, 127, -128, -116, 127, -5, -128, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 79, 127, 127, 63, 127, -128, 127, 127, 127, 127, 127, -128, 127, 87, -128, 127, 127, 127, 127, 127, -128, 127, 127, 81, 127, -128, 127, 127, 127, 127, 127, -10, -128, 127, 127, 127, -128, 108, -70, -3, -95, -128, 127, -112, -128, 127, -128, 127, 16, -128, -7, -128, -128, 95, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -27, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -128, -128, 79, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, -13, 127, -128, -128, 127, 80, 127, -128, 42, -128, -128, 127, 127, 127, -128, -128, 118, -128, -128, 127, -128, -121, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 34, 127, 127, 127, 127, 127, -128, -44, -128, 127, -128, -128, -3, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -117, -128, 127, 127, 127, -128, -128, 127, 127, -70, 127, 127, 127, 12, 127, 127, -128, -128, -128, -12, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -101, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, -128, -65, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 1, 127, -128, -128, -128, 127, 127, -128, 113, 127, -63, 127, 127, 127, -128, 127, 127, -128, 37, 127, 127, -128, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -26, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, 121, 127, -128, 127, 127, -128, -128, 39, 127, -128, 7, 127, -44, 66, -128, 127, 118, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, 127, 127, -54, 49, -39, -128, -128, 16, -128, -128, 124, 127, 127, 127, 127, -128, 127, 71, 127, 127, 127, 127, -128, -128, -64, -128, -128, 127, -69, -128, -128, 127, 80, -128, 127, 127, -128, -128, -128, -128, -50, 127, 127, 127, 127, 81, -128, -128, -128, -128, -128, -128, -128, -128, 12, 127, -128, -128, -128, -128, -128, -128, -128, 73, 127, -128, 127, -128, -128, -2, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, -128, 127, 127, -52, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -71, -53, -29, 127, 127, 127, 127, -128, -128, 127, 127, 13, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -81, 127, 127, -128, 127, 111, 127, 127, -128, 127, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -2, -128, -128, -128, -128, -111, -128, 127, -53, -128, -128, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, 127, 95, -128, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 71, -76, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, -128, 127, -128, -128, 127, -44, -128, 80, 68, -128, 127, 127, 127, -128, -128, -128, -118, -128, -128, 55, 127, 127, -128, 127, 127, 127, -128, -128, 127, -49, -128, -128, -128, -128, 127, -78, -52, 127, 127, 71, 86, 127, -128, -128, 127, -86, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 127, -98, -128, 127, -128, 127, -71, -128, 127, 127, -128, 127, -128, -128, -128, 127, 21, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -28, -128, -128, 127, 127, -128, 127, 127, -128, 27, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -11, -12, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -69, -128, -128, -128, -92, -5, 127, -128, -128, 127, 127, 108, 127, -128, 8, 127, -128, 127, 127, -128, 0, 127, -128, -128, -128, 127, -128, -128, 127, -128, -16, 102, -128, -128, -128, 127, 127, 127, 127, 127, 127, -54, 127, 127, -128, 127, -128, -128, -128, -128, -128, -128, 127, -128, -128, 127, 32, -128, 87, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 87, 127, 127, 127, 127, 127, -128, 127, -90, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -109, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, -93, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, -27, 127, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, 49, 23, -128, 127, 127, 127, -128, 127, -38, -128, 127, -128, -128, 127, 101, 127, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, 127, 127, 71, 127, 127, 127, 127, 127, -128, 53, 127, 127, 127, -128, -57, 127, -128, -128, 127, -128, -128, 36, 127, -39, -128, -128, -128, -65, 127, 127, -128, 127, -128, -128, 127, 112, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -6, -128, -128, -128, 102, -128, 96, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, -34, -128, -128, -128, -128, 127, -16, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 100, 127, 127, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -44, -128, 127, 127, 127, 34, -128, 127, -112, 127, 127, -128, 127, -128, -128, -28, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -48, 87, -5, -128, 127, -128, -29, 127, 127, 127, 127, 127, 127, -128, -128, 127, -128, -48, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, 47, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -52, 127, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -66, 127, -1, -52, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, 127, 127, 127, 127, 127, 127, -27, -128, 127, 127, 69, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 3, -128, -128, -128, 127, -75, -128, 48, -128, -128, 127, 127, -128, -128, -108, 127, -128, -128, 127, 127, -128, -31, 127, -128, 49, 127, -128, -128, 127, 87, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 28, 127, -128, -128, 127, 6, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 24, 127, 127, 121, 127, 127, -128, -58, -128, -128, 127, -106, 127, 127, 127, 127, -27, 127, -128, 127, -128, -128, -128, -128, -128, -128, -128, 127, 0, -128, 127, 31, -128, -128, -128, -128, -128, -128, -111, 127, 127, 127, 127, -128, 127, -98, -128, 127, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 34, 127, 127, -128, -128, -128, -128, -128, -17 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
