-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            108, 104, -76, -80, 9, 70, -13, -115, -108, 17, -62, 78, -3, -88     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -119, 2, -23, -81, -57, -91, -34, 74, -55, 106, 93, 14, 51, 111, -45, -97, -102, 70, -56, 79, 55, 59, -58, -126, -66, 117, -16, 38, 6, 44, 35, 16, -68, -39, 82, 63, 113, -125, 13, 67, -70, -28, 93, 50, 61, -27, -124, -39, -61, 17, 59, 44, -117, -1, 99, -37, 18, -69, 43, 8, 11, 108, -122, 62, 19, 55, -64, 75, -47, -108, -127, 84, -70, 80, -22, 18, -114, -115, -61, 119, -94, 22, 105, -19, -3, -104, -90, 37, -97, 29, 30, -75, -113, -116, -77, 82, 120, 49, 17, -35, -21, 77, -40, -83, 116, -60, -23, -106, 13, 83, 114, -124, 114, -16, 117, 14, -73, -93, 35, -35, -111, 60, 17, -16, 19, -34, 61, -20, -118, 95, 41, -8, 111, -127, -4, -51, -68, 97, 52, 121, 17, -115, 4, -116, -30, 71, 97, 11, 86, 72, -83, 49, 10, 48, -88, 125, -35, -59, -75, -4, -96, -83, 53, -94, -28, 65, -64, 52, 13, -90, -60, 46, 56, 18, 81, -44, 101, 52, 97, -29, 127, -12, 69, -75, -1, 59, -109, -33, 104, -40, -6, 126, -108, -45, 88, 122, 41, -53, 22, 82, -116, -13, 94, -79, -83, 118, 92, -54, -24, -96, 46, 90, 57, -52, 36, 50, 56, -85, 62, -108, -71, 5, 80, 10, 29, -47, -49, -28, 105, -123, -23, -77, 10, -20, 100, -74, 96, -72, 17, -88, 83, 73, -73, 87, 82, -89, 79, -115, 88, 62, -91, -20, -16, -28, -65, -80, -4, 114, -93, -6, -45, -57, 13, 80, 10, -70, -128, 54, -35, 101, -1, -14, 35, -51, 90, 127, 49, 88, 53, -127, 76, -104, -61, 6, -76, 39, -97, -92, 26, 37, 102, -31, -17, 100, 18, 64, -4, 38, -125, -48, 43, 42, -89, 4, 33, 93, -17, -92, -6, 89, 15, 74, -36, -109, 84, 83, 6, -123, 42, -108, -124, -111, -10, -50, 86, -1, -95, 5, 0, 23, -7, -109, 105, -118, 30, -37, 116, 15, -101, -96, 111, 43, 27, 54, 123, 65, 35, -29, -104, -1, 42, -37, -108, -17, 11, 67, -12, 118, -38, -27, -123, -79, 9, -26, 43, 21, 80, 22, -38, 98, 107, -114, 101, 46, 27, 100, 63, 99, 9, 36, -25, -57, -30, -69, 72, -45, -109, -53, 54, -14, 39, -36, -15, -47, -34, -15, -80, 88, 38, 82, 105, 64, -39, 45, 39, 55, 51, 83, 42, 106, 118, -84, 41, -77, -29, 28, -87, -12, 74, -40, 86, 7, 85, -79, -47, 39, 40, 76, -113, 81, -46, 10, -127, -25, 123, -7, 66, 96, 93, -50, 106, -64, 3, 34, 1, -5, 113, -36, -127, 74, 39, -111, 87, 58, 113, -77, 121, -115, 118, -53, 33, -32, -77, -73, -8, -58, -74, -1, -53, 27, 35, -126, 91, -61, 66, -120, -94, 25, 119, 67, -25, -33, -102, 74, 85, 58, 33, -81, 44, -72, 17, 26, -52, 29, -68, -112, -14, 69, -3, -40, 37, -1, -54, -124, 27, 46, -93, 101, -98, 40, -91, 126, 92, 84, 41, 69, 108, 109, -18, 61, 114, 10, 27, 127, -48, 21, -37, 71, -6, 30, 31, -63, 23, -110, -47, -80, 127, 105, -6, -63, -51, -25, 35, 47, 17, -34, 114, -49, -116, -21, 61, 10, 9, 27, 112, -100, -104, 92, 76, -109, -57, 49, 11, -112, 30, -63, -95, 117, -6, -41, 47, 23, 59, -74, 108, 54, 125, -46, -122, -86, 55, -3, -49, 83, -118, -116, -67, -68, -22, 8, -58, -14, 28, -109, 51, 19, -109, -6, 52, 5, 74, -94, 101, 38, -5, 99, -2, -85, -73, -70, -55, -87, 53, 112, -71, 92, -106, 27, 122, 4, -12, 103, 17, 100, -120, 22, -86, 74, -116, -23, 28, 83, -77, -43, -102, 46, 64, 40, 37, -44, -102, 81, 121, 120, -87, 12, -76, -125, -126, 112, 18, 86, -55, -63, 127, -32, -54, -110, -71, 42, 82, -16, 68, 27, 54, -13, 10, 43, 104, -41, -63, 64, 21, -41, 1, -106, 27, 109, 45, 43, 81, 110, 50, 46, -30, 58, 83, 87, -120, -57, -125, -115, -33, 12, -93, 45, 61, 64, -27, 28, 29, 119, 65, -30, -50, 0, 32, -96, -20, 44, -62, -96, -103, -9, 55, 51, -95, -44, -57, -65, 126, -106, -68, -110, -49, -18, -92, 125, -108, 104, 104, -67, 54, -100, 108, 23, 1, -100, 61, 104, 35, 100, -42, 62, 71, -5, -49, 25, -8, -125, -34, 35, 68, -74, -7, -109, -35, -119, 118, 14, -114, 121, -61, 124, 72, -52, -19, 54, 70, 73, 108, -57, -119, -61, -118, -5, 63, 104, 51, 28, -78, 84, 54, 12, -101, -9, -23, -111, -13, 97, 44, 3, -73, 23, -81, -82, -60, 17, 65, -68, 8, -65, 98, -48, -28, -95, -115, 115, 80, 59, 27, 105, -9, 53, 86, -110, 83, 15, 127, 118, 102, -114, 2, 18, -89, -40, 71, -5, 54, 83, 15, 63, -87, -90, 113, -36, -9, -65, 79, 119, 85, -17, -44, -119, 87, -97, 15, -98, -38, -75, 1, -109, -84, 71, -93, 34, 59, -87, -83, 61, -107, 97, -43, -86, 32, 109, 5, 117, -73, -57, 0, -8, -48, 28, -84, -59, -24, -16, 121, 75, -93, -48, -122, -84, 49, -124, 98, 92, -11, 7, 31, -121, -112, 57, -109, -110, 39, 78, -111, -68, 23, -115, 6, -1, -46, 52, -8, 85, -126, -50, -89, 79, 106, 52, -123, -125, -67, -11, 59, -64, -33, 110, -101, 33, 103, -39, -108, -72, -107, -41, -48, -98, 110, -87, 16, 92, -125, -121, 21, 7, 5, -24, 126, 37, 118, 92, -70, 85, -54, 49, -66, -63, 122, 93, 15, 49, 121, -19, 7, 80, -60, -19, -87, 47, 118, -10, 78, 1, -43, -54, 47, -65, 105, -41, -81, -18, -94, 34, 76, -76, 99, -33, 107, -85, 89, -17, 127, -82, 14, -41, 19, 122, -74, 99, -110, -90, 32, 94, -108, 105, 97, 33, -127, 54, 93, -127, -89, 8, -98, -87, 53, -124, 5, 35, -89, -94, 92, 102, -88, -63, -33, -100, -102, -3, 15, 84, -78, -7, 0, -10, -78, 93, 80, -55, 70, 66, 56, -52, -82, -20, -91, -41, -76, 46, 118, -87, 23, 14, -93, 68, 2, -3, -28, 86, -102, 11, 0, -41, -61, -37, -93, -84, -8, -105, 121, 15, -120, 73, 45, 70, 91, -3, 70, 44, 112, 73, 30, -43, -46, 61, 67, 109, 28, 98, 79, 74, 34, 44, 81, -92, 123, -75, -59, -38, -29, -86, 21, -13, -7, 12, -117, 25, -128, 21, 73, -35, -109, -62, 26, -24, 24, 103, 82, 5, -71, -118, -89, 87, 57, 97, 76, 41, 29, 18, -4, 106, -106, 7, 0, 25, 67, -78, -125, 98, -39, -52, -32, -66, -84, 47, -4, -70, 12, -35, 74, 9, -30, -9, 11, 0, 61, 93, -26, 95, 112, -31, -73, 91, -88, -27, -97, 80, -59, 120, 57, -113, 66, -50, 18, -43, 29, 29, 90, 115, 92, 0, 113, 106, 72, 109, 106, 24, -40, -97, -68, -116, -120, -73, 4, 79, -30, 24, -52, 68, 67, 90, 86, -62, 127, 44, 54, 21, 111, -107, 68, -38, -65, -98, -125, -110, 26, 49, -11, 11, -103, 32, -109, 17, -25, -60, 27, -82, 84, 127, 23, 16, 5, 30, 95, 35, -84, -31, -73, -29, -48, -8, 97, 48, 81, -45, 41, -15, -100, 75, -38, 41, -52, 50, -117, 94, 7, -35, 46, -17, -36, 95, 32, 102, 11, -38, 53, 37, -39, -105, -43, 3, 30, -30, -1, -91, 85, -79, -16, 86, -99, -48, 22, -57, 75, 27, 54, 79, 97, -69, -119, -45, -61, -44, -75, -14, -93, -21, 60, -17, -99, 81, -11, 81, -4, -75, 87, -93, 79, 118, -19, -90, -123, 98, 51, 86, 39, 101, 88, 16, 57, -57, 26, -69, -4, 61, -104, 60, 72, -82, -14, -78, -76, -46, 42, 106, 108, -55, -67, -101, 40, -114, 127, 10, -23, 56, 102, -121, -81, -47, 31, -6, -24, -75, -105, 53, -3, -21, 29, 108, 53, -28, -50, -30, 52, 39, -26, 74, -112, -56, -85, 12, -99, 33, -80, -4, -3, 60, 15, -39, -38, -115, 61, -66, 51, 20, 121, 82, -27, -70, -112, 86, -75, -108, 107, 97, -24, -2, -120, 66, 21, 77, -120, 27, 82, -44, -108, -29, 27, -5, 114, 16, 102, -12, 63, 12, -29, 5, -21, 26, 76, -109, 116, -101, -95, 92, 27, 72, -20, -4, 125, -69, -90, 66, -43, 82, 30, -87, 85, -111, -2, 39, 57, 36, 77, 40, 60, 92, 41, 102, -61, 101, 65, -25, -41, 53, 117, -13, -91, -121, -126, -47, 118, -120, -90, 88, 33, 123, 120, 73, -10, 32, -100, -55, -7, 13, 72, 73, -45, 120, -73, -60, -100, -111, 60, 11, 49, -9, -96, 5, -116, 18, 127, -80, -66, 70, 5, 15, 57, -45, 64, -53, -20, 112, -84, -73, 84, 2, 109, -38, 0, 21, 70, -28, 65, -80, 58, -9, -13, 72, -59, -32, -106, 19, 11, -100, 7, -60, -57, -113, -54, -24, 26, -25, -1, -21, -48, 18, -112, -63, -63, 18, -3, -12, 61, -78, 48, -123, -24, 105, -65, -23, 124, 24, 124, -91, -83, 103, -20, -68, -2, 110, 56, 61, -59, 9, -11, 61, -80, 8, 54, -120, -43, 100, 91, 48, 57, -115, -111, 6, 119, 74, 54, 110, 110, -92, 98, 87, 31, -31, -56, -123, -72, -63, 84, 28, 63, 79, -82, 35, -91, -6, 4, 5, 8, -92, -19, 63, -22, 99, -122, 3, 116, 80, 26, -80, -35, -122, -109, -111, 49, -43, 115, 14, 106, 79, 60, 99, 38, -46, 73, -26, -79, 68, 116, 65, -58, 68, -34, -99, 55, 118, 79, 46, -21, -61, -36, -62, 5, -60, -82, 56, -118, -112, -75, 31, -49, -38, 123, -31, -55, -96, -46, -53, -50, -27, 22, -80, -105, 11, 29, 88, -110, 2, 21, -31, 110, 97, -89, -119, 58, 58, -85, 55, -14, -20, 98, 35, -11, -68, -54, -111, -92, 79, -115, 83, 107, 37, -31, -81, 42, -105, 110, -44, 73, 47, -75, 78, -53, 117, -62, -68, 40, -92, -27, 117, -32, 23, -119, -107, -84, -115, -86, 110, 111, 63, -59, 121, 100, 4, 114, -23, -115, -118, 120, -125, 49, -128, 83, 35, -30, -38, 81, 70, -22, 44, -84, -116, 82, -54, 65, -50, -23, 123, 105, -121, -30, -67, 50, -23, 82, -72, 43, -117, 60, -5, -50, -34, 94, -81, 51, -11, 24, -112, 10, 70, 44, 23, -61, -117, 75, -97, 102, -7, -54, 95, -42, -95, -39, 48, -67, 98, 96, -48, 42, 40, -6, -98, 17, -82, 74, 18, 35, 90, -31, 5, -90, -119, 92, -127, -42, 64, 15, -122, 92, 60, -70, -61, 87, 55, -1, 119, -24, -56, 125, 3, -112, -113, 77, -93, 37, -65, 23, -27, 62, -42, 106, -11, -23, -105, -75, -43, -65, 36, 50, 10, -30, 13, 95, 62, -65, -81, 113, 75, 119, 118, 57, 44, -53, 32, -58, -115, 7, -123, 2, -51, 74, -114, 16, -108, 41, -33, 19, 37, 69, -115, -42, 127, 111, -95, 33, -9, 101, 68, 98, 15, 6, -21, -70, -65, -85, -34, 120, 64, 65, -12, -96, 104, -9, 49, 94, -94, -46, 126, 54, 38, 86, 3, -101, 4, -85, -51, -104, -15, 81, 65, -97, 99, 97, 61, 28, -96, 18, -99, 70, -27, -23, -46, 19, 68, -53, -51, 34, 99, -45, -87, 37, 25, 49, 89, 15, -110, 72, -65, -79, 44, 35, -38, 89, 55, 92, -119, 117, -93, -94, -32, -124, 61, -46, 11, 85, 62, -3, 92, 44, 111, 103, 124, -5, -6, 18, -5, -10, -113, 25, -6, -120, 26, 33, -122, 108, 97, -43, -17, 47, 8, -17, 30, 59, -60, -61, 13, -46, -118, -35, 7, -105, 2, -118, -70, 118, 26, -120, -45, -118, 17, 113, 7, -57, -108, -119, 123, 24, -20, 18, 114, 47, -32, 109, 68, 28, 91, 117, 38, -71, 25, -45, -54, -29, -30, 82, 59, -120, -126, 58, -26, -37, -109, 48, -48, -123, -108, -74, -16, -75, -78, 32, 55, -77, 56, -49, -33, 81, -33, -68, -31, -33, -124, -54, 19, -59, -83, -96, -12, -57, -65, 60, -111, -90, -18, -1, 112, 70, -23, 126, -64, 30, -75, 113, 111, -114, -105, -104, 21, 61, 78, -67, 70, 55, 20, -8, -102, 103, 102, 109, 16, 109, -5, 1, -96, -107, -11, 57, 115, -83, -89, 59, 47, 104, -112, -63, 15, 21, -68, 60, -126, 81, 74, -14, -111, -126, 99, -83, -11, 54, -96, 39, 20, 70, -103, 72, 124, -128, -54, 71, -13, 37, 35, -57, -55, -94, 109, 73, 123, 108, 86, -124, 73, 43, -103, 39, -117, 29, 58, -70, 94, 101, -74, 46, -81, -3, 40, -61, 108, -117, 51, -39, -79, -23, -107, -95, 51, 62, -53, 73, 87, 107, 27, -62, -89, 12, -52, 88, 33, 111, -48, -97, 113, -54, -85, -112, -46, -125, 41, 70, 77, 60, -121, 97, 103, -92, -27, 14, -100, -93, 92, 86, 82, -105, -112, 65, -98, -57, 5, 64, -1, 2, 66, -106, -53, 116, 46, 78, -11, -86, -43, 57, -23, -67, 66, 123, 19, -119, -126, 46, 50, -38, -97, 33, -86, 3, 121, -42, 18, -125, -10, 15, 96, -72, -77, 50, -102, -67, 93, 46, -89, 58, 82, -38, 12, -128, -4, -117, 25, 49, -29, 94, -62, 42, 39, -74, 41, -124, 43, -13, 5, 62, -122, 11, -15, 30, -101, 74, 18, -53, -112, 74, 69, 106, 120, -126, -1, -11, -35, 112, 62, 118, -97, 42, -31, 52, -46, -92, 94, -90, -128, 103, 3, -69, 86, -33, -112, -44, -27, -96, -119, 112, -50, -46, 2, 81, 48, -39, -65, 80, -108, 62, -64, 50, -97, -19, -7, 61, 125, 69, -24, 69, 127, 40, -105, -69, -121, -112, 49, -92, 33, -10, 4, -24, 25, -96, -63, -54, -15, 0, -113, 92, -43, 71, -60, -62, -107, 21, 7, -28, -31, -68, -73, 31, -14, 87, -32, 45, -36, 62, -119, -80, 47, -108, 74, 85, 89, -107, -23, 29, -128, 89, 50, 50, -43, -17, -51, -123, 91, -98, -113, 114, -84, 18, -63, 114, 45, -42, 101, -8, 5, 107, -10, -47, 59, -96, 65, -121, -73, 32, 4, -79, 127, -12, -63, 70, -85, 10, -62, 123, -33, 7, 114, -69, -77, -57, -128, 51, 85, 92, 48, -48, -96, 65, 42, 108, -98, -36, -44, 120, 39, 23, -4, 3, 71, 97, -62, 37, 93, 1, 79, -125, -7, 71, 112, 81, 94, 7, 99, -66, -120, -10, 113, 41, 68, -51, 89, 18, 109, 21, 88, -66, -60, 33, 106, -107, 60, 4, -6, -29, -118, 44, 103, -111, 91, 39, 104, 47, 86, -46, 36, -85, 54, 17, -47, 101, 115, 49, -47, 80, -1, -30, 39, 38, -38, 52, -59, -16, -111, -97, 83, -85, 62, -91, 47, 82, -6, 60, 42, -116, 79, -42, -59, 40, 55, 108, 125, -114, 54, -91, -13, -60, -23, 122, 20, 31, 19, -91, -85, -12, 19, -31, 59, -13, 78, -114, 13, 77, 14, 67, -62, 31, -67, 21, -72, 95, -84, 4, -104, 47, -86, 123, -33, 103, -10, 88, 97, -71, -44, -104, -128, -62, -72, -19, 15, 115, 52, -104, 97, -126, -21, 40, -4, -107, 116, 76, -83, -111, 125, -47, 43, 78, 72, -54, 57, -24, -24, 67, 21, 55, 127, -101, -42, -32, -22, -125, 68, -114, -90, -35, 30, 1, -37, -43, -59, 114, 118, 51, 0, 64, 92, 109, 38, 85, 36, -4, -91, 21, 67, 40, 19, -112, -98, -6, 15, -6, -123, 2, -117, -35, -99, 26, -28, -63, 0, 99, -119, 79, 114, -14, 88, -23, 59, 57, 50, 104, -127, 104, 92, 22, -63, -23, 81, 94, 25, -27, -108, -90, -2, -1, 32, -51, 94, 67, -31, 35, 78, 48, 24, -110, 80, -6, 9, 15, 69, 57, 20, 37, 90, 36, -55, -111, -56, 54, -108, 109, 124, 99, -12, -24, -114, -95, 61, 126, 123, 96, -83, 77, -58, -8, -118, -88, -51, 83, -10, 39, -124, -32, -77, 92, -63, -7, 38, -28, 6, 46, 71, 92, -22, 68, -76, -16, 19, 38, -64, 63, 73, 94, -13, -66, 33, 82, 28, -120, -58, 21, -87, 30, -35, 120, 91, 107, 108, -108, 90, -97, 6, 96, 82, -69, 97, 33, -46, -36, -124, -64, -119, 76, -20, 118, -71, -52, 96, 80, 90, -52, 86, 93, 121, -3, 22, 90, 59, -114, -9, 9, 73, -43, 50, 65, -9, -107, -58, -39, -38, 15, 28, 37, -100, 62, -63, -73, 111, 89, -101, 99, 13, 71, -125, -83, -49, -117, 22, 78, -29, 6, 115, -87, 48, -98, 87, -85, -128, -85, -61, 97, 58, 123, -109, -90, 116, 10, 81, 91, 24, 59, 76, -104, 100, -6, -56, 81, -68, 57, -54, 107, 8, -100, 48, 107, 14, -122, -111, 7, 103, 69, 17, 22, -66, -125, 24, -75, -16, 43, -118, 117, 124, 68, -44, 73, -74, -43, -122, 2, 37, 28, -119, 10, 36, 87, -1, -85, -83, 16, -64, -13, -49, 117, 76, 120, 103, -1, 65, 86, -87, -84, 20, 40, -113, 125, -20, 12, 58, -77, -112, 60, -53, 115, 40, 14, 53, 50, -35, -68, -107, 46, -16, 12, 40, -107, 65, -36, -76, 120, 66, 25, 46, -104, -65, -55, -94, 64, 33, -13, -5, 115, -45, -37, 26, -64, -81, -1, 16, -116, 65, 82, -45, 34, 14, -96, -83, -122, 62, 5, -84, -6, 34, 114, 68, -81, 54, 60, -10, 124, 19, 109, 117, 41, -78, -85, -92, -66, 35, -100, 11, 41, -16, -7, 78, 73, -93, -92, 29, -27, 120, 87, -28, 40, -5, -12, 113, -108, 114, 41, -93, -73, 46, 66, 39, 89, -117, -84, -17, -40, 110, 61, 69, 32, 71, -28, 50, -47, 87, 1, -126, 76, -108, -122, -46, 106, 107, 81, -86, 61, -13, 94, 9, -12, 57, 1, 9, 99, 33, -94, 9, -92, -17, 86, 85, 46, 17, -89, 13, 36, -97, 58, 43, -102, -36, 78, 48, -6, 39, 119, -16, 2, -46, -122, 39, -28, -96, -71, 115, -88, 38, 64, 10, -107, 74, 121, -58, -64, 30, 80, 119, 114, 116, -65, 81, -88, 16, 31, 16, -121, -54, 94, -6, -81, 8, 94, -113, -125, -56, 78, 89, -54, -51, 44, -89, 6, 77, -22, 46, -116, 67, 44, 63, 87, 86, -92, -22, -16, -108, 72, 64, -3, 21, -87, 70, -114, -58, -105, -108, -43, -101, 119, 58, -87, -10, 125, 117, -100, 43, -47, 81, 123, 104, 52, -60, -2, -72, 6, 43, -124, 52, -12, 96, -128, 86, -76, -81, -94, -53, -90, 108, 114, -4, 2, -125, 34, -23, 51, 67, -16, 96, -125, -126, -59, -3, 94, -84, -47, -124, -8, 42, -71, 124, -50, 54, 94, -8, 68, 85, -23, -8, 105, 30, -41, -89, 87, -83, 117, 23, 58, -101, 125, 126, 94, -27, -75, 63, 4, 56, -93, -99, 93, -86, -72, -117, -41, -54, 38, 68, -65, 40, 5, 113, -45, 52, 127, -55, 36, -88, -46, 108, -45, 13, 21, 33, -106, 70, -127, 56, 81, 104, -82, 51, 110, 123, 79, 106, 77, 94, -44, -35, -91, -35, -115, 116, -120, 81, -103, -86, 121, 72, 23, -103, 73, 74, 8, -108, 2, 76, -13, -53, -60, -92, -27, 90, 15, -122, 11, -58, -32, 102, 91, -128, -81, 22, -86, -84, -80, 22, 41, 105, 42, -122, -73, -49, -57, -74, 93, -102, -10, -62, -61, 127, 54, -26, 17, -34, 5, 107, 83, -66, -89, 22, 0, 49, 25, 102, 42, -77, 98, 17, 34, -90, -120, 54, 45, 9, 38, 27, -2, 97, -23, 88, 3, 96, -65, 67, -61, -75, -77, 86, 67, 40, -9, 82, -83, 103, -19, -93, 12, -33, -4, -38, 76, 107, 39, 102, -84, 55, 124, -77, 108, -25, -96, 17, -7, -114, -66, -95, -64, -21, 85, 24, -68, 4, -11, -27, -110, -62, 6, -49, 44, 12, -23, 46, -120, 82, 106, -28, -126, 123, -27, 44, -29, -68, 14, -32, -81, -106, 25, -2, -17, 94, -3, -69, 0, 109, -52, -33, 113, 74, 9, 89, -93, 79, 43, 73, -6, 51, 125, 32, 97, -88, 127, 1, -116, -128, -71, -89, 111, 6, 82, -21, -45, -34, -26, 16, -47, -62, -76, -21, -118, -69, 54, 64, -72, 81, -18, -9, 81, -12, 0, -38, 13, 85, 17, -116, 16, -39, -85, -71, 126, 45, 1, 73, -33, 2, -51, -45, 112, -59, -56, 63, 5, -28, 35, -45, 3, 20, 63, -99, 21, 24, -52, 19, 87, -95, -67, 41, -43, -72, 116, -51, -73, -26, 23, 50, 74, -69, 71, 85, -83, -49, -69, -28, 19, 49, 1, 85, 79, 87, -63, 8, 43, -51, -110, -47, -80, -66, -69, 121, 106, -11, 58, -59, 28, -2, 61, -107, -109, 47, 111, -23, -70, 33, 25, -15, -92, 75, -90, -41, -70, 125, 89, 60, 35, -103, 9, -67, 106, 47, 11, -52, -77, 93, 58, 5, -14, 97, 3, -79, -54, 12, -26, -34, 115, 103, 55, -5, 119, -86, 88, 87, 87, -95, 103, -125, 127, -92, 19, 113, -65, -7, -116, 71, 31, -43, 26, 21, -109, -33, -18, -34, -74, -52, 38, -128, 75, 79, -5, -121, 62, -33, -25, -63, 71, -34, 34, -7, -24, 107, -11, 93, -73, -48, 12, 21, -126, -63, -101, 114, -50, 38, -101, -82, -106, 32, -37, -79, -28, -102, 31, -50, 75, 38, 104, -48, -4, 32, -116, -15, 110, -64, -62, -33, -21, -51, 98, 30, 118, 21, 56, -54, -117, 36, 4, 32, -41, -20, -81, -18, 90, -32, -24, -25, -25, -125, -108, -59, -96, 85, -120, -65, 50, -15, 96, -106, -52, -53, -102, -44, -33, -79, 52, 106, -46, -43, -53, -77, 3, 9, -72, 18, -89, -119, 109, -123, 118, -102, 64, 116, 82, 103, -91, -96, 30, -65, -2, 124, 113, 90, 48, 18, -6, 32, -80, -115, -1, -9, 92, 97, -49, -18, -38, 74, 68, 121, 22, -77, -92, -53, 89, 57, -16, -44, -49, 53, -55, 92, -41, 54, -101, -35, -50, 11, 44, -79, -7, -123, 115, -89, -76, 61, -113, 57, 106, 102, 79, -97, 11, -103, -108, -128, -29, 20, -84, -77, 73, 54, 12, 122, -60, 65, -103, -125, 114, 110, -107, -41, -4, 102, 34, 118, -26, -121, -106, -103, -121, 55, -105, 37, -74, 54, 114, -33, -76, -37, -88, 57, 121, 72, 49, -62, -41, 68, -116, -49, 29, -95, -73, 123, -27, 19, -10, -65, 102, -81, 90, -45, -67, 78, 78, 50, 112, 101, -115, 95, 50, 27, 77, -44, 44, 9, -107, 10, -81, -105, 47, -55, -47, 104, -28, 50, -46, -13, -75, 77, -119, -8, -49, -79, -47, -8, -14, 40, -69, -77, 99, -28, 126, 107, 49, 92, -70, 10, 44, 75, -41, 86, -29, 127, -60, -76, -121, 26, 83, 60, 24, 17, -44, -89, 108, 113, 18, -95, 47, -54, 64, 58, -40, 122, 127, -24, 62, -78, -33, 7, -74, 100, -84, 81, -111, -72, -79, 82, -48, -17, 48, -106, -39, -67, 32, 53, 60, -93, -127, 76, -48, -87, 109, 26, -52, -7, -34, 28, -69, -101, -17, 94, -109, 55, -22, -121, -21, -33, -53, 118, -4, 63, -119, 88, 63, -125, 67, 77, 17, 34, -96, 117, 52, 59, -127, -112, -5, 66, -97, 58, -51, -127, 111, -122, 63, -38, 28, 74, -128, -32, -123, 42, 113, 94, -122, -29, 127, -69, -126, -14, -44, -55, 107, 97, 49, 51, 56, -50, 77, 121, -18, -21, -87, 109, 5, -109, -84, -99, -72, -128, -9, -8, -48, -16, 19, 1, 68, 68, -37, 98, -23, 25, -58, 34, -6, -79, -43, 35, 62, 65, 82, 6, 20, 6, 33, -56, -107, 94, -68, -75, -74, 96, -75, 98, -22, -17, 98, -48, 40, -39, -99, 79, -47, 100, 115, -124, -7, -59, 34, 79, 28, 30, 75, 18, 78, 96, 104, -17, -12, 27, 104, 15, 79, 45, -128, -20, -96, -35, 104, 67, 18, -1, 96, -103, 117, 49, -89, 125, 83, -70, -123, 3, 30, -105, 98, 41, -20, 47, 12, -34, -109, 101, -105, -109, -77, -32, 107, 12, 62, -44, 57, -36, -67, 40, 26, -32, -56, 36, 85, -111, 56, 90, -33, 40, 114, 68, -40, -87, 113, -42, -54, 34, -16, -8, 7, 122, -38, -95, 121, -20, -73, -26, -42, 37, -122, -95, -96, 12, 96, 106, 54, 115, -79, 26, -9, -9, -4, -109, -45, -5, 108, 118, -29, 113, -1, -32, 65, -42, 114, -87, -25, 73, 19, 89, -87, -111, -50, -120, 115, -14, 22, -112, -115, -25, 69, 47, -87, -35, 121, 64, -90, 23, -66, -120, -76, 33, -106, -52, 2, 124, 13, 71, 32, 33, -20, -50, 122, 38, 80, -13, 11, 76, 122, 69, -30, 21, -22, -26, -94, -114, -24, -126, 9, 10, 70, -81, -25, -87, -7, -20, -46, 118, 6, 2, -24, -45, -102, -111, 29, -119, -17, -62, -24, -120, 56, 101, 103, -9, 67, 51, 70, -35, -66, -84, 111, -24, -109, 9, 52, 103, 79, 1, 24, 8, 27, 107, -53, -60, -28, 32, -26, -116, 76, -82, 81, 77, -76, -119, -64, 92, -110, -24, 45, -47, 29, -41, 20, -84, 93, 121, 51, -105, 76, -81, 120, -109, -65, 101, -72, -74, 21, -46, -64, -2, -118, -104, -64, -101, 110, -111, 68, 52, -5, 108, -94, -122, 12, -33, 9, 42, 18, -12, -30, 54, 44, 120, 127, -4, 81, -123, 76, -68, -110, 125, 53, 53, -6, -44, 116, -38, -22, 70, -8, -80, 54, -120, -103, 119, -79, -128, -18, -94, -12, -65, -114, 36, -42, 74, -5, -87, -93, -96, -116, -105, 20, 95, 106, -9, -23, 94, -96, 124, -57, -63, 106, 15, -33, -36, -52, -66, 48, -84, 53, 29, -115, 68, 7, -83, 116, 72, 8, 88, 54, -24, 29, 4, -88, 42, -121, 50, -107, 127, -54, -84, 79, -71, 40, 105, 102, -88, -117, 71, -51, -109, -73, 105, 71, -126, -91, -10, -127, 78, -3, 96, 8, 70, -55, -35, -72, -124, 34, -87, -40, 82, 102, 127, 123, -1, -8, -13, 67, 39, -71, 51, -112, -113, 93, -51, 43, -7, 77, -29, 27, -116, 26, 74, 94, -48, 93, 71, 4, -73, -44, 3, 38, 45, -19, 44, 90, 36, -29, 63, 124, 16, -98, 78, 7, -91, -28, 38, 32, -43, -22, 111, 84, -109, -65, 12, -96, 43, 118, 93, -31, -110, 110, 16, -72, 123, -10, 76, 62, -53, 124, -118, -117, 50, -77, 52, -124, 65, -66, 55, -101, 1, -53, -73, -22, -77, 106, -78, 30, -45, 13, -57, -92, 5, -87, -74, 87, 97, 67, -40, 12, 10, -70, -44, -110, -109, -101, -58, -95, 103, 63, 23, -104, -49, 77, -76, -70, -116, 29, 4, -76, -81, 81, -11, 106, 47, -28, 97, -44, 26, 31, -126, -103, -60, -44, 54, 66, -75, -103, 127, 101, -108, 98, 41, -126, -72, 5, -98, -85, 78, 67, -38, -48, -123, -13, 35, 60, 89, -54, 25, 55, -40, -104, -90, 97, 74, 42, -94, 45, -106, -18, -54, -75, 17, -55, -74, -105, -64, 30, 47, 122, -8, 97, 30, 113, 117, -20, -32, -17, 89, 122, -13, -59, -83, -119, -66, -33, 29, 108, 102, 67, -74, 77, -74, 105, -108, -124, -61, -93, 91, -49, 88, 89, 72, 34, -76, -11, 97, -101, 14, -46, -13, -34, 66, 117, -84, 37, -33, 53, -58, 68, 82, 78, -15, -52, -44, -22, 101, -66, 33, 48, 6, 102, 82, -24, -35, 58, -83, -5, 66, -8, -51, 9, 124, -29, -91, -128, -128, -126, -70, -20, 41, 15, 10, -123, 76, 88, 74, 109, 102, -96, -83, -30, 109, 104, -82, -89, -38, -29, 27, 121, 41, -9, -67, -111, -4, -7, 82, -127, 56, -109, 80, 107, 88, 50, 54, 19, -86, -115, -8, -14, -111, 118, -82, -79, -13, -18, 120, -32, -128, 107, 66, 82, -24, 99, -94, 65, 17, -67, -45, -122, -93, 9, 84, 51, 5, 52, 62, 120, 90, -99, -2, -113, 78, 124, -70, 29, -2, 90, -36, 48, 71, 15, 69, -43, 127, -124, -68, 79, 79, 3, 84, -122, -84, 69, -112, 124, 51, -85, 125, -16, -41, -121, 76, -19, -106, -46, 115, 86, 101, -49, 63, 76, -42, 23, -67, -83, 77, -10, 115, -35, 36, 43, 21, -126, 23, 106, 53, 54, 42, -32, 109, -118, 64, -59, -94, 106, -37, -77, 15, -57, 17, -28, -79, 16, -99, 60, -3, 54, 9, 81, -71, 60, -20, -112, 85, 73, -9, 89, 21, -58, 77, 99, 102, -80, 60, 77, -49, -118, 27, 95, 109, -114, -118, -32, -103, 61, -94, -90, 30, 53, 124, 45, 60, -40, 96, -71, -48, -3, 43, -18, -27, 35, 120, -54, -51, -95, 63, 118, 113, 0, -70, 57, 59, -47, -110, 18, -96, -114, 52, 45, 43, 87, -19, 42, -39, 87, -24, 117, -79, -102, 15, -29, -3, 126, -81, -63, 120, -115, 61, 118, -63, -99, -21, -49, 99, 84, 124, -19, -69, -75, -44, -90, -8, 117, 43, -82, 30, -64, 1, 0, 101, 98, 33, -63, 89, -66, 57, -82, 4, 41, 83, -22, -1, 84, -28, 20, -31, 12, 9, 122, 85, 101, -35, -107, -103, 83, 59, 35, -33, 108, 105, -6, 11, -119, -113, 35, 125, -108, 108, -92, -124, 27, -84, -125, -31, -126, 29, 54, -1, -18, 50, 53, 89, -73, -93, 1, 40, 32, -7, -98, -8, -111, -118, -65, -49, 50, 63, -77, 76, -56, -101, -26, -95, 98, -89, -59, 71, 16, 57, 45, 52, -27, 8, -21, 11, 1, -15, -97, -10, -12, 20, 26, 0, -125, -54, 80, 35, -62, 15, 120, -20, 99, 106, -46, -88, 25, -24, 68, -114, -93, -61, -90, -111, 59, -16, -31, 101, 57, 60, -35, -14, 8, -81, -100, 124, -19, 12, -1, 11, 124, -14, -105, -34, 51, -86, -25, -54, 49, -116, -114, 119, 66, 97, -46, 85, 62, -126, -66, 44, 126, -92, -83, -106, 79, -48, -90, 12, 48, -9, 44, -76, 62, -5, -105, -109, -103, -119, 41, 97, -91, -79, -46, 16, -108, 105, -28, -122, -128, -34, 100, -36, 91, 25, -75, -68, 41, -46, 32, 43, 56, -124, 110, -17, 126, 28, -44, 111, -59, 28, -123, 39, 104, 39, 11, 49, -69, 17, -100, -38, -127, -72, 62, 80, 59, 60, -127, -94, 58, -43, 23, 72, -15, -71, -81, -11, 31, -52, 108, 36, 66, -9, -126, -107, 33, 95, 117, -71, -56, 1, 71, 60, -95, -123, 87, 52, -55, -95, 58, 102, -89, 52, -51, 120, 15, -15, 4, -115, 5, -53, 68, 6, 25, 87, 2, 20, -31, -30, -97, 80, -122, 0, -125, -111, 113, -24, -85, -78, 102, -36, 94, 122, -34, 36, -7, 83, 85, 97, 92, 42, -79, -106, 120, -112, 93, 70, -43, -1, 31, -26, -37, 18, -17, -94, 97, -25, 107, -85, 66, 65, -6, 30, -5, -101, 88, -61, -18, 37, -90, -85, -7, 48, -113, 126, 40, 4, -3, 15, -57, 51, 18, 7, -101, -37, -125, -87, 127, -126, -22, 88, 102, -40, -9, 122, 10, 89, -62, -49, -21, -23, -107, 110, 123, 29, 72, 61, 88, 23, -56, -58, 29, -19, 104, 60, -78, -90, 58, -30, 6, 18, 75, 8, -88, 25, -60, -124, -88, -26, 101, 56, 25, 104, 56, -123, 103, -85, -39, 36, 106, 93, -93, -47, -12, 6, 70, -34, -17, -91, 98, -13, -71, 92, -91, -31, 95, -68, 119, -116, 39, -101, -123, -91, -117, -44, -39, 77, -6, 116, -82, -12, 35, -28, 117, -100, 37, 78, -35, -48, 99, -69, 16, 42, -23, -28, -104, -88, -10, -66, -34, 93, 95, -31, -25, -67, 59, 68, 96, -96, -11, -21, 33, -17, -94, -84, -123, 45, 33, 99, -62, -75, -42, -93, 25, 58, 33, -8, 88, -118, -48, 34, 35, 11, -89, -21, -37, 23, -2, 74, -66, -54, -76, -5, -37, -64, -5, -17, -68, 121, -90, 18, -116, 26, 13, -128, -113, -61, 64, -75, 32, -32, 35, -65, -50, -31, -23, -40, -77, 100, -60, 123, 19, -80, 125, -47, 42, -109, -34, -64, 31, 112, -69, 4, -10, 56, -110, 12, 72, -4, 70, 1, 59, -95, -101, -49, -37, 23, -76, -21, 52, -53, 111, 4, -60, 81, 117, -113, -87, -42, 1, 56, 52, -74, 42, -23, 29, -98, 35, 115, 78, -84, -33, 79, 87, -30, -54, 81, -4, 15, -20, -49, -12, 76, -25, 113, -88, 32, -65, 88, 17, -97, 78, -74, -40, 119, 84, 112, -48, 34, -55, 24, -71, -56, -37, -7, 22, -59, 117, -68, 72, -9, -54, -40, -50, -62, 120, -101, -52, 29, -100, 69, -16, -33, -40, -121, 116, 61, 38, 59, -125, -86, 20, 120, -29, 2, 124, -85, -104, 111, 8, 40, 121, -65, 16, 114, -61, -69, 65, 103, -104, -110, -2, -37, 28, 104, 70, -75, -82, 12, -29, -91, -40, -63, 73, -12, 3, 90, -7, -12, 87, 40, 36, 68, -111, 108, -102, 93, 67, -116, 74, -91, -24, -29, -113, -120, -8, -96, 40, -1, -57, 83, -45, -51, -57, -76, 33, 44, 45, -78, 42, 12, -18, 81, 48, 93, -13, -45, 7, -69, 45, -65, 17, 88, 113, -17, -64, -113, -8, -29, 123, 22, 64, 63, 74, 0, -43, 82, 68, -47, -68, 35, 48, -94, -33, 61, 66, -123, 104, -77, 91, 31, -42, -10, 76, -10, 31, 68, -41, -104, 57, 75, 11, 96, -29, -13, -56, 15, -122, -23, -11, 96, 6, 122, 40, 62, -43, 125, 97, 63, -24, -29, -1, -1, -4, 109, 37, -43, -14, 7, -111, -94, 64, 115, 27, 124, 0, 63, -108, 6, -63, -43, 107, 38, 1, -20, -125, 16, 101, 59, -108, -37, -74, -76, -75, -53, -26, 97, -10, 58, 53, 93, -120, 5, 104, -122, -40, 75, -13, 126, -117, -41, 108, -122, 8, 94, 52, 83, 105, 52, -18, 36, 80, 124, 94, 101, -80, -120, 53, 38, -51, 121, -82, 68, -25, 113, -94, -80, 68, 46, -10, 107, -8, -119, 28, 117, 124, 114, -120, -30, 116, 0, 104, -21, -58, -71, 68, 51, -67, 25, 48, -22, 29, -88, 105, -1, -46, 59, 18, 118, 54, -111, 49, 109, 19, 114, 42, -90, 99, -108, -87, -17, 100, -102, -104, 95, -11, 90, -79, -5, 3, 40, 85, 44, -37, -95, 99, -65, 14, 107, 82, -44, -10, 109, 48, 122, -125, 117, 91, 32, -75, 28, 46, -19, 66, -10, -83, -56, 108, -44, -126, -99, -57, -53, 75, -34, 68, 37, -84, 29, -117, -127, 29, -127, -65, -80, 21, -15, -12, 71, 19, -5, 80, 97, -69, 12, -52, -24, 57, 6, 73, 62, 7, 54, 42, 46, 40, -28, -64, -63, 127, 9, 0, -73, 110, -51, 25, 104, -24, -97, 46, 110, -52, 80, -6, 15, -116, -14, 29, -95, -31, -17, -24, 5, -55, 20, 86, 39, 52, 21, -70, -101, -10, -36, -36, -2, -2, 47, -95, -74, 50, 57, 40, 63, 22, 83, -54, 115, 2, 56, 12, 19, 54, -35, 32, -59, 52, -86, 9, 18, -42, 56, 44, -75, -100, -98, -76, -116, -7, 23, 61, -32, 92, -58, -106, 100, 84, 89, 118, 103, -28, 34, -102, 71, 11, -61, 89, -10, -47, 36, 96, 17, -102, -34, 91, -13, 86, -25, -127, 85, -3, -44, 103, -26, -11, -96, -27, -34, -90, -21, 26, -98, -87, -48, -51, 32, 66, 62, 77, 15, -56, 107, 59, -19, 26, -100, 44, 84, 107, -29, -60, -100, -72, -1, 120, 46, 38, -30, -118, 32, 78, 73, -2, 111, 85, -73, -40, 9, -31, 61, -42, 36, 8, -108, -92, 30, 63, -43, 19, -48, -20, 90, 28, 67, -38, -59, 1, -109, 49, -63, -83, 7, -121, 51, 3, -57, -97, -3, 92, -38, 27, 93, -13, 19, -103, -119, -92, -101, 104, 24, -30, -18, -3, 93, -75, -28, -66, 7, -13, -103, -61, 117, 74, 13, 82, -78, -68, 84, -80, 17, -86, 37, -49, 30, -61, -71, 118, 78, 27, 0, -120, 87, -102, -6, -122, -81, 97, -15, 101, 51, 116, 96, 7, 14, 61, -122, 83, -112, 63, -85, -24, 59, 23, 103, -70, 5, 69, 13, 4, -67, 102, -45, 47, 86, -89, -14, 9, 9, -100, 84, 11, -107, -47, -91, 85, -66, 88, -105, 87, 119, 79, 23, 17, 94, -92, 110, -120, 113, 98, -93, 54, 31, 44, 83, 99, -30, -108, 70, 24, -118, 41, 16, -126, -123, 1, 41, 100, -111, 110, -5, -115, -78, -68, 63, -24, -17, -97, 110, 98, -83, 37, 50, 124, 3, 79, 119, 75, -116, 5, -7, 102, 107, 92, -93, -8, 120, -94, 93, 91, 84, -17, -55, 106, 79, 102, -7, 68, 88, 17, -112, -27, -21, -83, -67, 79, 28, 46, 26, 127, 93, 71, -99, 42, -37, -49, -5, 1, -92, 24, 104, 106, -2, -15, -125, -54, -118, -127, -63, 65, -91, 102, -85, -38, -9, -99, 15, -8, 67, -90, 2, -101, 13, 112, -98, -108, 72, -31, 68, 36, 68, 97, -71, 26, 51, -120, -99, -70, 56, 51, -115, -40, 72, 5, 59, -33, -36, 127, -82, 68, -83, -109, -59, 63, -118, -27, 77, -61, 27, -125, -114, -10, 1, 12, 110, -110, 39, -6, -106, 21, 40, 127, 122, -111, -40, -128, -1, -18, 112, -10, 76, -121, 127, -123, -41, -120, 40, 2, 84, 28, -44, 11, 100, -58, -39, -19, -57, -28, -5, 86, -52, -40, -73, -10, 61, 85, -23, -5, -51, -102, -43, 120, -18, -110, -13, -29, -52, -76, 118, 52, -92, -114, -1, -17, -60, 69, -69, 26, 59, -99, 27, -35, 8, 122, -22, -59, -123, 4, -42, -104, -96, -48, -102, 85, -6, 20, -117, -82, -37, 17, 60, 110, -45, 59, -98, 109, -9, -77, -39, -39, 78, -95, 7, 125, 52, 30, -98, 91, -80, -38, 62, 65, -74, 90, -51, -60, -75, -99, -101, 103, -56, -37, 99, -96, -111, -70, -115, -100, 101, -25, 101, -52, -45, -102, -62, 103, -20, -22, 15, -73, -67, 59, 55, 0, -98, 70, 10, 45, 96, 100, 118, 123, 114, 37, 68, 28, 71, -4, -54, 24, 91, 47, -64, 2, 53, 0, 89, -93, 49, 110, 20, 67, -112, -101, 99, 7, -115, 125, 104, 45, -116, 84, 112, -50, 95, -118, 47, -100, -126, -114, -67, -86, 2, -80, 101, 46, -38, -30, 61, 95, 73, 71, -96, 87, -95, -110, -20, -115, -100, 14, 2, -19, -126, -15, -78, 48, -31, 123, 28, 61, 68, 88, 118, -11, -76, 50, 88, -47, 64, 45, -10, -117, 42, 117, -124, -74, -13, 88, -29, -39, 15, -75, -122, -121, 108, 99, 124, 24, 51, -105, -96, 107, -14, -57, -3, 44, -80, -114, -15, 75, -62, -120, -98, -25, -14, 63, -82, -29, -5, 76, 127, -7, 8, -22, -102, -100, 76, -117, -26, 23, -75, -94, 18, -102, -103, -29, 42, 89, 119, 22, 11, 115, 28, 0, -20, -66, -15, -44, -18, 17, 55, 36, 111, -109, 6, -126, -29, -114, 66, 14, 21, 81, -15, 24, 35, -93, 17, 114, 105, -69, 108, -74, -34, 53, -107, 82, -75, 30, 117, 120, -85, 30, -75, -37, -123, -103, -11, -5, 93, -70, -5, -122, -125, -53, 121, -103, -19, 19, -51, -38, 86, 35, 95, -109, -108, -99, 98, 81, 34, -31, 3, 32, -38, 108, 13, -26, -42, -95, 57, 18, 9, -86, 114, -6, -4, -39, 52, 105, -110, -125, 101, -70, 12, -9, 64, 51, -28, 116, -109, -81, -61, -106, 115, -51, 93, 51, 37, 6, 113, -103, -23, 92, -48, -79, 34, 123, -5, 25, 68, 37, 44, -117, 98, 13, -91, 33, 43, 28, 107, 19, -61, -72, 39, -118, -55, 30, 34, -96, -79, 47, -87, 90, 24, 126, 20, -80, 87, 102, -112, 87, 106, -86, 127, -99, -17, 78, 0, -87, 71, 80, -70, -31, -40, 125, -91, 28, -52, -125, 111, -63, -30, 46, -47, -111, 34, -6, -114, 119, -46, 104, -80, 5, 11, -89, 4, -36, -38, 111, -53, -98, -111, 42, 76, -90, -55, -32, -20, -123, -10, -122, 20, 40, 83, 8, -116, -81, 74, -22, -58, -39, 72, 8, -41, 38, 110, -107, -28, -4, -91, 20, -5, -24, -98, 106, 33, -76, 114, -106, -29, -97, -107, 6, 59, -45, 33, 83, 48, 34, -66, 82, -57, -66, 95, 43, -26, -39, 83, -21, 53, 23, 106, -14, -76, 51, 85, -115, -59, 19, 29, 115, -1, 84, 48, 53, -76, 54, 30, 38, -97, 110, 103, 121, -36, 48, 62, 42, 79, 102, 84, -74, -110, 57, 122, 51, -18, 85, -42, 39, -128, -23, -64, 25, -58, -33, -64, 27, -27, -20, -35, 110, -11, 13, -41, -127, 64, 107, -39, -48, -42, -22, -31, -49, -58, 72, 27, -71, 63, 59, -103, -12, 105, 85, -62, 95, 87, 5, 7, -24, 71, -31, -37, -12, -122, 54, -13, 13, -98, -115, 71, 34, -83, -46, 68, -72, -14, -83, -39, -92, 52, 57, 41, -68, 115, -108, 61, 107, 63, -55, -69, -60, 86, -16, 120, -40, -100, -102, 98, 122, 11, 4, 17, -128, -49, -72, 112, -20, 120, -93, -77, -86, -95, -3, -126, -90, -21, -41, 24, 38, 124, -92, -44, -18, 43, 82, -103, -52, -62, -91, -50, 53, -51, -49, -99, 86, 108, 92, 32, 61, 92, 115, -3, 65, 104, -5, -52, -65, -55, 67, 59, -113, -87, -85, -35, -36, 89, 122, -66, 32, 111, 82, 97, -101, -82, 127, -101, 118, -98, -121, -33, 24, 64, 46, 38, 19, -66, -91, 27, 85, 97, -14, 56, -122, -9, -81, -117, 112, 55, -48, 77, 12, 84, 36, 33, 66, -56, 99, -29, -88, 68, -87, -99, -58, 113, 98, -52, -45, -59, 115, 5, 94, 55, 126, -110, 82, 44, -14, 70, 57, 68, -29, -26, -100, 113, 48, 75, 84, -83, -27, 35, 29, -112, -40, 42, -80, 74, 50, 45, 19, -73, 84, 97, -23, 68, 32, -52, 15, -3, -125, -9, -106, 43, -72, 25, 6, 85, 12, 45, -90, 82, -21, 126, 86, -20, 50, -53, 66, 119, -10, 84, -85, -127, -46, -128, 90, 43, 117, -58, -97, -72, 46, -65, -14, -31, -27, -84, 48, 9, 21, -47, -28, 116, -96, -74, -70, 45, 115, 52, -75, 90, 85, -23, 26, -75, 44, -41, -8, -116, -38, -106, -41, 41, -88, -117, -127, 112, -22, -122, 18, 69, -103, 85, -108, 9, 54, -125, 24, -45, -14, -27, -78, -12, 96, -81, 112, -16, 113, -54, 101, -6, 53, -14, 74, -70, 22, -31, 23, 67, 118, -11, 87, 66, 125, -33, -68, -9, 87, 99, 24, 13, -106, -26, 11, -94, 91, -103, 40, 16, 101, 17, -70, -92, -77, 93, 1, 115, -110, 13, 92, -59, -65, -2, 100, 50, 110, -62, -68, 81, -58, 45, -104, -21, 0, -125, 47, -83, -95, 59, 91, 20, 40, 38, -14, 2, 82, -96, -94, 59, -65, -128, 52, 73, 17, -126, 67, -4, -16, 98, 60, -104, -39, 10, -59, 27, -106, -56, -62, 81, 73, -9, -59, -40, -4, 27, 117, -80, 21, -55, 111, 121, -15, -16, -95, 70, -18, -82, 45, 114, 25, -119, 8, 126, 23, 38, 68, 31, 109, 91, 95, -31, 76, 64, -87, 27, 23, 0, -91, 47, 28, -16, 123, -42, -1, -124, -75, -97, 98, -97, -45, 16, -23, 25, -111, 75, -34, -55, 55, 70, 37, -39, -37, 94, 63, 5, -55, 29, -87, -15, -40, 105, -60, 27, 33, -109, 6, 11, -113, -109, 124, -45, -19, -24, -123, -45, -118, -48, -115, -96, -77, 92, 52, 122, -67, 59, -49, 113, -19, -68, -109, 61, 3, -76, 38, 39, -63, -57, 76, 106, -91, -24, -102, -95, -39, -72, -105, -16, -88, -59, -102, 125, -118, -114, -97, -94, 61, -33, -5, 114, -128, -6, -109, -60, 48, -61, 21, 46, -11, -80, 6, 106, -1, 41, 117, -15, 89, -6, -72, -106, 47, -36, -61, -35, 40, 124, 98, 107, 125, -88, 103, -35, 41, 50, -22, 50, 48, -103, -119, 99, 16, -43, 50, 81, 64, -72, -128, 41, -87, -68, -50, 50, 43, 12, -3, -21, -91, -111, -10, 59, 107, -71, -84, 3, -75, -12, -122, 123, 52, -11, -19, 69, -24, -49, -70, 81, -92, -84, 106, 95, -89, -3, -57, 99, 12, -72, -82, 48, 70, -119, 122, -62, 113, -66, -22, -125, -97, 64, -33, 20, -114, 74, -11, -81, 93, 73, 78, -96, 27, -56, -68, 28, 3, 19, -61, -19, 107, -61, 95, 82, -6, 80, -52, -44, 43, 111, 48, -74, -90, 11, -124, -82, 46, -106, 3, -115, -50, 110, -89, 113, -23, -21, 22, 82, -86, -115, -76, 17, -69, -99, 27, -91, 20, -21, 126, -66, 120, -22, -76, 17, -12, 12, 24, 38, 108, -10, 12, 80, -123, -55, 8, 28, 126, -115, -128, 113, 6, 114, -31, 78, -104, 110, 49, 6, -26, 32, -7, 86, 89, 19, 6, -11, 84, -66, 98, -78, 75, -19, -111, 122, -110, 98, 108, 36, -60, -9, -82, 98, 35, 98, -31, -67, 92, 23, -75, -119, -81, 19, -125, -65, -20, -110, -106, -124, 61, -98, 107, -9, 121, -45, -85, -103, -58, 5, -76, 6, -7, -72, 87, 95, -110, 127, 50, -111, 61, 44, 85, -117, -105, -90, -41, -42, 2, 48, -46, -60, -36, -18, -30, 119, 37, -3, 72, -65, -89, 119, 88, 15, -116, -13, -54, -17, 56, 82, 7, -97, -66, -29, 33, -16, -34, -69, -48, 105, 77, -10, 35, 95, -32, 118, -52, -47, -112, 58, -91, 108, -31, 16, -9, 19, -35, -17, 82, 49, -15, 92, 18, 69, 50, -13, -41, -44, 78, 25, 48, 33, -85, -79, 80, -80, 91, -46, 41, 28, -59, -120, 74, -127, -91, -86, 96, 37, 49, -31, -50, 58, -66, -108, 88, -126, 111, 34, 32, -15, 93, 20, -108, 55, 28, -5, 75, -24, 112, 38, 15, -87, 65, -42, 49, 64, -87, -102, 12, -83, -83, 102, 100, 96, -8, 2, -38, -110, -32, 67, 48, -62, 29, 8, 58, -4, -32, 34, 35, 83, 22, -38, 124, -85, 16, -118, -13, -103, -13, -38, 50, -89, -35, -94, -50, -110, 127, 108, 95, -38, 126, 0, -86, -85, 25, -111, 113, -84, -119, -2, -44, -126, 23, 61, -69, -50, -80, 17, 91, -30, 115, -8, -15, 52, 5, -81, 40, 92, 33, -98, -64, 6, -69, -86, 30, -41, -119, -37, -35, 9, 29, -3, -96, -42, 51, -90, 56, 34, 117, 120, -15, -78, -119, -91, 124, 50, -80, -84, 30, -8, -11, 127, -120, 108, -23, -121, -6, -51, -28, -2, 2, -35, 57, 68, -91, -59, 27, 101, 122, -105, -96, 45, -125, 101, -33, -53, -116, 10, 91, -44, 89, -15, 31, -27, -83, -28, -7, -122, -51, 11, -17, -45, 78, -110, -11, -32, 21, -51, -15, -25, 95, -23, -28, -35, 107, -80, 108, -85, -54, 84, -58, -57, -33, 126, -39, 16, -16, -25, 109, -29, -43, 33, 2, -37, -114, -72, -96, -39, 47, -21, 106, -1, -82, -90, 94, -24, 62, -68, 50, 110, 1, 119, -10, 111, -120, -51, 68, 81, 118, -28, 69, -62, -54, -75, 7, 14, -32, 103, -43, -5, -127, -71, -85, -91, -36, 37, 14, -92, 93, 85, -108, 26, -19, 32, -52, -94, 113, -67, -42, -25, -122, 81, -59, -93, -22, 88, -80, -107, -87, 98, -92, 111, -107, -117, -72, 83, -111, 84, 112, -118, 19, 101, 121, -5, 104, 93, -67, 69, -91, -5, 70, -79, 91, 110, 39, 65, -8, 70, -41, 60, -35, -31, 23, -125, -111, -43, -66, 49, -86, -109, 117, 73, -99, 7, 13, 88, -8, -104, 112, -94, 18, -88, -25, -65, 41, -11, 89, 24, 58, -109, -2, -72, -4, 61, 126, -79, -98, -72, 90, -92, 125, -86, -74, 94, -25, -87, 11, 19, 87, 13, -85, 7, 29, 64, 120, -34, 45, -92, 18, -117, -78, -32, -34, -76, -41, -71, 56, -80, 71, -97, -46, -35, -9, -74, 31, -36, -6, 8, -74, -93, -94, 53, -5, -16, 50, 48, 30, -86, 42, 91, -120, -31, 24, 22, -121, -16, -112, 97, 88, 62, 79, -93, -125, -58, -70, 113, -77, 30, -66, 57, -25, 121, -111, 54, 34, 49, -105, 74, 119, -107, -51, -54, 48, 89, -109, -14, -100, 72, 87, -97, -84, 100, 66, -62, 52, -128, 69, -27, 46, 4, -60, -101, 57, -117, -112, -61, 125, 110, 70, 86, 122, -125, -21, -34, 31, 4, -44, 64, 100, 17, -88, 14, 53, -32, 115, 101, 40, -32, 33, -81, -105, -71, -77, -117, -8, -92, 96, 43, -127, -26, 44, -109, 28, 12, 105, -82, -82, 30, -39, -4, -90, -83, -34, 124, -21, 47, -16, -30, -92, -86, 116, 4, -64, 17, -71, -38, -105, 42, -111, -111, 35, -56, -92, 9, 33, 120, 39, -78, 124, -83, 41, 2, 79, 122, -30, 6, 22, 32, -49, 56, -71, 127, -128, -102, -51, -120, -98, 121, -116, 111, -99, -36, 17, -110, -83, -3, 38, -117, -1, 75, 33, -75, -82, -119, -116, -13, -118, 32, 61, 92, 61, 88, 19, -125, 91, -13, -104, -23, 41, -125, -100, -59, 67, -1, -58, 77, -87, -102, 17, 126, 107, -76, 106, 104, -58, -70, 27, -86, 52, 44, -32, -104, -125, -78, 113, 70, 5, 51, 94, -90, 18, 113, 100, -23, 86, 122, 123, 33, -128, 96, -12, -56, -31, -4, -30, -124, 76, 29, 83, 32, -66, -122, 4, -60, 39, -127, -128, -75, -75, 41, -22, -22, 31, -109, -127, 66, -28, -14, -27, -107, -8, -109, 10, -89, 72, -43, -99, -9, 127, 122, -42, 88, -115, 76, -7, -88, -61, -102, 67, 78, 110, 67, 1, 106, 74, -35, 37, -101, 81, 38, 110, 33, 4, -113, 40, -21, -120, -104, 112, 104, 125, 48, 9, -16, -47, 56, -55, -111, -49, -97, 6, 11, -69, -115, 8, 104, 52, -18, -54, 35, 32, -64, 17, -23, 65, -49, -8, -34, -28, -101, 78, -119, -55, 50, 8, 16, -112, -118, -43, -115, -80, 117, 72, -99, 1, -93, 118, 115, 94, 83, -54, -54, -35, 100, -19, -45, -50, -74, 36, 123, 25, 75, 120, -51, -48, 42, -106, 71, 77, -103, -26, 6, -6, 92, -21, -61, -39, -128, 20, -107, 109, -112, -125, -91, -43, -74, -42, 53, 116, 13, -101, 120, -39, 75, 6, -8, -81, -128, -27, -126, 103, -127, 87, -100, -72, -59, 73, 103, -102, 69, 120, -128, -85, -94, -64, 6, -5, -93, 90, 33, 124, 119, 125, 70, 76, 49, 68, 107, -125, 53, -40, -93, 102, 64, -43, 88, -42, -6, 84, -83, -26, 102, -108, -118, 9, -13, 49, -75, 93, 75, -117, 33, 86, -7, -40, 28, 89, -97, -44, 15, 43, -61, -116, -80, 87, 47, 17, -106, -117, -125, -68, 62, 90, 34, 31, -62, 117, 72, -22, 113, -124, -47, -7, -115, -118, 102, 68, -75, -17, 72, -82, 5, 67, 80, -68, 114, -124, -1, 16, 65, 5, -49, 98, -110, 63, -103, -87, 64, 112, -68, -102, -126, 99, -73, 6, 67, -21, 14, 110, -101, 102, 20, 35, -122, 80, -44, 84, -102, 102, -116, -25, -106, 117, 122, -76, 43, -12, -9, -119, -27, 45, 111, 118, -117, -72, 125, 97, -66, 124, 2, 73, 13, 42, 116, -47, -114, -67, 44, 24, -77, -7, 108, -30, -32, -77, 68, -97, -128, 110, 44, 70, 126, -91, 113, 112, -25, -71, 79, -82, -70, 86, -16, 89, -27, -50, -25, -34, 28, -85, -23, 76, -69, -101, -17, -14, -12, 82, -12, 127, -89, 45, 104, -93, -118, -114, -14, 62, 52, 34, -105, -45, -54, 82, 95, -41, -97, -81, -119, 32, 97, 126, -7, -48, -114, -74, 127, -114, -92, 99, -40, 34, 117, 81, 2, -76, 45, -19, 87, 26, -54, -54, -48, -47, 86, -70, -99, -48, 49, -113, 23, 68, -34, -40, 70, -83, 28, 92, 100, -53, 116, -41, -59, 77, 52, 11, 29, -25, -122, 15, -95, 13, -21, 11, -117, 0, -53, 52, -42, 47, -27, -91, -96, -96, 30, 27, -112, 14, -117, -6, -122, 77, -108, -42, -23, 114, 1, -99, 93, -68, 26, 28, 30, 30, -62, 0, 51, 99, 111, -124, 65, -57, 51, 91, -3, 48, 74, -7, -64, -51, -68, -101, 9, 92, 16, 53, 118, -78, -54, 77, 86, -71, -37, 7, 35, -29, -43, 86, -121, 103, 60, -116, 31, 81, -9, -59, 67, -40, 104, -71, 123, 14, -34, -123, -46, -75, -18, 118, 69, -102, -37, 35, 122, -48, 70, -29, -120, -24, -86, -55, -102, -100, -37, 26, -24, 13, -50, -88, -97, 12, -98, 124, 118, 86, -6, 119, 125, -79, -12, 8, 0, 126, -79, 49, 85, 93, 48, 14, -49, 21, 106, -9, -60, -113, 80, 72, -36, -91, -7, 67, -17, -80, -95, -64, -7, -126, 45, 76, -31, -71, -17, 72, -113, -104, -22, 2, 60, -45, -44, -46, 3, 63, -6, 70, -78, -68, -71, 9, -61, 77, -55, -82, 42, -31, 46, 75, 84, -57, -45, -31, -51, -5, 27, -42, 104, 52, 68, -94, 22, -75, 93, -122, 67, 100, 73, 94, -104, -39, 28, -15, -33, 40, -101, 17, 58, -7, 27, 7, -43, -87, 72, -56, -26, -71, -29, 29, 115, 77, -39, -63, 112, 37, 53, -97, 77, 2, 50, -82, -116, 30, 43, -11, -59, -51, -33, 12, 31, 113, 32, 107, 96, 3, -83, -73, 43, -81, -107, -13, -121, -96, 31, -23, 88, 0, -59, 83, 78, -55, 32, 28, -72, 127, 31, 1, 102, -54, -13, 95, -121, -6, 14, 38, 98, 65, 52, 44, 123, -91, 55, -81, -92, -103, -100, -79, 94, 5, 35, -15, 118, -125, -2, 105, -102, 7, -65, 102, -4, -47, 66, 34, -29, -35, 116, -46, -119, -38, 51, -79, 3, -8, -23, -107, -38, -32, -82, -43, -59, 42, 28, 91, 43, 61, -85, -61, 8, 8, -23, 69, 51, -89, 54, 8, -50, 54, -104, 13, -46, 55, -10, 51, -47, -120, -98, 2, 108, -76, -97, 105, 72, -122, -94, -64, -29, -55, -117, 55, -86, -62, -85, 97, 6, 93, 113, -62, 111, -23, 41, -45, 38, -12, 61, 15, 105, -4, 121, -81, 27, 4, 73, 97, -49, 34, 52, -68, -28, 26, -96, -36, -37, 11, 9, 105, 120, 27, 56, 62, 40, -15, 74, -24, -8, 28, 57, -28, -53, -10, -103, -34, -115, 26, -63, 123, 15, -11, 75, 97, 77, 51, -30, -88, 87, 92, -8, 96, 101, 121, -106, -80, -111, 83, -34, 64, 70, 33, -31, -4, 39, 115, -57, 111, 121, 64, -106, 24, 51, 19, -109, 25, -125, 98, -94, -54, 7, -108, -55, 114, -19, -103, -54, 19, 20, 93, -24, -24, -58, -15, 32, -52, -13, 110, 119, 12, -66, 88, 3, -16, 83, 106, -5, 14, -20, -56, -6, -64, -17, 74, -2, -18, -63, 109, -14, 126, 27, 80, -22, -105, -126, -117, -76, -79, 0, -36, 110, -30, -96, 77, -105, 1, -7, -3, 27, 127, 102, -110, 27, -19, 55, -6, 74, 5, -90, 30, -20, 19, 111, 44, -106, -111, 66, 99, 32, -112, -17, 100, -17, 117, -54, 41, 40, -1, 108, 112, 0, 35, 7, -124, 67, 62, -95, 60, 36, -33, 86, -115, 44, 76, -60, 34, -76, -9, -90, 0, 59, 78, -28, -44, -48, 12, -61, 100, -95, -41, 51, 82, 118, -109, -127, -72, 25, 123, 25, -79, 61, 101, -76, -111, 59, -56, 125, -94, -20, -2, -119, 125, -22, 16, -51, -21, 110, 98, -35, 106, -121, -70, 79, 57, -29, 13, -116, 22, -39, 14, 77, 34, 30, 80, -31, 61, 36, 70, -59, 15, -64, 62, -46, 43, -120, -104, -120, 9, 124, -13, 63, 84, 116, -52, 7, 11, -75, -77, 93, 83, 62, -120, 82, -30, 72, 29, 72, -23, 33, -11, 115, -40, 55, 6, -35, -42, -87, 111, -22, 32, 118, 37, 95, 93, -98, 35, -100, -16, 53, -113, -90, -95, 98, -20, 67, 124, -45, -124, -108, 116, 68, -9, -106, -101, -59, 94, 126, 126, 16, -125, 109, 107, -124, -4, -7, 10, 61, 81, 121, -65, -64, -90, -48, -114, 19, 77, 50, 4, 73, 27, 34, -53, -9, -29, -94, -105, 77, 45, 48, -21, 73, 47, 97, 111, -15, -95, -114, -68, -127, 117, 70, 119, 31, -84, -62, 60, 30, 86, 55, 61, 66, -111, 74, -120, -103, 89, 107, 45, -32, 86, 53, -61, 15, 102, -112, -67, -99, -118, 89, -107, 94, -80, -31, 15, 6, 97, -9, 120, -20, 59, 57, 35, 9, 44, 28, 24, 18, 14, -48, -112, -56, 75, -92, -9, 29, -92, -51, 3, 31, -115, 47, -25, -91, -50, 121, 124, -127, 32, -72, 117, -75, 112, 42, 33, 108, -96, -25, -19, -46, 13, 43, 56, 27, -79, 9, -18, 26, -82, -62, 38, -22, 63, -119, -72, -124, -87, -25, -67, -127, 117, -33, 39, 56, -73, 118, -88, 98, 15, -12, -3, -57, -11, 32, -72, -15, -86, -104, 117, 121, -103, -90, -51, 67, -72, 86, -85, -91, -62, -101, -60, 6, -44, 102, 18, -21, -84, -19, 64, -75, -69, 39, -26, -27, 43, -75, 53, -39, 22, -6, 56, 46, -44, 6, -106, 114, 18, -125, 110, -122, 105, 105, -109, -76, -12, -36, 84, 39, -98, -40, -32, -56, -104, -40, -70, -91, 9, 92, -50, 6, -113, -4, -29, 18, -45, 39, -94, -46, 20, 108, 52, 52, -122, -97, 80, 20, -4, -45, 10, 48, 14, -69, -70, -59, 71, 2, -60, -109, -7, -85, -52, 4, 116, -7, -19, -2, 63, 48, -26, 26, -29, -121, 19, -11, -65, -75, 74, 35, 51, -85, 94, -46, -123, -21, -12, 65, 61, 124, 123, 29, 25, 1, -15, -113, -92, 10, -36, -3, 124, -68, -34, 30, 124, 65, -108, 44, 124, -48, -77, -54, -37, -121, -27, 53, -30, -127, -40, 127, 72, -125, -106, -56, -91, 101, 113, 21, -50, -118, 38, 51, -92, -46, 5, 16, -59, 53, 124, -88, -103, -125, 55, -69, -50, 9, 84, -16, -89, 94, -83, 54, 112, 42, 65, -35, 0, 6, -99, -103, 44, -43, -2, -60, 100, 42, 114, -2, 104, -95, 87, 101, 25, 101, 19, -58, -5, 20, -47, -125, 34, 5, -67, -103, 55, -15, 34, 50, -77, -89, -73, -88, -72, -104, -16, -75, 15, -37, -41, 26, 26, 28, 5, 19, -96, 123, 51, -5, -95, 104, -40, 74, 31, 119, -97, -77, 11, 87, -26, -35, -90, -65, 7, 64, 45, -51, -116, -47, -18, 122, -11, -62, -73, -51, -54, 43, 42, 72, 80, 107, 24, 112, 42, 121, 100, 39, -34, -71, 11, -17, 108, 8, 70, 15, -123, 15, -37, 88, 108, -76, -128, -42, 67, -58, 41, 61, -116, 14, -95, 106, -16, -45, -103, -57, 125, 75, -79, 65, 17, 7, -9, -51, 47, -124, 95, -120, -50, -88, -29, 40, 117, 108, -70, 5, -75, -44, -73, 50, 41, -72, -94, 2, -116, -79, -102, -22, 90, -101, 33, -51, -52, 34, 14, -32, -1, 19, -126, -56, -91, 71, -66, -57, 10, -127, -38, -89, -94, -8, 40, -76, 20, -87, -25, 123, -13, 72, 69, 56, -13, -127, 88, 41, -24, -100, -55, -29, 79, -71, 106, -71, -43, 70, 58, -89, 61, -32, -77, 20, 10, -41, -63, -47, 40, -5, 122, -76, -75, 3, 111, 118, 103, 60, -57, -95, 114, -46, -88, 51, -53, 25, 38, 126, -58, -57, -89, 20, -116, 85, -61, -46, 16, 109, -53, -22, -43, -62, -23, -14, -32, -101, 23, -124, 4, -84, 123, -101, -35, 110, -110, 66, -106, 123, 61, 26, -118, -61, -95, -87, -32, 53, -28, 53, 83, 31, 117, 20, -59, -46, -77, -43, 94, 0, -20, 76, -14, 32, -18, -55, 12, 123, 120, -57, -21, 93, 112, -14, 62, -44, -30, 126, 49, 76, 90, -7, -82, 92, -49, 46, 30, 47, 74, 18, -114, -38, 87, -95, -120, -102, 9, 5, 73, 102, 18, -97, 125, 50, -44, -33, 55, 90, 87, -124, 62, 82, 53, -69, 54, 8, 1, -123, -117, 62, 1, 93, 37, -33, -38, 59, -88, 54, 72, -128, -89, 60, 41, 102, 108, -29, -102, -35, -47, 78, 54, -67, 31, 78, 111, 59, 44, -71, 118, -72, 104, -93, -75, -60, -25, 84, 103, 23, 3, 61, -85, -23, 55, -59, 47, 69, -35, 14, -23, 79, -123, 104, 61, -69, 69, -77, -4, -30, -67, -107, 112, 5, 88, 98, -103, 60, 64, -115, -87, -67, 109, -116, 76, -7, 107, 123, 69, -31, -91, 17, 3, 69, 33, -80, 5, 0, 98, 35, 18, 15, 60, -128, -112, 127, -43, -26, -85, 68, 32, 62, -38, -118, 83, 112, -90, 5, -36, -51, -123, -1, 43, -126, 16, 103, 40, 40, -50, -91, 34, -38, -48, -29, 33, 32, 9, 91, 125, -14, 19, -37, 67, -41, -54, -124, -72, -39, -114, 92, -23, 22, 105, -105, 17, 44, -27, 80, -98, 109, -100, -106, -57, 89, 110, 5, -17, -19, -100, 90, -6, -111, 82, -44, -43, 18, 48, 31, 117, -47, 57, 18, -81, 107, -48, 56, -72, -23, -14, -128, 56, 11, 78, 99, -88, 92, 62, -92, -24, 16, -36, -34, 60, 8, -83, 93, -118, 124, 58, 16, -121, 35, -103, -84, 16, 53, -103, -116, 50, 21, -66, -28, -116, 104, -4, 14, 15, 95, 106, -89, 21, 45, 84, 76, 45, -87, 108, -109, -18, -18, 119, 111, -110, -8, 94, -121, -89, 55, -107, -53, -4, -97, -65, 88, 87, 8, -110, -44, -32, 81, -112, -125, -47, 109, 52, 75, 6, -122, 118, -123, 79, 90, 39, 20, 119, -117, -65, 88, 27, 124, -11, -126, 87, -89, -36, 123, 17, -65, -46, 72, 34, -56, 117, -128, -85, -30, -3, 6, 124, 28, -86, 27, 90, -95, 127, 109, 16, -92, -112, 68, 90, 13, 34, 78, 26, 104, -17, 25, -33, -59, 118, -72, -123, 37, 71, 115, 33, -2, 0, 20, -127, 2, -91, 107, -61, 21, -15, -92, -55, -18, -39, -3, 59, 70, -116, -119, 64, 81, -91, 16, -9, -31, 105, 124, 45, 76, 44, 58, 8, 62, 112, 87, 32, -7, 44, -112, -90, -42, 69, 112, 32, 112, -49, 91, 88, 126, -80, 18, -124, 45, 121, 46, 89, 94, -18, 55, -79, -33, 109, 99, -66, 39, -67, -69, 87, -43, 113, -105, -10, -16, -87, -21, -44, 52, 56, -104, 48, 69, 98, 70, 49, 48, -14, -42, -12, -81, -86, -34, 118, -50, 73, 115, -122, 19, 24, 88, 91, 3, 22, -42, 97, -20, 100, -73, -84, -38, -15, 26, 37, 15, 116, 51, -69, 36, -110, -8, 18, -14, 30, -65, 66, -93, 85, -107, -8, 58, 91, -92, 122, 52, -24, -60, 127, -9, 23, 43, -73, 99, -26, 122, 116, -93, 119, -112, -71, 16, 2, 20, 107, 34, -64, 108, 42, -18, -7, 33, 35, -96, -61, -107, 105, -96, -54, 58, -46, 113, -110, 82, 43, 90, 74, -47, 78, -91, 86, -124, 92, 88, -94, -16, 122, -74, 71, -100, 121, -109, 118, 112, -58, 93, -97, 84, 96, 90, 0, 20, -104, 113, -77, -111, 25, -49, -105, 9, 37, 103, -88, 32, -82, 20, 87, 116, -18, -60, -65, -21, -15, -88, -22, 40, -4, -10, 1, -123, -23, 88, 31, -118, -65, -94, -95, 29, -110, 23, -35, -43, 24, -40, -91, 7, 7, 93, -42, -26, -102, 4, -5, 37, 35, -17, -62, -118, 80, -45, -79, -60, 10, 20, 32, -41, -35, -10, 17, 0, 6, 109, 120, 57, -74, 67, 95, -68, 97, -5, -48, 101, 108, 94, 37, 19, 30, 5, -53, 21, -101, -105, -2, -43, -64, 103, -21, -37, 41, -124, -46, 94, 88, -121, -106, -40, 6, -22, 3, -102, 94, -113, 68, 46, -67, 127, 74, -54, -80, -73, -108, -128, -76, -19, 73, -104, 11, -19, -18, 125, -42, 80, -45, 97, -123, 91, -23, 80, -51, 73, -124, 1, -86, -73, 56, 74, -55, 100, 69, 75, -116, 19, 51, -122, -123, 15, 91, 11, 1, -4, 73, 127, 35, -104, -12, -14, 51, 115, 70, -66, 83, -52, 120, 98, 78, 34, -5, -54, -36, 23, 37, 99, -2, 25, 65, -19, -39, 64, 109, 90, -43, -38, -20, -127, -10, -19, 4, 118, 63, -46, 36, -18, 95, -24, 40, 111, 8, 127, -43, 37, -49, -61, 120, 4, -7, -28, -61, -109, -24, -17, -93, -21, -64, -33, -80, -60, 9, 59, -107, -7, 125, 90, 32, -88, -110, -72, 46, -104, 78, -58, 44, -61, 84, 51, -102, 10, -68, -43, -94, -6, -17, -81, 109, 67, -38, 12, -105, -45, 9, 3, -29, -23, -44, 26, -81, 35, -103, 25, 119, -37, 114, -112, 86, 78, 63, -80, -39, 8, 33, 124, -128, 32, 23, 46, -75, 65, -68, -31, 31, -38, 69, 93, -112, 3, 85, 126, -67, -126, -82, -84, -41, 109, 62, -34, 79, 6, -84, -32, -40, -6, 31, -123, 8, -85, -64, -24, -19, -3, -124, -55, 31, -123, -57, -35, -51, -102, 57, 33, 73, 31, 46, -105, 98, -59, -52, -87, 81, 119, -102, 47, -41, 36, 70, 12, 44, 93, -105, 44, 105, 80, 59, -121, -24, -70, 79, -15, 35, -46, -2, -77, -79, -7, -68, -30, 12, 83, -29, -80, 64, -126, 17, -85, -75, 113, 119, 120, 100, -65, -54, -119, -104, -51, 123, 105, -68, -56, 98, -120, -46, -36, -8, 65, -30, 88, -30, -58, -90, 26, 34, -32, -110, 89, 49, -32, -125, 72, 93, 97, -64, 10, -77, 35, -8, 8, -124, -46, 31, 78, -63, 67, -122, 113, -117, -12, -10, 126, 31, 113, -33, 72, 59, -37, 127, 74, -121, -42, 54, 59, 52, 123, 81, -125, 119, -98, 87, 36, 8, -43, 14, 67, -127, -60, 98, -59, 78, -98, -64, -80, -3, -69, 19, -61, -121, -58, -7, -51, -20, 53, 87, -36, 58, -11, 10, -29, 10, -117, -94, -105, 7, 41, -8, -4, 38, 22, -121, 80, 60, -125, 109, 85, -3, -104, -30, 100, 35, -93, -36, -105, -114, -92, 104, 49, -69, 109, -76, 73, 4, -40, -19, -86, 69, 36, 92, -25, 0, 17, -112, -56, -35, -59, 87, -44, -99, 62, 50, -7, 69, -15, -28, -99, -29, -99, 54, 9, 73, -44, -54, 57, 9, -112, -4, -25, -17, 32, -64, 29, 2, 83, 100, 7, -73, 95, 86, 38, 102, -89, 50, 122, -32, -22, -37, -9, 113, 17, -71, 66, -45, -121, 64, 47, -47, 29, 17, -30, 71, -98, -45, 29, -13, -66, -106, 65, -48, -10, 121, 84, 115, 67, -15, 115, -21, -10, -30, 92, 86, 65, -35, -101, -114, -117, 83, 51, -36, 115, -75, -79, -69, 0, 107, -97, -72, -44, -27, 94, -87, 125, 93, -76, 43, -118, 117, 43, 66, -46, 104, 67, 111, -115, 35, 115, 125, -107, -17, 33, -94, -113, -47, 104, -113, 24, -126, -66, -124, -115, 64, 15, -31, 117, -110, 111, 70, 91, 5, -101, -111, 4, 55, -18, -62, 68, 55, 59, 82, -102, -19, -49, 31, -75, -71, 69, 82, -85, 82, -47, -8, -72, -109, -72, 119, 122, 112, 13, -60, -15, 0, -35, -114, 62, -108, 87, 63, 75, 111, 30, 48, 51, -125, -36, 87, 91, -15, 25, -102, 90, -104, -46, 48, -127, -13, 44, 116, -77, 60, -104, 81, -12, -10, -70, -98, 8, 23, -52, 51, 23, 40, 79, -106, 112, -61, -14, 100, -48, -100, 123, -78, -16, 126, -109, -26, -112, 0, 112, 88, -79, -63, -61, 49, -34, 112, 91, -26, 48, -72, 52, -80, 66, 1, 10, 52, -114, 91, 51, 80, -88, 102, -125, -98, 31, 59, -41, -127, -24, 6, -115, 98, -93, 20, -24, 120, -108, -112, -95, -86, 19, 57, -73, -123, 26, -39, -2, -81, 59, 72, -84, 14, 54, 20, 115, -97, -49, 114, 110, -72, -79, 74, -27, -109, -101, 24, 126, 15, -88, 97, 42, 68, 40, -42, 124, -47, -12, -46, 58, -50, 82, -43, 97, -47, -49, -57, -71, -7, 47, -74, 17, 4, -86, -8, 56, -90, 19, 9, -14, -54, 88, 57, -61, -59, 51, 19, -73, 106, 8, 76, 70, 63, -107, 99, 48, 73, -36, 23, 77, 28, 19, -11, 103, 54, -29, 12, -64, -97, -22, 115, 28, -73, 62, -36, 54, -41, -122, 31, -9, 62, 32, -13, -29, -28, -41, 36, 32, -53, 103, -42, 32, 34, -110, -125, 90, -72, -123, 93, -55, -59, 125, 0, 108, -93, -88, -101, 88, -127, -38, -2, 37, -94, 33, 43, -101, -124, -27, -16, -93, 8, 90, 39, 83, -126, -98, 24, -56, -90, 104, -73, 108, -28, 111, 118, -92, 4, 95, 52, -43, 110, 107, -96, 18, -56, -128, -62, -41, -23, 44, 101, 38, -81, 56, 45, -110, -29, -47, 91, 43, -27, -18, -19, -123, 28, -62, -97, 98, -23, -104, 20, -78, -48, 12, 17, 117, 41, 89, -119, -110, 79, 97, -122, -124, -97, 65, 57, -7, -39, -91, -55, 46, -124, 75, 73, -113, 104, -12, 121, -63, 66, -30, -89, -51, -3, -75, -39, -37, 96, 80, 69, 14, 41, -79, 38, -108, 98, -67, 9, -69, 59, 9, -83, 77, -75, 12, 91, 23, 20, -11, 91, -121, -20, -34, -12, 82, -89, -122, -62, -16, -34, -112, -35, 76, -91, 6, 98, 66, -19, 45, 127, -105, -28, 125, 34, -47, -55, -116, 49, -68, -96, -14, 33, 127, 18, -27, -118, -73, -74, -54, 83, -73, -67, -58, -110, -71, 32, 84, -23, 5, 120, 49, -21, 34, 95, -67, -30, 123, -115, 14, -27, -15, -20, -90, 106, 65, -96, 52, 13, 96, -11, -20, -115, 110, -43, -14, -119, -19, 53, 109, -30, 21, -24, 36, -102, -38, 76, 13, -42, -100, 49, 58, -85, -27, 118, -19, 79, -65, 88, -4, 99, -108, -29, 29, -89, -30, -53, -81, 99, 120, 40, -82, 92, -104, 49, -8, 23, -33, -118, 96, 91, 124, 28, -20, 51, 77, -82, -94, -81, -39, 55, -61, 42, 0, -54, -80, 35, 9, 120, 33, 48, 35, 77, 99, -59, 10, -27, 45, -29, 113, 35, -50, 28, 80, -72, 53, 79, 2, 111, 111, -77, -23, -50, -74, -15, -26, 116, 7, -68, 54, 116, 1, 8, -66, 25, 28, -116, -116, 25, -76, 5, 109, 86, -13, -4, -76, 36, -41, 83, -119, -56, 109, -26, 55, 124, 26, -91, 115, -52, -101, -11, -10, -46, -102, 20, 42, 63, 74, 61, -47, -48, 103, -21, -91, 52, 16, -30, -115, 58, 52, 115, -52, -26, 29, 14, 107, -91, 74, -96, -50, 90, 109, -96, -42, 21, 73, 117, 104, 110, -93, 88, 32, 21, 43, -57, -33, -66, -112, 121, 30, 58, -68, 60, 2, 27, -89, -113, 77, -20, 105, -85, 2, 1, -25, 22, 76, 73, -105, -65, -102, 8, 126, 88, 103, 6, 54, -121, -64, -92, -41, 123, -3, 17, -38, 126, 39, 56, 101, -55, -16, 80, 95, -5, 63, -81, 47, -32, -119, 5, -99, -109, -34, -123, -110, -72, 40, 43, -126, 40, -41, -119, 42, 48, 39, 94, 84, 27, -104, 8, -32, 77, 100, -87, 119, -101, 104, -45, -38, 86, 0, -40, 109, 78, 20, -20, -127, -115, 43, 2, 57, 60, -32, 87, -47, 22, -12, 44, -117, -9, 124, 92, -86, -37, -48, -65, 52, 83, 81, 37, -36, -17, -83, -54, 28, 102, 111, 126, -14, 88, 125, -108, 36, -64, -35, -53, 72, -29, -101, -17, 20, 76, 54, 24, 19, -54, -95, 60, -63, -24, -69, 20, 63, 123, 100, -98, 84, -18, 51, 61, 111, 119, -108, 49, 45, 64, 100, 107, 22, -41, -116, -4, 21, -110, -110, -37, 80, 2, -15, -33, -73, -20, 110, 105, 14, 36, -47, -43, 81, 102, -116, 63, -95, -43, -88, -62, 21, -98, 35, 123, 60, -94, 116, 22, -127, 63, -112, -34, 113, 30, -7, 47, 31, 6, 57, -5, -121, -61, -23, -55, -99, -77, -43, -70, -23, 83, -12, -109, 118, -97, -52, 106, -35, 10, -25, -17, 46, -75, -32, 55, -117, 110, -107, 54, 53, -4, -123, 79, 122, -114, 13, 99, 19, 66, -119, 67, -84, -117, -43, 75, 67, 55, -60, -74, 100, 124, 118, -57, -55, 3, 64, -110, 107, 107, 41, -45, 43, -27, -50, 97, 89, -10, -25, -87, -118, -4, -24, -24, -57, -15, -72, 33, -38, -56, 96, 11, 77, -91, -51, 64, -20, 126, 58, 89, -91, -118, -97, -30, -9, -46, -63, 72, 21, -83, 123, -104, 45, -121, 105, -127, 119, -127, 41, -64, 44, 22, 11, 116, -14, -47, 42, 117, 83, -128, 121, 78, 112, 127, 123, 47, 6, -69, 52, 65, -67, 0, -16, -8, 70, -12, -12, -18, 80, -51, -50, -102, 107, 122, -118, -7, 69, 89, 43, -108, 29, -16, -117, 15, -88, -89, -60, -11, 114, -93, -38, 84, 36, 3, 11, 25, 16, 94, -23, -29, 94, 9, 35, 100, -1, -56, 110, 104, -56, 4, -26, 81, -28, 111, 122, 15, 18, 43, 60, -31, 28, -64, 30, -112, -127, 20, -31, -21, 8, 106, -39, -124, -26, -99, -43, 26, 4, -128, -32, -43, 96, -98, -19, 73, -23, -81, -59, -112, -107, -17, 55, -25, 43, -19, -82, -75, -46, -51, 109, 58, -98, 113, 47, 116, 15, -5, 0, -119, 75, 112, 127, -109, -69, 115, 58, 65, 55, 12, 53, 103, -60, -25, -15, 12, -122, -33, 56, -51, 5, -74, -112, 95, 14, 46, -122, -94, -125, 122, 39, 51, 114, 70, -110, 127, 1, 53, 47, 28, 61, 23, 125, 108, 62, 96, -88, -90, 32, 21, -95, -122, -108, 64, -32, 34, -62, -1, 75, 53, -115, 51, 7, 92, 42, 69, 32, -120, 83, 97, -68, 66, 125, -127, -39, -75, 12, 111, 50, -10, 30, -3, 70, -20, 123, 34, 34, -45, 19, 65, 34, -45, 66, -78, 114, 58, -86, -119, 116, 0, 46, -78, -5, 28, 65, -40, -61, -19, -57, -114, -115, -124, -41, -41, -77, 124, 105, 109, -90, -101, -78, 2, -97, 39, 51, 66, 94, 61, 74, -99, 65, 98, 26, -124, -4, -80, -41, -97, -121, -12, 72, 92, 58, -104, -70, 1, 19, 98, -127, -14, 10, 50, 20, 64, 49, -20, -83, 12, -1, 110, 3, 68, 23, 72, 6, -19, -38, 35, -117, -46, 95, 106, 121, -33, 98, -79, 64, 25, -51, -128, 78, 70, -39, 86, 25, 68, -71, -97, 50, -84, -15, 29, 83, -70, 104, -22, 120, 39, 63, -60, -113, -84, -102, 77, 70, -76, -104, -22, 60, -104, -12, 108, -37, 65, 57, 105, 116, 103, -99, 14, 19, 3, 118, -31, 122, 97, -1, -66, 41, -128, 65, 124, -82, 9, 54, -100, -102, -95, 33, -118, -9, 49, -103, 30, 84, 52, 45, 121, 116, -58, 52, 81, -75, -107, 30, 29, 5, 71, -28, -91, 103, 126, 106, -67, 114, -58, -124, -27, -28, 86, -34, 63, 107, 4, 31, 9, -11, -34, 100, -7, -114, -65, -28, -68, 112, -12, -122, -79, -61, -84, -4, 86, -127, -56, -103, -90, 96, -113, 33, -58, -70, 67, -9, -1, 77, 17, -32, 48, -119, 71, -24, 93, -80, 10, 100, 41, 104, -88, -116, 55, 15, -104, 44, 90, -23, 97, 88, 68, -86, -119, 41, 91, 38, -3, -123, 58, -56, -47, -91, 63, 85, 99, -61, -20, -50, -48, -33, -30, 23, -80, 20, 53, 49, -109, 83, 24, -26, 107, -72, 62, 55, -41, 49, 106, 6, -2, 60, -33, 45, -31, -91, 110, 75, -80, -94, -15, -46, 37, -95, 124, 55, -68, 19, -107, 106, -108, -127, 4, 27, -23, 100, 92, 76, -115, -14, -14, 4, -33, -127, 29, -99, -66, -115, 124, 81, -110, -127, 13, -79, -115, -92, -54, -36, 38, -114, 6, 119, 41, -46, 109, -127, 126, 87, 53, -41, 23, 23, -89, -7, 80, -22, -60, -101, -23, 20, -68, -33, -6, 91, 2, 83, 14, -36, 127, 127, -30, -43, 109, 118, 40, 115, -15, -1, 110, -98, 11, 110, -30, 114, 99, -41, 2, 115, 66, -57, -28, 90, -16, 73, -42, 2, -80, 14, 30, 94, -61, 118, 124, -57, -68, -1, -104, 19, 25, -7, 19, 6, 31, 17, 9, 86, -85, -105, -85, 117, -40, 64, 19, 12, -35, -79, 9, -93, -10, 37, -63, -25, -44, 16, -99, 71, 3, -124, -125, 28, 78, 119, -91, -114, 27, -9, 50, 89, -103, -84, 93, -108, 31, -42, -105, -30, -114, 5, -103, -78, -51, 122, -29, -30, 30, -126, 69, -50, 22, -35, -108, 101, 64, -94, 24, 73, -119, 111, -44, -21, 62, 49, 113, 47, 0, -22, 106, 120, -53, 44, 10, -70, 112, -18, 70, 90, 9, -11, -43, -59, 39, 19, 22, -31, -22, 48, 63, -87, -58, -34, -78, -109, -111, 67, -27, -109, -6, -26, -62, 99, -102, 5, -101, 92, 4, 65, 74, -26, 25, 10, -53, 39, -108, 113, -73, -21, -92, -40, 69, -42, -105, 111, -54, 5, 19, 98, 16, 15, 62, -41, 18, -36, -41, 111, -49, -69, 93, 19, -38, -118, 35, -18, 64, -79, -36, -57, -66, -4, -59, -117, -24, -20, -48, 119, 27, -65, -71, 125, 110, 15, -45, -47, -50, -34, -99, 27, 83, -114, -82, 79, 106, 94, 124, -8, 19, -71, 13, 83, -25, -7, -35, 101, 61, 58, -48, 70, -35, -6, 44, 7, -77, -3, 1, -91, 102, 15, 11, 99, -127, -42, -83, -7, -1, -48, -54, 34, 26, 108, -113, -54, 62, -78, -56, 107, -30, 74, -96, -92, -88, -92, -3, 26, -37, -31, 42, -44, -94, 32, 78, 106, -55, 79, 19, 50, -35, -32, 32, -71, 85, 98, -80, 96, 46, -13, 14, 99, -36, 19, 112, -63, -33, 43, -73, 80, 120, 31, -2, -30, -87, 26, -109, 121, -106, 121, -99, 106, 38, -10, -77, -4, -111, -76, 36, -63, -3, -101, 105, -54, 97, 101, -2, 117, -93, 116, 102, -27, 50, -45, -68, -16, -60, 23, -125, -85, -111, 51, 39, 69, -65, -69, -42, -124, 34, -59, 7, -25, 98, 23, 34, -124, 83, 99, 25, -115, 63, 34, -114, 124, 32, -82, 54, 6, 125, 66, -104, 121, 9, 94, -43, -23, 33, -92, 82, -98, 41, 69, -22, 40, -128, 52, -10, 0, -126, -82, -66, -24, -28, -24, -40, -21, -54, -121, 24, 3, -84, -89, -37, -65, -116, 57, -44, 57, 9, -15, -99, -75, 74, -78, 76, -59, -37, 51, 127, -57, 82, 47, 92, 4, 0, -18, -100, -33, 9, -17, 33, 31, -86, -71, -62, 34, 77, 108, 116, 27, 104, 94, 123, -54, 100, 3, 3, 54, 52, -48, 2, -81, -87, 24, 12, -49, -78, 58, -59, -24, 20, 4, -63, 104, -82, 119, -69, -20, 121, 14, 77, -29, 89, 89, 111, -106, 49, -29, 74, -25, -97, -43, 13, -48, -84, -5, -107, 126, -41, 17, 15, -23, 86, -74, 4, -73, 58, -103, -31, 112, 105, -10, -97, 26, 36, 121, -41, -61, 21, 81, -95, -41, -59, -99, 82, -43, -63, -49, 107, 26, -27, 23, -22, -27, 97, 35, -88, -22, 42, -28, 73, -111, 90, -121, -43, 115, 104, -100, -40, -99, -15, -66, 31, 115, 52, 19, -77, -3, -19, 45, -118, 34, -43, 27, -85, 49, -114, -118, -67, 122, 70, 39, 37, -41, -18, -104, 38, -54, 89, -71, 20, 39, -37, -79, -44, -65, 72, -9, 110, -17, 103, 96, 98, -47, 32, 113, -50, 79, -83, 10, -36, -83, 8, -42, -15, 14, 118, 13, -36, 90, 62, 23, -67, 92, -54, -29, -71, -47, -76, -64, 13, -66, 22, -107, 1, -7, -41, -15, -3, 42, -63, 45, -61, 125, 24, -90, -4, 45, 47, 49, -51, -88, 82, -69, 30, 31, -113, -60, 112, 62, -28, -88, 68, 38, -40, -94, -114, 102, 20, -54, -11, -116, -91, 22, 100, 89, -67, 54, -55, 60, 75, -46, -64, 125, 97, -91, -86, 95, 90, -26, 41, 115, -128, -49, -86, 110, -16, -109, -81, -51, -56, -19, -93, -41, 66, -46, 77, -100, 33, -39, 82, 0, 33, 127, 86, -1, 91, -101, -6, -122, -67, -51, -105, 110, -78, -59, 1, -17, 64, -34, 25, -116, 22, 48, -104, -84, 77, -125, -82, -91, -125, 7, 22, 28, -10, 2, 6, 48, -116, 62, 49, 96, 74, -16, 19, 93, 24, 61, 63, 49, -80, 35, 21, 81, -1, 28, 112, -94, -34, -123, 24, 74, -90, 95, -113, -19, 49, -52, -79, -102, 81, 53, 109, 86, -85, 108, -52, 71, 67, 47, 36, 56, -31, -37, -50, -24, 65, 77, 14, 16, 40, -114, 24, 2, -33, 37, -76, -10, -103, 77, -70, -21, -9, -22, -14, 53, -19, -35, 50, -94, -87, -120, -55, -43, 25, -28, -88, -79, 98, 26, -45, -92, -15, 37, -4, -127, -20, -31, -72, -47, -36, -128, 32, -95, -24, -91, 126, -46, -77, -88, 102, 88, -78, 122, 14, 11, 70, 9, 80, 36, 114, -126, 24, 64, -50, -57, -61, -14, 54, 107, -72, 30, 38, 53, -45, 21, -70, -43, 30, -46, -106, -105, 66, 17, -74, 48, -28, -76, -25, -86, 30, 10, 54, -34, -110, -72, 74, -60, 105, 8, -21, 56, -71, 120, -24, 63, -44, 6, -18, -24, 94, 19, 19, -23, -49, -60, -2, 61, 56, -69, 18, 16, -59, -43, -9, -10, 64, -12, -6, -103, 127, 67, -69, -81, -34, -117, -4, -53, -43, -62, -75, 43, -2, 45, -3, 41, -84, -9, 110, 67, -57, 111, -23, 94, 8, -94, -105, -57, 87, 82, -97, -9, -18, 21, -94, -87, 66, 26, 51, -67, -55, 22, 112, -86, 45, 119, -63, 13, -76, -23, -98, 51, -80, -2, -3, 12, -90, -59, -77, -19, -87, 18, 109, -98, 9, -74, 81, 29, -70, -28, -79, 43, 31, 53, -26, 29, -12, -90, 82, -94, 95, 70, -123, -70, 117, -47, -14, 46, -117, 106, 45, -93, -49, 1, 124, -32, 122, -84, -99, 100, -22, -79, -3, -31, -108, -51, -22, 17, 38, 71, -71, 38, 58, 60, 123, -31, -97, -83, 98, -5, -116, -3, -22, -97, 84, -12, 40, -66, 65, 44, 53, 2, 71, -84, -71, -118, 4, -42, -84, -75, -2, 120, 29, -28, -66, 120, -43, 30, 115, 81, 79, 38, 124, -33, -119, -13, -48, -82, 30, 62, -61, 20, 80, 46, 48, -32, -100, 24, 44, -29, 1, -118, 114, -75, 85, -90, -78, -119, 22, 31, 13, 11, 63, 106, -70, 92, -91, 26, 102, 126, 104, -14, -45, -40, 127, 76, 49, 6, -88, 103, 35, 82, -97, 107, 72, -30, -79, 109, -6, -7, -127, -54, -121, -88, -1, 94, -14, 81, -71, 31, 38, -99, 111, 37, 54, 30, -53, -50, 86, 126, 127, -5, -101, -18, -51, -79, 97, -60, -22, -19, -34, 35, 31, -17, 17, -26, -96, -80, -88, -44, 67, -77, -92, -57, -109, -18, -105, 108, 19, -13, -101, 9, 41, -54, -74, 27, -14, -68, 116, 51, 118, 107, -3, -119, -50, -113, 81, -46, -111, 7, 82, 119, -20, 43, 85, -98, 72, -85, -85, -94, 62, -79, -73, -70, -9, 44, 109, 58, 48, 39, 111, -96, 117, 110, 84, -112, -42, -21, -103, -6, 72, -35, 68, 39, 88, 35, -26, 81, 32, 10, 114, 42, 77, -50, -91, 100, -101, 108, 18, 8, -15, 70, -68, 12, -30, -54, 91, -76, -76, 37, -33, -68, -107, 12, -66, -115, -29, -48, -44, 30, 75, -53, 6, -97, 102, -54, -124, 81, 120, -113, 34, -22, -98, -113, 69, -99, 105, 110, 99, -124, 106, -95, -49, 57, -11, -28, 115, 50, -50, 62, 62, -86, 9, 86, -13, 77, 112, -29, 101, 12, -50, 66, -20, -50, -58, 45, -121, -116, -46, 31, 29, 123, -86, -122, -3, -1, 0, -99, -99, -66, -88, -93, -87, -95, -96, 93, 52, 21, -18, -3, -73, 118, -121, 84, 75, -47, -7, -12, 123, -58, 62, -34, -122, -52, -68, -49, -122, 31, 62, -68, 85, 40, 4, 12, 79, 117, 25, 2, 64, -42, -108, 40, -60, -120, -20, -81, -46, 118, -15, -125, 29, 122, -77, 31, -123, -15, 93, 126, -76, -72, 72, -42, -97, 89, -72, -123, -109, -107, 1, -43, -71, 29, -34, -83, 41, 96, 72, -93, -7, 124, 122, -76, -79, -121, 60, -40, -92, -103, 119, 71, 115, 42, 23, 85, -65, -43, 17, -5, 27, 44, 0, 19, 46, 110, -125, 35, -78, 42, 124, 8, -85, -50, -57, -72, -22, -96, -53, -67, -63, -41, -81, -26, 76, 76, -100, -118, -14, -121, 85, 51, -41, -26, -60, -93, -126, 102, 79, -61, -52, -35, 84, -111, -39, 77, 107, -45, 15, 115, 86, 83, -21, 42, 20, -38, 57, -52, 11, 62, -113, -61, -106, 123, 17, 54, -16, -19, -124, -97, -14, 52, 34, -11, -98, -20, 71, 108, 123, -63, 93, 123, 42, -43, 11, -42, -35, 55, -4, 41, -85, -95, -51, 40, 90, 112, -124, -96, 88, -103, -79, 1, -124, 104, 35, -50, 43, -63, 106, 66, -65, -81, 72, -50, 71, 1, -64, 0, -113, 51, -97, -60, -90, 19, 3, 65, 69, 56, 11, 33, -88, 30, -19, 115, 56, -84, 20, -22, 116, 4, 15, 71, -121, -26, -28, 43, 121, -124, 13, 69, -90, 46, 32, -80, 112, -77, 53, 57, 54, 25, 40, 49, -51, 1, -55, -8, -119, 23, -69, -26, -45, -69, -63, 13, -24, 83, 124, -115, -46, -44, 22, 79, -91, -77, -125, -113, -50, -105, -119, 88, 118, 8, 118, 16, -6, -47, -11, -49, 35, -93, 98, 111, 50, -65, 36, 29, 22, 93, 32, -7, 112, -43, 102, -95, 107, -118, 41, 102, 23, -62, -20, -42, -62, 112, 91, 123, 27, 67, 106, 69, 30, -51, -27, -34, 58, 62, 32, -68, 111, 84, 7, -125, -108, 87, 70, -18, 78, 35, -70, -74, 110, 68, 14, 32, 37, 29, -81, -59, 36, 73, 13, -59, -74, 107, 110, 76, 111, 80, -39, -104, -75, 44, 2, -21, -14, 96, 90, 63, 63, 94, -54, 14, 90, -66, 36, 73, 110, 98, 54, -11, -81, 91, 19, 30, -108, 103, -89, 17, -45, -30, 105, 53, -123, -47, 31, -16, 64, -30, -109, 12, -76, -32, -41, 36, 2, -74, 68, 75, -98, 13, 119, -60, 62, -3, -50, -117, -63, 45, 113, 33, 95, -5, -49, 31, 127, -25, -119, -125, -113, -14, 23, 83, -124, -55, -45, 36, -85, -23, 98, -78, 104, 44, 116, 58, -10, -5, 76, -83, 15, -45, -106, -74, -103, 73, 56, 47, -54, -21, 9, 6, 14, 106, -62, 14, 108, 43, -113, 75, 13, -30, 73, 120, -125, 21, 25, -80, 3, 116, 13, 89, -10, -38, 102, -76, -67, 68, -39, -69, 57, -89, -20, -106, -75, -53, 116, -38, 37, -23, 28, -100, -83, 98, -98, -74, -43, -74, 23, -26, 67, 39, 40, 101, -44, -10, 11, -11, 62, 35, 49, 99, -87, -112, -9, 30, -13, -121, -56, -72, 25, -32, -32, -83, -103, -127, 85, -105, -3, 47, -75, 58, -119, 123, 64, -14, -22, 48, 123, 120, -66, -24, 96, -16, -26, -98, -111, -6, 3, -28, 81, -58, 64, -98, 32, 123, -50, -98, -90, -11, 38, 97, -76, 73, -5, -101, 90, -105, -94, 67, 74, 17, 58, -71, 120, -64, -42, 32, -78, -93, 118, -50, 53, 82, 44, -117, -17, 2, -108, 71, -88, -31, -14, 54, 110, 81, -8, -101, -17, -85, 15, 92, 93, 82, -68, 91, -50, -1, 5, 121, 112, -55, -64, -120, -49, -90, 121, -45, 119, -104, -28, -101, -46, -122, -11, -36, -2, -120, -58, -128, 7, -108, 26, -63, -63, 84, 23, -85, 32, -11, -80, -31, -44, -22, -124, 65, 4, -108, -15, 124, 35, 1, 96, 80, 12, 96, 39, -60, -48, -1, 59, -119, -6, 79, 31, 10, -76, -82, 18, -84, 17, 30, 47, 40, -54, 78, 1, -21, 32, -1, 121, -119, -60, 36, 109, -86, -92, -67, 45, -58, 107, -77, -27, 93, -111, 59, -120, 52, -79, 109, -62, 59, 57, 100, 66, 96, 31, 39, -101, 14, 80, 35, -95, -35, 79, 13, -107, -50, 2, -17, 59, -32, 15, -7, 45, 47, -12, -8, -96, -120, 123, 98, -57, -1, 76, -60, 20, 31, 51, 10, 127, 88, -52, -126, 56, 101, 55, 4, 94, -44, -9, -121, 70, 102, -41, -97, 11, 4, 18, 35, 4, 98, 114, -65, 91, -46, -17, -22, 88, 89, -73, -119, 9, -60, -25, 38, 115, -119, -51, 123, 82, 21, 100, -55, -3, 114, -20, -115, 102, 106, 85, -122, -118, -33, 80, -36, -99, -111, 109, -94, -121, -125, 95, -81, 78, 83, 1, 75, 84, -62, -39, 94, -21, 68, -3, -30, -2, 30, -57, 97, 74, 87, 55, -74, 113, -86, -97, -126, 31, 34, -103, -72, -14, -14, 61, 65, -85, 67, -57, -67, -107, 90, 51, 118, 57, -77, 48, -31, -13, 19, -56, -44, 39, -37, 43, 103, -24, 96, 45, -92, -57, -45, 113, -44, -106, -68, -120, -16, -30, 43, 39, 17, -104, -48, -123, 64, 32, 23, 121, -83, 43, -61, -17, -59, -64, -4, 72, 13, 92, -99, -24, -28, 80, -49, 99, 45, -75, -83, 86, -87, 71, -30, 10, -102, -109, 39, -86, 74, -29, -61, -95, -90, 106, 9, -63, -54, -58, 3, 7, 48, 89, -90, -24, -87, -80, 97, -34, 38, 104, 21, -103, -72, -59, -115, -128, 51, -69, 52, 20, -64, -8, 66, -91, 77, -112, -111, 84, 90, -16, -54, -26, -70, -108, 46, -32, 100, 71, 31, 2, 58, 90, -50, 27, 106, -60, -128, 11, 72, -125, 80, 97, 112, -110, -104, 91, 26, 103, 121, 43, 103, 97, 106, 34, -55, 5, -68, 23, 98, 82, 44, -120, -35, 33, 33, 91, -121, -9, -106, 34, 22, 30, 62, 20, -22, 31, 24, 14, -35, 23, 8, 16, 50, -19, 71, 47, -61, 81, 98, 18, -39, 18, -9, 106, 38, -59, -47, 39, -79, 68, -33, -67, 95, 110, -80, 14, 83, 39, 32, -103, -11, -39, 15, -38, 17, -10, 21, 109, -15, -25, -105, -128, -24, 85, 26, -18, -14, -90, -40, 62, 67, -103, 53, -109, -26, -126, -59, -58, -104, 107, -40, -15, 99, 35, 38, -15, 14, -122, -115, 83, -73, 48, 45, -74, -54, -70, 111, -22, 30, -1, -75, -8, 61, 62, 79, -32, -64, 84, -4, -64, -86, -21, 87, 9, 112, -26, -72, 20, 86, 85, 68, 84, -64, 94, 70, 102, -68, -19, -93, -33, 126, 48, 35, 10, -66, -97, -111, 124, 98, -40, -91, -12, 81, 90, -66, 88, -77, 41, -28, -51, 17, 60, 98, 31, -6, -76, 27, 23, 77, -115, 95, -112, -54, 54, 5, 120, 19, -111, 118, 115, 11, 87, 57, -9, -47, 57, 36, -84, -89, 90, -16, 105, 126, -13, -77, -89, 107, 45, -105, 51, -79, 85, -12, 70, -86, 63, 7, -30, -101, -35, -12, -117, 88, 55, -120, 59, 36, 56, 100, -117, -97, 48, 58, -34, 15, 79, -114, -99, 56, 86, 78, 29, 33, 127, 98, -16, -36, 19, -89, -22, 101, -85, 110, -100, -76, -101, 113, -71, -89, 80, -77, -91, 62, 52, 58, -22, -41, -105, -15, 118, -3, 87, 19, -14, 82, -78, -122, 70, 4, -19, -52, 16, -25, -18, 48, -15, -100, -98, -57, -106, 85, 62, -71, -127, -74, -113, 0, -96, 49, 98, -4, -114, 64, 16, -102, -90, 51, -74, 15, -121, -38, 28, 63, 99, -48, 60, 46, -39, -76, 7, 90, -23, 9, 111, -124, -29, -75, 78, -18, 20, 27, -94, -20, -100, 64, -4, -115, -30, -31, -51, -41, 120, -35, -34, 86, 49, -33, 16, 24, -35, -90, -91, -79, 18, 112, 91, 112, 15, -22, -47, 75, 74, -15, 45, 50, -127, 117, -67, 95, -61, -97, 50, -51, -122, 4, 106, 112, 65, -90, 101, -94, 5, 68, 17, 110, 97, -58, 114, -50, 5, 114, -114, -101, 123, -32, -126, -62, -62, -65, 63, 95, 10, -74, -53, 79, -6, 124, 118, 46, -90, 60, 67, 35, 17, -111, 102, 13, 25, -100, -118, -21, 81, 115, 21, 69, -68, 9, 107, 5, 72, -62, -14, -54, -128, -108, 49, -94, -44, -86, -13, -106, 53, -57, -17, -26, 118, -123, 96, -115, 95, -114, -78, 87, 63, -91, -35, 10, -70, -107, 22, -43, 6, -66, -12, -91, -40, -38, -15, 6, -26, -121, -102, -94, -125, 74, 48, -7, 84, 127, -79, -13, 108, -31, -13, 41, 80, 28, -68, -83, 107, 46, -37, -109, 52, 114, -27, -92, -76, 8, 55, 110, -39, 87, 113, -30, -76, 10, 88, 20, -113, 47, -87, -24, -39, -20, -113, -2, 56, 29, -100, 116, -74, -82, 101, 92, -73, 13, 108, -32, 65, -121, 13, -115, 96, 8, -54, -119, 87, -76, 35, 8, 36, -98, -116, 45, -77, -51, -69, -5, 60, -88, 24, 103, 79, 50, 114, -63, -54, 103, 78, -95, 7, -96, -119, -85, -53, -23, 98, -41, 115, -117, 31, 23, 93, 31, -78, -54, -116, 70, 9, 103, -11, 47, 5, -50, 24, -25, 69, 18, -79, -86, -47, 55, -61, -76, -46, -94, 103, 55, 110, 22, -106, -53, 110, -1, 77, 12, 16, 5, -6, -108, 72, -71, 74, -79, 82, 20, 106, -9, -91, -54, -74, -5, -16, 30, -68, 18, -48, 20, -2, 66, -18, 90, 123, 32, -8, -86, 56, -24, 17, -7, 118, -68, -124, 35, -43, 33, 24, 35, 62, -18, 112, -75, 19, -45, -12, 33, 66, 21, 78, 54, -80, 118, -74, 26, -80, 107, 99, -89, 119, 8, 4, -28, 82, 19, 28, 47, 35, -17, -19, -119, 120, -82, -54, -114, 68, 123, 7, 75, -105, 1, -44, 89, -44, 59, 64, -104, 61, 36, 88, 59, -29, -44, 71, -74, -120, 107, -80, -63, 17, -106, -39, 118, -95, 127, 89, 73, -71, 77, -87, -33, 83, 87, -65, 60, 66, -17, 67, -64, -55, 73, 9, -127, 47, -27, -122, 123, -77, 94, 15, -54, -11, -68, -98, -48, 94, -57, -71, 10, -44, 71, 12, 10, -72, -15, 71, 38, -10, -104, -25, -45, 17, -126, 15, -100, -29, 8, 48, -29, 111, -53, -127, 127, 36, -37, 27, -53, -39, 116, -98, 21, -14, -54, -74, -35, 112, -90, -123, -10, -4, -128, 125, -95, -125, 23, -121, -59, -33, -102, -6, -33, 107, 6, 93, 52, -91, -114, -67, 44, 62, 33, 80, -4, -69, -112, 83, 85, -103, -125, -121, 82, 22, 3, 10, -82, -68, 29, -9, 27, -36, -30, -36, -48, 118, 58, 33, -71, 56, 51, 52, 42, -108, -76, 5, -47, 2, 47, 25, 48, 29, -33, 61, 112, -58, 10, 69, 86, -3, -79, -124, -55, 11, -45, -8, 12, 9, 75, -8, -99, -36, 18, 77, -16, -109, -114, -27, -49, 65, -108, 15, -113, 78, 69, -73, 114, -106, 27, -104, -73, -4, 50, -67, -14, 67, -67, 73, 112, -125, -29, 77, -4, -106, 72, 5, -47, -14, -110, 39, 99, 41, -69, -26, 5, 126, -50, -7, -13, -85, -52, -47, -118, 124, -1, -102, -39, -28, -61, -90, -28, -39, -64, -4, -95, -3, 29, 61, -87, -111, -85, -60, -102, 104, -118, 113, -16, 110, -58, -34, 33, 86, -40, 104, -91, 74, 15, -81, 113, -102, 120, 40, 103, 41, 41, -35, -24, 103, -122, 101, 29, 122, 94, -83, 96, 112, -105, 94, 82, 72, -65, -6, 107, -58, 28, -96, 119, -12, 102, 120, 9, 127, -98, 21, 122, 95, 83, 118, -80, 114, 3, -9, 68, -8, 121, 117, -27, 98, -48, 91, 62, -33, -55, -118, 20, 22, -64, 11, 114, -52, 127, -111, 60, -119, 41, -92, 58, -87, 12, 8, -117, -106, -17, 53, -101, -124, -46, 91, 104, -24, -50, 74, -50, 32, 63, -91, 64, 107, 15, 16, -42, -115, -99, 73, -9, -125, 34, -128, -74, -114, 92, -86, 21, 84, -81, 12, -53, 13, 78, -14, -23, -52, -79, 74, 66, 30, -48, 88, 84, 43, 10, 2, 13, -106, -38, 97, -1, 90, 105, 105, -117, 54, 27, 2, 20, -93, 111, 118, -96, -19, -31, -44, -80, 102, 41, -85, 94, -112, 105, 22, -78, -88, 65, -99, -86, -39, -112, -109, -8, -61, -61, 93, 125, 85, -5, -50, -113, -46, -31, -23, -65, 37, -107, -54, -89, -39, 98, -51, 35, 54, 41, -8, 119, -22, 6, -37, 57, 90, 95, -85, -91, -113, 29, -94, -52, 61, 50, 78, -109, -107, -111, -34, 15, -75, -11, -108, -42, 78, 36, 60, 4, 101, -110, 69, -21, 84, -73, 50, -114, -77, -81, 117, -95, 109, 63, -73, 102, 101, 69, 102, 54, 80, -93, 68, -83, 39, 14, 52, 31, 39, 27, 71, -83, -31, 79, 22, -53, -111, -1, 83, -37, 91, 12, 79, -51, 92, 58, -79, -102, -87, -90, 59, 118, 56, 20, 76, 4, 80, 34, -108, -26, 126, -62, -127, 74, -92, 41, 49, 108, -68, 42, 1, -4, 8, -65, 20, 56, 37, -54, -64, 41, 2, 19, 87, -84, -36, -95, 46, -43, -12, -46, -4, -57, -35, 49, 63, 90, -5, -18, 69, -6, -65, 109, -128, 122, 9, -82, -36, 26, 38, 12, -114, 44, 14, 68, 7, 96, 50, 59, 127, 20, -46, -61, 64, 99, 98, 123, -62, -57, 123, -68, 111, -103, 59, 0, 125, -124, -88, 122, -106, -126, 72, -106, -93, 15, 41, -118, -127, -87, -64, -108, -122, -98, 121, 100, 104, 32, -24, -42, -70, -46, -27, -97, -15, 39, 12, 71, -88, -41, 50, -115, 109, -106, -22, -82, 46, 39, -20, 29, 84, -128, -78, 22, 46, 7, -64, 44, 76, -7, -84, 26, -43, -6, 33, 124, 41, -93, -106, 9, -32, 124, -65, -31, -27, -77, -88, -87, 91, 25, -52, 17, 69, 24, 26, -30, -98, 45, -47, 55, 83, 68, 43, 78, 18, 93, -23, -21, -28, -121, -42, 60, -41, 9, -26, 19, 46, 57, 87, 59, 69, 7, -20, -40, -12, -57, 106, -50, -101, -118, -111, -125, -43, -101, -29, -98, -118, 47, 63, -6, 53, 125, -85, 122, -42, -51, 91, -92, -83, -44, 105, -125, -49, -64, -45, 35, -73, -67, -23, -3, 107, -6, -57, 99, 103, -83, 24, -119, 38, 59, -80, 122, 50, 69, -100, -82, -94, 96, -24, 51, -124, -31, 16, -26, -122, -18, 112, 32, 92, 117, 95, 122, -92, -106, 82, -92, -116, 87, -22, -68, 103, 98, 87, 127, -58, 86, -66, -48, -63, 105, 122, 104, 25, 33, -31, 20, -61, -6, 41, 54, -13, 124, 38, -64, 115, -92, 119, -30, -44, 28, 116, -5, 22, -28, -19, -101, 82, 125, -120, -2, 123, 76, -126, -101, 104, 74, -60, -60, 33, 89, 121, 68, -30, 113, -53, 62, -10, -60, -63, 10, 38, -9, 67, -80, 38, -20, -94, 123, -72, -128, -40, 93, -123, 16, 43, -20, -103, 54, 63, 8, -43, -87, 5, -66, 15, 102, 41, 117, 38, 48, 116, -95, -113, -70, 28, -51, -68, 120, -56, -91, -73, -20, 11, -111, -24, -87, -98, -92, 30, -58, -42, 94, 114, 35, 91, -77, 72, 57, 29, -50, -123, 93, 126, -44, 79, -101, -58, 97, -89, 36, -55, 10, 99, 72, 106, 28, -81, 117, 29, -21, -65, 81, -93, -107, -64, 44, 70, 50, -93, 88, -37, -50, 105, -107, -78, 105, -109, -64, -73, -40, 112, 79, 114, -100, 113, 78, 102, 110, 105, 127, 52, 23, -69, 80, -63, -19, -47, -85, -91, 42, -59, -15, 34, -34, 44, -20, -69, -36, 84, 57, -13, 33, -77, -37, -3, 94, 32, -83, 6, 44, -59, -73, -80, 127, -18, 103, -56, -26, -95, -41, -125, 5, 115, -107, 89, -118, 50, -50, 89, -109, -80, -3, -7, 60, -25, 102, -37, -31, 117, -98, 63, -80, -38, -13, -69, 20, 16, -44, 106, -75, 52, -87, 88, -2, 114, 84, -95, -80, 99, 49, 30, 1, 71, 99, -30, -87, 109, 32, 26, 121, 49, -1, -4, -25, -75, -14, -3, 111, -17, -118, 42, -60, -60, -45, 31, 36, 103, -49, 114, -56, -123, -36, -118, 10, -55, 43, 31, -51, 97, -26, 100, 30, -63, -31, -56, -116, 68, 37, -81, -115, 45, 24, -49, 103, 7, 49, 97, 2, -84, -96, -23, 119, -20, -55, -78, 94, -8, 68, -86, -66, 61, 60, 13, 53, -87, 93, -56, 102, -99, -18, 100, -34, 3, -57, -40, 65, 43, 46, 85, 101, -111, -84, 54, -94, -119, 87, 65, 96, -92, 53, 56, -20, -80, -36, 113, -46, 114, -116, 95, -2, -127, 26, 25, -3, 45, 38, -128, 123, -102, 30, 58, -61, 58, -25, -119, 14, 108, -27, -88, 77, 66, -72, -112, 25, 19, 103, -103, -50, -113, -8, 11, 52, 32, -66, -44, 102, 46, 12, -45, 28, -62, 20, 73, -61, -43, 122, 53, -37, -25, 0, 90, 78, 108, -72, -105, -26, 42, -98, 38, 93, 0, -121, -61, 11, 19, 113, 72, -48, 99, -60, -37, -18, 55, 5, -70, -14, 55, -34, 70, 65, 23, -47, -41, 87, -43, -84, 53, 69, 119, 37, -24, 99, -55, -22, 35, -100, -108, 28, 20, 104, -16, -114, 28, -32, -37, 82, -75, 63, -27, -69, -9, 58, -16, -60, -6, 106, -75, -75, 5, 2, -110, 65, -82, -5, 90, 60, -35, 17, 52, 116, 120, -30, -93, -101, -88, -64, 46, 20, -27, -84, -80, 21, 115, -127, 121, 45, 38, 40, -17, 26, -88, 105, -91, 45, 15, -107, -90, 61, -128, -75, -69, -21, -56, 31, 72, -12, 96, 122, -94, -52, -107, -68, -4, -108, -25, -51, -65, 83, 100, 90, 103, 45, -115, -68, -1, 73, -36, -25, -13, -93, -114, -45, 62, 3, 80, 21, 71, -2, -105, 49, 40, 60, 94, 67, -39, -23, -122, 16, -22, 72, -101, -91, -104, 48, -128, -79, -123, -19, 126, -57, -43, 89, 37, 15, -114, -15, -80, -47, -38, -18, 42, 98, -123, 124, 95, 5, -96, -54, 31, -87, -64, 111, 98, -125, 14, 86, 88, -74, -54, -121, 3, -10, 105, -49, -69, -107, 98, -92, 35, 19, -32, -81, 55, 37, -116, -5, -73, 97, 61, 104, -103, 85, -89, -77, -64, -99, -99, -4, -96, 105, 47, -87, 118, -119, 79, -88, -113, -13, 49, 94, 78, -80, -80, 75, 53, 78, 22, 15, 18, -113, 56, -106, 48, -77, 0, -38, -19, 4, 0, 64, 28, 110, -91, 87, -117, 65, -67, 21, 41, 72, -35, 97, 109, -83, -39, 108, -22, -117, 5, -6, 101, 76, 72, -71, -116, -2, 89, 66, 73, 18, -21, 20, -98, 72, 14, -3, -126, 58, -35, 71, -125, 54, 59, 81, 33, 5, 40, 93, 118, -66, 90, -32, 31, 19, 102, -120, 25, 112, 122, -83, 60, -90, -115, 119, 0, 57, 18, -73, -35, 96, 67, 66, -88, -75, 113, 83, -70, -38, -84, -124, -12, -20, -78, -15, -111, 50, -20, -36, 66, -58, 107, -74, 80, 109, -45, -51, -108, 94, 54, -54, -33, 22, -88, 119, 24, 71, -27, -60, -74, -124, -6, -86, 13, -13, -7, -100, 90, 31, 38, -57, -18, -74, -81, -123, 103, 57, 30, 4, -98, 76, 39, 57, -90, 29, 87, -41, 57, -64, 126, 32, -74, -91, 118, -57, 123, 116, 26, 99, 101, -70, -86, -91, -117, -88, -31, -108, -86, -11, -52, 116, 108, -9, -34, 118, -95, -43, -7, -57, -59, -27, 44, 84, 105, -21, 31, 67, -111, 112, 91, -75, 77, 43, -89, 27, -84, -4, 91, 0, 71, 53, -95, -118, -114, -15, 17, 76, -32, 36, 106, -59, 98, 39, 46, -22, 85, -21, 123, 61, 98, 40, 74, -28, 28, -86, -63, 96, -98, -114, -108, -45, -33, 54, -65, -2, 36, 53, -31, 3, 106, 16, 123, -43, 73, 13, -98, -55, 98, 9, 31, 64, 57, -84, -7, -35, 0, -84, 107, -54, -51, -94, 51, -125, 63, -114, -18, 55, -24, 81, -77, 14, 72, 51, -26, 104, 119, -67, -60, 75, -124, -110, 89, 58, -70, -27, -6, -27, 21, -102, -42, 66, -65, -73, -58, 20, 99, -50, 54, -23, 69, 103, -118, -106, -53, 14, 51, -107, 50, -94, 64, -103, -18, 66, 7, 38, -45, 100, -17, 106, 10, 24, 42, 103, -101, -51, -104, -78, 87, -52, -26, 41, -12, -100, -82, 4, -6, -28, 1, 93, -2, 14, 93, -33, 77, -83, -56, 66, -10, -43, 7, -7, 22, -56, -71, -49, -97, -14, -96, 63, 21, 59, -78, 56, 123, 13, 89, -87, 7, 23, 84, -99, -6, -63, 71, -99, -13, -102, -64, -7, 111, -107, -86, -81, 78, 100, 86, 115, 95, 34, 102, -109, 17, 29, -124, 96, 39, 95, 95, -35, -92, -12, 70, -7, 117, 24, 127, 62, -41, 116, -59, -112, -83, 26, -120, 15, -81, 78, 51, -2, 8, -28, 89, -18, -97, 75, -23, -102, -102, 73, -57, 100, -85, 88, 17, 76, 66, -81, 33, 86, -99, -29, 15, -26, 11, 124, -16, 25, 113, 91, 78, 54, 57, -79, -69, -70, -71, 73, 119, -103, -121, 56, 56, 23, -99, 104, 26, 110, -20, -27, 71, 110, -9, -29, 50, -43, 36, -23, -54, 2, -13, -126, 111, -57, 80, 125, -48, -4, -72, -13, 77, 120, 51, 23, 66, 92, -39, -111, 55, 110, -35, 24, -20, 64, -126, 86, 56, 105, 83, -57, 108, -15, -60, 44, 113, -4, -70, -101, -111, 7, -57, 113, 27, 27, -60, -77, 53, 19, 125, -128, 101, -32, 16, 126, -13, 3, 59, -21, -77, 119, -90, 62, 16, 25, -107, 33, -24, -123, -66, -98, -64, -107, -116, 74, 53, 21, 42, 112, 116, -83, 21, -119, -24, 125, -61, -40, 43, -118, 45, 114, 28, -115, 23, -46, 30, -124, -62, 59, -8, 7, 109, 62, -57, -108, 76, -54, -39, -38, 60, 101, 68, 62, 24, 53, -43, -31, 21, -106, 88, -50, 126, -82, 82, -34, 73, 89, -58, -119, -25, 60, -123, 113, -11, 127, -45, -18, -44, 91, 25, 122, -80, 80, -50, 58, -60, 43, 13, 115, -120, -53, -3, -75, -55, 86, -37, -91, 74, 88, 81, 77, -9, -42, 17, 95, -14, -128, 44, -90, 20, -92, -78, -12, 54, 5, 72, 86, 18, -42, -116, 7, -29, 24, 58, -123, 57, -94, -53, 109, 38, -61, 74, -111, -29, -103, 111, 12, 88, -51, -55, 66, 65, 58, -49, -114, -74, 46, 61, 63, -126, -69, -11, -32, -128, 9, 108, -111, -28, -47, -2, -36, -86, 3, -82, -98, -24, -104, -44, 90, -34, 41, -127, -31, 13, 115, -83, -8, 70, -96, 34, -8, 45, 108, 115, -18, 107, -83, 47, -33, 25, -83, -99, -48, -104, 21, -55, -16, 2, -116, -122, -85, -32, -69, -105, 102, 38, 4, 34, 102, -21, 84, 78, -119, -4, 56, 3, 65, 98, -40, -61, 62, -12, 1, -93, -89, -38, 126, -34, -59, 99, 74, -117, -93, -100, -31, 30, -106, -58, -78, -14, -100, -54, 27, 84, 124, 18, -124, -59, 67, -79, -34, -43, 118, -76, -107, -59, 75, -11, -109, -106, -23, -115, 94, 1, -7, 17, -6, -90, 77, 41, 1, -127, -70, -127, 90, -84, -91, 41, -66, -81, -76, -14, 107, 104, -16, 79, -111, 81, -18, 35, 124, 95, 96, -120, 118, -99, 126, 39, 40, -60, -41, 109, -53, -125, 76, 109, -103, -66, -93, 103, 55, 111, -55, -4, 113, -41, 95, -6, 30, -102, 37, 89, -91, -23, -77, 0, 119, -56, 4, 42, -107, -11, -69, 44, 76, 38, -66, 121, 119, 77, -34, 12, 32, -37, 36, 110, -69, -15, 92, -10, 23, 79, 121, 3, -87, -117, -60, -99, -3, -123, 76, -105, 102, 50, -56, -122, -122, 64, -43, -11, -82, 88, -58, -95, 3, 37, 92, 21, 79, 11, 39, -15, 19, 124, 90, -39, -73, -65, -78, 60, -127, 39, -98, 42, -35, -72, -48, -40, -87, -26, 77, 127, 114, -63, -85, 65, -10, -111, 13, -72, 38, -41, 106, -26, 77, -48, 39, -57, -57, -2, 16, 8, 14, 11, 79, -62, 126, 20, 115, 4, -122, -89, -47, -68, -75, -89, -40, -32, -80, -119, 39, -81, 117, 83, 68, 44, -55, -96, -7, 127, 74, 76, -60, 64, 106, -123, 71, 35, 33, -110, 126, -25, -102, 12, -78, 122, 18, -110, 24, -66, 39, 18, -63, -127, -26, 67, 112, -61, -5, -55, -126, 51, -23, -100, 39, -32, 10, -76, -2, -47, -96, 63, 7, 103, -74, -33, 120, -76, -94, 114, 96, 23, -93, 69, -18, -68, 81, -112, 123, -86, 122, 62, 122, 4, -9, 24, -94, -37, -77, 112, 82, -77, -20, 69, -1, -60, 105, 90, 66, -98, -48, 9, -10, -96, 67, 34, -90, -8, 107, -93, -99, 4, 19, -24, 94, -56, -45, -106, 124, 107, 102, 11, 48, -33, 97, 40, 108, 15, 74, -49, -25, 58, -84, -88, 20, -42, 55, -98, 5, -77, -35, 101, 59, 89, 122, 49, -1, -61, -74, -85, 43, 46, -115, 86, -73, -22, -54, -26, 11, 10, 16, -29, 7, 106, 82, 55, 18, 101, 45, 20, -79, -35, 66, -53, 95, -74, 87, -23, 91, -124, -90, 120, -75, -19, 82, -76, -42, -64, -43, 24, -67, 115, -105, 73, 80, 66, 122, -18, -72, 14, 15, 37, 80, 39, 27, 54, -118, 112, -29, -3, -37, -87, -120, -85, -6, 95, 43, -22, -91, 1, 55, -69, 50, 43, 39, 23, 115, 74, 62, 46, 32, 108, -8, 30, 116, -55, 20, 118, 36, 111, -95, -1, 1, -121, 5, -51, 52, -73, -8, -15, -122, -100, 19, 22, 101, 34, 107, 79, 59, 49, -21, 107, -107, 20, -47, 52, -24, -52, -27, -79, -83, -93, -15, 35, 11, 116, 80, -120, -3, -111, 25, 87, 109, 121, -67, -89, -25, 32, -88, -62, 26, 125, -73, 103, 50, 78, 46, -107, -54, 50, -49, -52, 88, 69, 66, 34, -15, -93, -72, 106, -101, -116, -101, 91, 19, 26, -22, -102, -79, 11, 69, 47, -95, -41, -83, 19, 93, 20, -9, -46, 29, 87, -22, -116, -35, -102, -5, 87, -77, -125, -97, 114, 41, -120, -99, -85, 11, -12, 33, 37, 77, -127, -90, -36, -78, 63, -15, 43, -61, -38, -20, 94, 30, -86, -6, -19, -119, -126, -31, 45, -40, 105, 106, 113, -109, -68, -114, -21, -57, -102, -89, -105, 61, 2, -1, -6, -118, 66, 114, -66, -95, -42, -27, -61, -71, 60, -57, -16, -21, 57, 55, 112, -31, -93, 20, 30, -55, -90, -25, -115, -110, 118, 94, -82, -89, -23, 127, 15, 0, 70, 127, -72, -80, -14, 126, -6, 90, 40, -9, 14, -73, -45, 84, 81, -26, -52, 119, 84, 28, 20, 89, 48, -88, -116, 24, 11, 45, -90, -73, -46, 123, -63, 91, -14, -43, -127, 78, -1, 107, -93, 69, -2, 70, 80, -22, 69, -59, 124, 9, -35, 102, 102, -59, -91, 111, 62, 5, -42, -43, 113, -103, -10, 12, 38, 27, -2, 14, -95, -48, 15, -36, 94, -55, -3, 124, 40, -103, 8, 40, 83, 9, 102, 119, 53, -83, 57, -75, -113, 27, -108, 107, -47, 34, 2, 61, 10, 1, -4, -98, -59, 119, 100, -91, 34, -64, -64, -15, -83, -55, 81, 49, 76, 79, 123, -44, -80, 77, -77, -107, 95, -40, 74, -11, -54, 38, 21, -17, 93, -108, 86, -58, 9, 39, 58, -76, -45, 20, -102, 4, -69, 97, 119, 24, 78, 59, -101, -26, 32, 116, -101, -60, -49, 5, -77, -85, 112, 74, 37, -48, -44, 91, 55, -7, -81, -9, -4, -98, 17, 106, -91, -34, -52, -13, 43, -1, -99, -94, -59, -39, 79, 3, -111, -23, -70, 50, -61, -30, -100, -86, -9, 68, 121, 78, -60, -116, -45, -4, 35, -39, 21, -26, 21, -66, -55, 9, -127, -21, 115, -121, 21, -87, -15, -102, -60, -8, 106, -16, -25, 115, 29, 73, -40, 83, 59, -66, 116, 111, 29, -74, -46, 83, -5, -93, -91, 7, 114, -14, -36, -124, -38, 123, 123, -53, -33, -113, -37, 108, 19, -97, -1, -61, 38, -109, 117, 29, 24, 2, -93, -89, 124, 72, 3, -63, 75, -13, 70, -104, -119, 116, 7, 68, 44, 5, -97, 62, 72, -38, -16, 103, -116, -4, 108, 9, -22, -48, -61, 5, 57, 126, 39, 61, 20, 68, 45, -19, -29, -40, -8, -43, -105, 2, -114, 3, 117, 34, 82, 73, -19, -22, -59, -104, -93, 112, 103, 80, 126, -68, -19, 41, -46, -22, -100, 21, 36, -47, 127, -27, 58, -4, 73, 44, -63, 13, 21, 14, -40, 0, 85, -105, 67, 105, 0, 118, 126, -74, -6, 100, 71, 106, 17, -12, -60, -127, 55, -16, 9, 10, 107, 6, 37, 80, 31, -7, -101, 94, 19, -76, -48, 22, -73, -78, 41, -25, -8, 21, 110, 96, 31, 60, -124, -84, 75, 50, 54, -43, -93, -20, 14, 57, 64, -18, 100, 56, 114, -99, -80, -63, 88, -40, -108, 62, -68, 76, 122, -40, -95, -105, -74, 25, -79, 107, -18, 107, 30, 98, -13, 30, -101, 71, -18, 37, -80, -96, -119, -74, -59, 40, 84, -88, -91, -62, 5, 12, -123, 88, -84, 121, 11, -94, -87, -64, 86, -26, -24, 88, 12, -87, -92, 39, -11, 12, 107, 84, -63, -110, 123, 7, -77, 93, 0, -114, -76, -61, -128, 76, -84, 53, 84, -111, -58, 103, 101, -65, 47, -80, 40, -79, -51, 24, -27, 66, -54, 76, 80, -69, 89, -62, 109, 1, 122, 120, 13, -81, -124, -109, 104, 48, 53, -92, 66, -72, -108, -125, -98, -97, -108, -45, -122, 39, 98, -123, 75, 91, 58, -52, -106, -29, 35, -109, -123, -10, 101, -5, 34, 18, 16, -43, 103, 83, -98, 111, -73, 35, 73, 17, -120, -93, -106, -4, -106, -108, -104, 79, -49, 105, -83, -73, -30, 103, -32, -47, 55, -114, 40, 127, -26, -11, -48, -92, 112, -110, -128, 66, -32, 95, 22, 73, 68, 78, 9, 78, -76, 14, -36, 102, 101, -74, 5, -29, 21, -61, 61, 60, -78, 100, 112, 114, 34, -68, -13, -87, 108, -16, -3, -49, -102, 66, 110, -10, -100, -11, -89, 80, 0, 5, -125, 58, -11, 15, 115, 3, 49, 52, 69, 73, 5, -109, -57, 67, -42, 92, -101, 82, -92, 93, 126, 21, 42, -49, 108, 29, -25, -22, 115, 115, -37, -102, -16, 73, 77, 29, -52, -84, 53, -28, -68, 118, -59, 23, 34, 110, 87, -95, 70, 61, -75, -95, 109, 113, -128, -40, 106, -3, -32, 32, 22, -72, 117, -45, -69, -90, -81, -122, -59, -28, -34, -101, -25, 75, -96, -87, -99, -7, -33, -82, -53, 47, 112, 16, 118, 60, -27, -2, 108, 34, 86, -94, 107, 43, -30, -88, 43, 25, 89, 104, -19, -88, 120, 73, -94, -120, 76, 29, -121, 44, 1, -92, -40, 82, 19, 8, 84, 19, 33, 25, 57, -118, -124, -14, -116, 53, -12, -88, -41, -70, 25, 119, -125, 48, -115, 3, 89, -107, -98, -91, -125, 26, 80, 117, -88, -108, 23, 97, 30, -17, -118, -37, -20, 57, 81, 38, -108, -105, 1, -83, 91, 70, -60, 125, -7, 114, -19, 120, -76, -80, 85, 126, 120, -20, 126, -17, 48, 95, -37, -72, 53, 75, 63, -97, 58, -21, -6, 111, 2, 105, 118, 39, 47, 68, 113, 112, 123, 45, -30, -53, -28, 46, 61, 56, -83, 117, -39, -64, 16, 57, -108, 29, 18, -96, -125, -108, 111, -90, 90, -37, -59, 40, 62, -93, 35, -14, 4, -50, -39, -79, -18, 16, -1, -30, -14, 40, -53, 124, 54, 105, 125, -18, -86, -124, 84, -40, 92, -75, 76, -69, -56, 111, 54, 118, 121, -59, -64, -67, -98, 46, 93, 79, -44, -48, -99, -42, 8, 112, -106, -4, 58, -78, 123, -77, -63, -14, 33, -20, -85, -46, -101, -32, -97, 37, 8, -42, -12, -128, -53, 91, 26, -22, -89, 18, 91, -60, -92, -20, -117, 47, 99, -93, 8, -24, -30, 98, -114, 2, -54, 114, 106, 99, 44, 50, 7, -44, -102, 11, -75, -67, 57, -6, -8, -25, 97, 53, 123, 121, 23, 118, -36, -1, 25, 110, -10, -105, -42, 13, -23, -55, -28, 126, 115, -95, 126, -39, 96, -125, -33, -124, 47, -49, 19, -113, 18, 88, -102, -82, -60, 70, -9, -47, 92, -84, 60, 26, 90, -123, -52, 111, -97, 7, 51, -88, 75, -118, 0, 89, -127, -52, 31, 71, 52, -15, 21, 47, -20, -21, -35, 124, 8, 4, 77, -125, -124, 5, -22, -4, 62, 48, -108, 87, 115, -79, 126, 52, -15, 3, 36, 108, 124, 2, -91, -21, 61, -48, -58, -25, 92, 63, 113, -112, -68, -117, 75, -17, -57, -33, -88, -42, 79, -84, 102, -7, -128, 96, -92, 97, 51, 99, 91, 76, 77, 43, 84, 50, -43, 47, -119, -120, -73, -15, -48, -5, 108, 74, -104, -54, 57, -41, -116, -99, -100, 110, -43, -31, -81, -75, 28, 9, 34, -81, 50, -5, 4, 0, 20, -90, 67, -29, 103, -123, -93, -90, -54, 25, -109, 16, 112, -96, 107, -60, 125, 12, -28, -7, -88, 78, 36, 55, 34, -90, 32, -20, 72, 63, -13, 27, 63, -29, -48, -67, -47, 16, -43, 25, -57, 88, -46, -71, -90, 85, -99, 98, 69, -79, -51, -101, -118, 74, 105, 39, -53, -125, 119, 51, 53, 31, 19, -22, 84, -4, -123, -3, -91, -1, -44, -83, 119, 69, 107, -26, 70, 49, 94, -106, -105, 2, -122, -35, -85, 102, -46, -94, 119, -92, 65, 32, 38, 67, 58, 5, -17, -22, -77, 36, 27, -50, -38, 82, 31, -50, 73, 96, 78, 60, -1, 97, -22, -36, 34, 116, -54, 5, 67, -46, -65, 50, -79, -71, -7, 22, 27, -119, -72, -43, -47, -50, -73, 44, -32, 67, -106, -90, 52, 8, -124, 116, 23, 89, -108, 119, -24, -87, -92, 45, 125, -82, -34, -69, -47, 112, -113, 47, -65, -1, 81, 89, -85, -44, -86, 122, -36, -90, 103, 15, -79, 5, 5, -97, 74, -52, 53, -63, -8, -104, -126, -89, -64, 53, -53, 14, 95, 10, 96, 64, -108, 103, 40, 69, 31, -1, 3, -93, 34, 93, 20, 104, -86, -34, 101, -8, -46, -128, -126, 44, 14, -72, -68, 95, 7, -29, 56, 125, -125, 12, 28, 72, 110, 32, -27, -101, 35, 109, 97, 102, -36, 76, 105, 62, -83, 104, -125, -33, -32, -102, -116, -62, 65, -11, -99, 104, 101, 26, -36, -120, -40, -11, 66, 26, 46, 10, -32, 109, -62, -7, 24, 102, -1, 114, -18, -87, 51, 83, -116, 76, 114, 35, -20, -29, 126, -10, 18, -93, 34, -32, 72, -101, -118, -1, 68, 54, -31, 33, -97, -23, 31, -8, 1, -40, -99, 25, 44, 126, 102, 45, -72, -118, 4, 25, 118, 85, -97, -114, -19, -99, -98, -70, 9, -24, -93, -23, 69, -11, -82, 51, 25, -70, 103, -26, 8, -120, -125, 45, 33, -18, -115, -84, -101, -104, 43, 108, -116, 99, -93, -45, 30, -48, -127, -41, 61, 113, -112, 52, 70, -94, 69, -5, -70, 79, 56, -81, -44, 87, -45, 118, 96, -17, -44, 116, -8, 23, -114, -68, 93, 113, 82, -125, -50, 88, -42, 117, -109, -15, 74, 54, 31, 125, -31, 60, -90, 1, 14, -51, -87, 87, -86, -103, -125, -60, -62, -35, 44, -48, -118, -94, -62, 1, -26, 32, 2, 5, 14, 19, -13, -120, 67, -78, -40, 117, 43, -97, 99, 19, 93, -90, 27, -29, -92, -74, 15, 69, 42, -21, 27, -11, -86, 59, -117, -105, -16, 108, -121, 73, -98, -53, 76, 80, 51, -53, -24, -47, -33, -52, 74, 55, 66, -83, -53, -2, -119, 90, 116, -24, -50, -77, -105, -85, 2, 8, 115, -38, -1, 67, -110, -81, -11, -110, -48, 101, -50, 55, 49, -117, -27, -7, -102, -83, 75, -57, 79, -79, -48, -91, -24, 98, 13, 46, -50, -48, 99, 69, -8, -127, -31, -75, 47, 80, -124, -103, 62, 111, -69, -12, 87, 16, 76, 47, -18, 27, 53, -64, 35, -66, 26, 35, -112, -103, 49, -78, 36, -127, -51, -89, -99, 28, 107, -40, -25, 37, -96, 26, 96, -75, -13, 6, -22, -86, 59, -36, -46, 127, -14, 56, 52, 90, 66, -124, 115, -105, 36, -8, -113, 74, 26, 74, -96, -103, -125, 14, 52, -110, 87, 88, -3, -29, 122, 62, 69, 117, 84, -27, -105, 48, -24, -31, -122, 20, -82, -105, 87, 97, 97, -98, 93, -38, 60, 89, -51, -90, 93, 60, -74, -64, -97, -126, -19, -34, 82, -40, -53, 46, -41, -82, -37, -14, -13, -57, 126, 7, -34, -85, 60, -102, 84, -30, 44, -57, 58, -36, -25, 0, -66, -56, -5, -61, -69, -96, -124, -110, 74, 112, 81, -75, 60, 16, 24, 69, -71, 13, -15, -70, 65, -110, 48, -8, -68, -12, 71, -39, 58, -67, -22, 72, -11, 29, -76, 96, -39, 44, 12, 114, -73, -122, 24, 124, 3, 96, -54, 12, 119, 8, 59, 102, 32, -67, 61, -46, 25, 58, 29, -58, -98, 24, -55, -49, -57, 121, 37, 43, 17, -45, -71, 29, 67, 20, 104, -124, 3, 90, 39, 104, -122, 37, -112, -42, -69, -104, 35, -73, 9, 122, 31, 104, 88, -77, 70, -83, -105, 73, 77, 112, 21, 57, -67, -11, 96, 116, -36, 125, -81, 40, 91, -6, 115, -73, 78, -93, -46, 106, -115, 97, 103, 103, 93, -123, 110, 94, 21, -37, 112, -61, 56, -36, 2, 24, 33, 117, -15, 72, -122, -10, -69, -8, 24, 78, 51, 11, 125, 107, 123, 20, -46, 83, 29, 26, -68, -115, -12, -105, -113, 11, -63, -23, 126, -59, -9, -1, -61, -111, -43, -88, -59, 58, 6, -74, 68, 22, 110, 61, -70, -121, -22, 35, 96, -24, -8, -63, -96, 45, -59, -2, -73, -23, 114, 123, 52, 18, 61, 109, 81, -23, -20, 83, -93, 39, 30, -99, 90, -7, 69, 56, -25, 45, 25, 118, -71, -100, 13, -11, 124, -28, 66, 79, 82, -52, -85, 64, 125, -19, -93, 87, 54, 76, -107, 102, -114, 60, 101, 84, 38, -42, 20, 102, 100, -125, -35, -118, -40, 24, 70, -50, -126, 105, 87, 34, 86, -51, 111, -58, 51, -3, -11, 105, -27, 68, -49, -15, 77, -102, 39, 33, -125, -72, -40, 52, -119, 4, 24, 0, 97, -73, 113, -27, -81, -1, 87, -102, -57, -105, -110, 53, 93, -34, 60, -81, 7, -35, -94, -37, 114, -62, -111, -74, 17, 23, 99, -6, -50, -49, 113, -50, -15, 88, 2, 88, -62, 13, 29, 63, 40, 22, -66, -106, -7, -42, -68, -67, -32, 97, -111, -112, -115, -19, -34, -40, 74, 87, -65, 83, 89, -89, 26, 16, -47, 17, 121, 123, 99, -126, -58, -63, 92, -51, -75, -25, -82, -79, -83, -86, -77, -99, -104, -69, 27, -24, -123, -45, -66, -73, 114, 95, 83, -39, -86, -45, 17, 64, 116, 118, -71, 28, -57, -64, -37, 50, 15, -40, 39, 23, 8, -54, -124, -43, 85, 122, 92, 50, -127, 113, -34, 92, -10, 111, -50, -30, -116, -89, 112, 31, 65, -82, 62, 41, -107, -108, -68, -57, -50, 24, -2, 121, -3, -98, 118, -35, -123, 87, -66, -77, 106, 21, -16, 74, -93, -104, -103, -24, 72, 49, 12, 85, -128, 75, -126, 6, -67, 85, 125, 52, 15, 104, -36, 96, -8, -99, 115, 127, -70, 10, -112, -67, 74, 100, 52, -71, 44, 25, -115, -65, -40, -125, 43, 71, -2, 44, 38, 59, -104, -118, 15, -113, 127, 96, -104, -34, 55, -55, 115, 34, -33, 26, -23, 77, 91, 67, 116, -50, 7, 109, -34, 68, 16, 122, 120, -81, 108, 106, 93, -7, -44, 90, -38, 111, 24, -101, -123, -58, -85, 16, -108, -82, 56, -94, -62, -121, -49, -52, 108, -100, 124, 3, 69, 101, 64, -12, -63, -3, -82, 27, -102, -16, -79, 70, -55, -103, 99, 27, -72, -105, -79, 68, 113, -37, 64, 68, 50, -73, -31, -90, -59, -38, -17, -96, -105, 111, -45, -103, -98, -99, 96, 87, 61, 101, 84, -81, 59, 66, -104, -21, -24, -98, -82, -16, 81, -73, -21, -97, -1, -71, 8, -8, -7, 95, 117, -101, -102, -42, -41, 106, 84, -124, -10, -68, -8, 34, 65, -18, -12, -72, -45, 79, -61, 16, -27, 45, 72, 3, -27, -84, -15, -26, 8, 76, 126, 69, -86, 5, 13, 78, -69, 24, 92, 33, -11, -8, 78, 27, -92, -59, 101, 49, 32, -10, -96, -42, 103, -9, -111, -113, 23, -64, -26, -123, -18, 95, -61, 100, -121, -125, -117, -62, 23, -48, 36, 13, -6, -45, -118, 18, 10, -22, -80, -125, -72, -10, 47, 110, 74, -85, 45, 53, 89, -59, 67, 18, -119, -82, 63, 81, 41, 102, -3, 58, -7, 103, -67, 74, 106, 12, -60, -75, -34, 1, 93, 33, -57, -1, 4, 124, -84, -42, 57, -57, 79, 53, 69, 87, 64, -13, -76, 97, -54, -18, -98, -104, -77, -39, 119, 63, -16, -54, -23, 50, 0, -90, -34, 101, -58, -120, -42, -42, -45, -59, 1, -38, -120, -83, 111, -46, 70, -79, -82, -59, 93, -65, -16, -114, -34, 104, 3, -89, 96, 76, 114, -15, 53, 108, 72, -94, 100, -89, 6, 29, 47, -31, -99, -119, 105, 18, 70, -38, 58, -65, -3, -125, 119, -32, -72, -54, 34, 117, 61, -18, -74, 55, 37, 63, -107, -44, -114, -7, 77, 112, -99, 69, 108, 91, -6, -59, -83, -6, -91, -93, 73, -105, -99, 61, 47, 16, 80, -82, 58, 17, 2, 75, 57, 105, -99, 93, 18, 50, 55, 101, -70, 99, -57, 5, -27, 68, 98, 68, -60, -37, 78, 119, 107, -49, 31, -21, 78, 40, -35, -85, 25, -55, 124, 123, 121, 68, -83, 93, 68, -126, -82, -71, 53, -108, -57, 40, 17, -125, -31, 115, -113, 28, 50, 28, 89, 71, 69, -58, -77, 116, -93, -45, -86, 29, 14, 57, 90, 40, 26, 74, 115, -28, -118, 77, 72, -108, -37, 100, 91, 30, -23, 69, -49, -11, 69, -120, 27, 34, -27, -104, 19, -22, 8, -52, 71, -115, 84, 23, 79, 58, 103, 29, 66, -113, -117, 80, 57, -41, -119, -60, 87, -118, -80, 119, -100, -42, 35, 56, -29, 67, 69, -56, 0, 11, -21, 127, 104, -39, 65, 117, 12, 85, 110, 51, 105, 7, -20, -125, -113, 60, 108, 59, -85, 13, -10, 54, 92, -28, -69, 7, -50, -82, 6, -8, -97, 26, -87, 42, 120, 115, 107, 4, 33, -24, -117, -1, -39, -77, 31, -44, 68, -42, 119, 112, -111, -89, -15, 90, 4, 84, 74, -53, -39, -38, 29, -26, -114, 9, 34, -113, 13, -55, -80, 92, -74, -83, -45, -106, -6, 29, -125, 114, -97, -118, 76, 88, -26, -19, -57, 61, 72, 85, -50, 121, -15, 52, -115, -93, -29, 94, -35, -81, -125, 119, -29, -96, -47, 56, -77, 42, 31, 19, -118, -30, -29, -87, 18, 109, -58, 41, 114, -30, -32, 126, -6, 79, 60, -123, 50, -28, -35, -32, -25, 29, -36, 120, -70, 69, 87, 25, 58, -70, -6, 67, 113, 12, -42, 7, 51, 94, -126, -67, -37, 111, -118, -109, -72, 64, -70, -21, -33, 121, -84, -67, -84, 54, 73, 80, -44, 115, 10, 86, 17, -51, -93, 22, 39, -112, -43, -92, 103, 93, 49, 83, -15, 62, -85, 100, 81, -3, 119, 84, -81, 6, -15, 98, 3, -67, 34, 124, 30, 1, 36, -39, 34, 103, 71, 50, 2, 33, -100, 82, 9, 64, 100, 79, 10, 63, -66, 112, -85, 31, 29, -22, -53, 51, 125, -55, -39, -40, 102, -100, -73, 111, 44, 51, 52, -59, 106, -79, 38, 18, -122, -30, -51, -40, -58, 53, 112, 105, 25, 36, 54, -12, 2, -5, 61, 35, -3, -56, 77, 42, -68, -76, -102, 17, 102, -21, 111, -126, -81, -9, 109, -112, -49, -38, -55, -24, -66, 110, 73, -124, 16, 119, 13, -50, 37, -110, -106, -63, -60, 4, -93, 22, 90, 16, 121, -53, -84, 55, -117, 103, -55, -90, -65, -63, 37, -82, -30, 111, 58, -21, -75, -72, -57, -63, 93, 97, -99, -68, -24, -90, 101, 48, -107, -123, 78, 10, 29, -6, 126, 84, 49, -50, 35, -80, -76, -68, 127, 6, 12, 97, -33, -36, 58, 6, 103, 65, 63, -64, 86, 107, 43, -9, -20, 120, -105, 34, 22, 12, -59, 78, -77, -31, 33, 65, 66, 60, -24, 126, 6, 26, -128, 17, -8, 103, -101, 108, -128, 98, 33, -113, 110, -8, 120, -38, 52, 4, -33, 24, -21, -35, -58, -26, 27, 53, 4, -114, -57, 94, -49, -24, 10, -114, -123, 124, -49, -9, -78, -68, -71, -70, -19, 111, -85, -60, 114, 72, 49, 25, 43, 16, -29, 117, -41, 59, 45, -120, -40, -30, -103, 53, -74, -107, 74, 21, 120, -22, 75, -122, -3, 106, 100, 15, 108, -28, 73, 33, 40, -103, 126, -70, 77, -48, -24, 60, 60, -20, -127, -16, -54, -71, -97, -98, 97, 2, 108, -99, 58, -56, 121, -107, -1, -12, 61, 66, -86, 5, 90, 112, 19, -8, 95, -41, -6, 23, -63, 43, -109, -28, -47, 48, -56, -84, -57, 13, 0, 108, -103, 72, 109, -30, 27, -75, -32, 12, 111, 69, -34, -94, -39, -8, -86, -14, -106, 37, -29, 102, -20, -46, 89, 120, 46, -67, -40, 88, 91, 102, 125, -45, 115, -97, -96, -22, 115, -109, 1, 112, 78, -116, -35, -35, 61, 47, 10, 54, 52, 1, -16, 41, -14, 24, -16, -29, -99, 52, 74, 36, 122, 73, 1, 52, 68, -91, -78, -35, -47, -59, -119, 21, 126, -54, -39, 93, -63, 24, 42, -125, 0, 24, -33, -60, -20, -42, -63, 1, -5, 112, 15, 114, -51, 13, -64, -26, 24, -59, 69, -72, -44, -87, 91, 57, 29, 117, 14, 31, 89, -106, -81, -86, -15, 127, 33, 102, -65, 33, 9, 120, 114, 82, 123, 107, 120, -6, 54, -42, -103, -52, 80, -97, -77, -93, 78, -125, 115, -2, -93, 105, 1, -76, 57, -126, -98, 53, -114, 74, 70, 77, -18, 71, -23, -105, 27, -105, 107, -30, 78, -52, 82, -31, 76, -76, -29, 107, -31, 4, 51, 42, -78, 127, -66, -103, -11, -16, 78, -56, -5, -67, -79, 49, -93, -34, -112, 58, -106, -32, 127, 40, -125, -78, 109, -125, -99, -12, 43, 75, -53, 78, -96, 120, 17, 41, -24, 68, -117, 14, -16, 31, 40, -88, 127, 27, 68, -107, 17, -32, 100, -72, 68, -8, 92, -70, 23, 92, 68, 11, 23, 111, -52, 67, -42, 110, 40, 41, 0, 31, 50, -65, -79, 4, -94, 91, -98, -106, -86, -47, 12, 97, 121, 0, 35, -72, -116, 79, 122, -50, 105, -51, -1, 91, -38, -61, 80, 88, -126, -58, 27, -1, 1, -109, 113, 68, 62, -18, 29, -27, -56, -57, 123, 26, 107, -62, 26, -108, 87, 78, 74, -106, 76, -67, -119, 67, 47, 13, 20, 7, 26, 36, 51, 31, -62, 7, 8, 40, 75, 116, 61, -69, -103, -128, 65, 82, -87, -47, 105, -116, -68, -83, -9, -68, -32, 5, -68, -126, -72, 83, -10, 104, -23, -3, 37, 41, -36, -37, -56, -32, -52, 51, 89, -84, -15, 100, 16, -55, 92, -69, 51, 3, -87, 80, -42, 108, -93, -36, -87, 97, -68, 70, -2, -115, 101, 99, 12, 13, -10, 19, 61, 92, 6, -112, 77, -115, -29, -97, 15, 47, 19, 42, 121, -11, -89, -76, 24, -87, -87, 104, 59, 38, -87, -91, -20, 20, -46, 6, 46, 125, -42, -11, -50, 63, -73, -42, 21, -19, 7, -56, -97, -86, -96, 68, 32, 46, 17, 19, 15, -119, -38, 81, 0, -8, -86, -69, -63, 46, -19, 2, -81, 93, 36, -104, 106, -28, -103, -38, 23, 37, 99, 114, 124, -113, 109, -84, 84, -7, 98, 89, 105, 57, -47, -63, -92, -123, -12, -97, -49, -28, 43, -122, -3, 81, -95, -120, 37, -69, 57, -39, 122, -87, 126, 102, -37, -25, 52, -66, 79, -90, -112, -19, -113, 86, 45, 121, 91, 52, -123, 49, 73, 21, -44, -65, -61, -123, -125, -5, 15, -105, -28, -23, -5, -100, -27, -78, 119, 22, 71, 29, 116, 42, -100, -8, -111, -115, -71, -44, 60, -15, -6, 124, 45, -79, -119, 21, 39, -12, 112, 80, -61, 42, -54, -81, 31, -13, 106, 15, -69, -111, -125, -49, 48, -37, -88, 49, 12, -58, -22, -25, -44, 45, 36, 25, 127, 107, -98, -93, 115, -10, 71, 88, 110, -41, -39, 104, -108, -126, 51, -56, 55, 126, -32, 116, -41, 68, 61, 100, -111, -60, -116, 26, -59, -79, 42, 75, 84, 12, 102, -82, -24, 13, 14, 31, 90, -40, 110, 29, 86, 101, -87, -122, 99, -75, -34, 85, 50, -61, -11, -125, 88, 25, -115, 93, 87, -117, 76, -110, -110, -88, -103, -115, -12, -104, 77, 121, -106, 11, 92, 10, -65, -125, -60, -52, -68, 72, 79, -125, 104, 126, -128, 82, -21, 3, -2, -106, 97, 16, 67, 15, 124, 91, -124, 88, -48, 99, -80, -84, 93, 44, 127, 84, 96, -66, 2, 75, 59, -104, 123, -32, -43, 109, 41, -89, -22, -123, 81, 61, -20, -5, -6, 106, 61, -97, -11, -1, 55, 30, 60, 94, 35, -127, -101, -91, -45 );
    signal scenario_output : scenario_type :=( 127, 127, -128, 127, 127, 127, 42, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 8, 127, 127, -128, -128, 127, -128, 116, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -92, 127, 127, -63, 127, -128, -128, 127, 127, -128, -128, 127, 102, 127, -128, -128, -128, 127, 127, -128, 127, 23, -128, -128, 127, 127, -128, -128, 127, -128, -42, 11, 127, -128, -128, -24, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -103, -128, 127, 127, -128, -128, 127, -78, -128, 127, 127, -101, -128, -79, 127, -73, -128, -38, -128, -128, 127, -128, 127, 86, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 6, -128, 127, 127, -128, -68, 127, -128, -111, 106, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 53, 127, -128, 127, 127, 127, -128, 127, 127, -128, 50, 127, -128, 127, 127, -128, -128, -128, 127, -69, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -78, 59, 113, -128, 127, -128, -128, -128, 113, 15, 127, -128, -128, -128, 127, -128, 127, -128, 49, -128, 127, -128, 127, 127, -128, -128, 127, 55, -128, 127, 127, -74, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 2, -128, -128, 127, 127, 127, -128, -64, -128, 127, 127, 127, 127, -128, 23, -128, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -45, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -81, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 15, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 13, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 69, 127, -128, -128, 127, 127, -128, 127, 127, -128, 23, -128, 127, -128, 127, 127, -50, -128, -128, 127, 127, -128, -128, 127, -128, 127, -15, -80, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -42, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -32, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, -73, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 88, -54, -128, -128, 127, 127, -128, 95, -69, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -44, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 65, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 112, -128, 107, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 2, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -18, -96, -128, -128, 127, -81, -128, 127, -27, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 24, 127, 18, -128, 127, -128, 127, -128, 18, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -123, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 106, 127, 127, -128, -128, 127, 127, -128, -128, 75, 127, 127, 127, -128, -128, 127, -47, -128, -128, 127, 127, 127, -128, -128, 127, 127, -122, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -109, -128, -128, 127, 101, -114, 127, -128, 117, -128, 127, -128, 127, 127, -38, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, -114, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -54, 127, 34, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -118, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 24, -128, 127, 68, -128, -128, -128, -128, 127, -128, -128, -96, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 28, 127, -128, 127, 127, -128, -128, -128, 127, 127, -12, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -75, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 69, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 101, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 50, -128, 127, 127, -85, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 57, -128, 127, 127, -128, 73, 127, -128, -53, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 111, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -103, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -97, 127, -128, 106, 95, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -66, -128, 127, 127, -128, -128, -128, 6, 127, 127, 127, -128, -28, 127, 127, -128, 127, 127, -128, 122, 127, 63, -128, 127, -128, -17, 127, 101, -128, -128, -88, -81, 127, 119, 127, -128, -128, 127, 127, -128, 74, 127, -128, -128, -128, 127, 127, 127, -128, -128, 39, -128, 127, 127, 127, -128, -128, 5, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 76, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -68, 127, -10, 88, -128, 96, 127, 127, -128, 127, -43, -128, -128, 127, 127, -64, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -87, 21, 127, -128, 127, 0, 127, 127, -128, -128, -128, 127, -88, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 117, -128, 127, 127, -128, 127, -128, 127, 122, 127, -128, 127, -128, 44, 127, 64, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -43, -128, -128, 127, -128, 66, 127, -128, 36, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -3, 127, 127, -128, -48, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -112, -128, 127, 127, -13, -128, -75, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 59, -128, -128, -36, 127, -12, 127, -128, 93, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 90, -128, 127, -128, 127, -128, -128, -128, -12, 127, 127, 127, -128, 127, -128, -128, -128, 2, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -6, 127, 127, -128, -128, 127, 127, -128, -128, 111, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, -29, -52, -128, 127, -128, -128, 107, 127, 127, -128, -47, 127, -21, -128, -128, -128, 127, 127, -128, 127, -128, -128, 27, 127, 127, 127, -18, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 90, 127, -128, -128, 127, -128, -1, 81, 86, 127, 127, -39, -37, -128, -128, 123, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -91, -128, 127, 127, 127, -128, 111, 127, -128, -128, -37, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 92, 0, -128, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 3, 127, 127, 127, 34, -128, -128, -128, -128, 86, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -47, 127, 127, -128, -128, 58, 127, 127, -128, 127, 127, 68, -128, 127, -128, 127, -128, 127, -128, 29, 127, -128, -128, 127, 127, -128, -128, 127, -123, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 95, 127, -128, -128, 127, -73, -128, 127, 127, -128, -128, 127, 127, 103, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 73, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -49, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -98, 127, -128, 127, 96, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -18, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -71, -128, 127, 127, -128, -128, 127, -128, 81, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -44, -128, 127, 127, 127, 11, 127, -102, -128, -16, 127, 127, -128, -128, 127, 127, -50, -128, 127, -128, -128, 127, 127, -128, -128, 127, 96, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, 106, 127, 127, 127, -128, -128, -128, 127, 127, 88, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 116, 127, 127, -128, -8, -128, 96, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -6, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -23, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 96, -128, 127, 113, -128, -111, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 87, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -73, 86, -128, -128, 127, 127, -128, -128, -128, 127, 37, -128, 127, 127, -128, -128, 127, 127, 127, 108, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 117, -128, 127, 127, 127, 127, -128, -128, 127, 127, 91, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 86, 127, 123, -128, 127, 127, -128, -128, 127, -128, -108, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 0, 127, -128, 127, -34, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 52, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 29, -18, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -10, -128, -128, 127, 127, -128, -128, 127, 127, 16, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 0, 127, -128, -128, 127, -128, 127, -128, -79, 127, -116, 127, -128, -128, -128, 127, 127, -128, 127, 127, 109, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 112, -128, -34, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 98, -29, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -87, 127, -81, -128, 76, 127, 127, -128, 127, -128, 127, 127, -128, -128, -93, -31, 127, 127, 127, -128, 13, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -8, 91, 60, 127, 127, -128, -128, 127, -128, -128, 127, -71, -128, -128, 127, 5, -128, 127, -128, -128, 127, 122, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 48, 127, -8, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 76, 127, -128, 127, 127, -128, 127, 127, 11, -128, 127, -128, -128, 44, 85, -128, 127, 127, 127, -128, -128, 127, -7, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -47, 127, -128, 63, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -33, -128, 127, -128, 127, -128, 127, -128, 127, -128, 26, -128, -16, 127, -98, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 8, -128, -128, 124, 127, -128, 127, 79, -128, -128, 127, -128, -128, -128, 121, 127, 127, -128, -128, 127, 127, 127, -128, -128, 124, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -11, 127, -128, 127, -128, -128, -3, 127, 127, -128, -8, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 8, -128, 127, 127, -128, -128, -128, 127, 127, 127, 17, -128, -128, 57, 127, 127, -128, 127, -27, 127, -119, -128, -128, 127, 17, 127, -128, -128, -128, 127, -128, 127, 127, 1, -128, -128, -128, 127, -13, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -88, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -85, 127, 63, 127, -128, -128, 71, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 37, -128, -6, 127, 65, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 57, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 43, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 76, -128, -128, -24, -128, 127, 127, -88, -128, 127, -128, 127, 127, -128, 127, 127, 73, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 22, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 118, -128, 127, -128, -128, -114, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -122, 127, -128, -128, 127, 127, -128, 127, 127, -128, 70, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 118, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -86, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, 81, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -6, 127, 127, -128, -76, -128, 127, -128, 111, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 85, -128, 127, -22, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 22, -128, 127, 127, 127, -128, -128, -128, -38, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 93, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -45, 127, -128, -128, 3, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -80, 127, 127, -128, -128, -128, 127, 127, 127, -128, 54, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 47, -128, -58, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 29, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 87, -7, 127, 0, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 32, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 39, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -93, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 87, 127, 108, 95, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -33, 127, -75, -6, -128, 127, 127, -128, 127, 127, 6, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -106, 127, -71, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -54, -128, -128, 127, 127, 127, -128, 127, 127, -27, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -23, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -122, -128, 127, 127, 127, 49, -128, -128, 97, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -114, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -27, -44, 127, -128, -128, 127, 127, -128, 127, -75, -128, 127, 127, -128, 66, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 121, -128, 127, 127, -128, -128, 127, 127, -57, 127, -128, -128, 127, 127, -128, -128, -1, 127, -43, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -102, -128, 57, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -26, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -116, -128, 127, 127, 127, -86, -128, 39, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -93, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -71, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, -128, 127, -5, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -54, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -97, 65, 127, -98, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 69, -128, 127, -128, 127, -128, 127, -53, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -45, -86, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -29, -128, -128, 127, 52, 127, -128, -128, 127, 127, 127, 127, -128, -128, -17, 127, 127, -128, 117, 127, -128, 127, 127, -128, -128, 127, 127, 127, 107, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 124, -26, 122, 33, -128, 127, 13, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -109, -128, -128, 127, 127, -54, -128, 127, -128, -128, 8, 127, 127, -128, -128, 73, 127, -128, -128, -128, 127, 127, 127, -128, -128, -63, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -100, -128, 3, 127, -63, 127, 12, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 107, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -101, 127, -128, 127, 127, -45, 127, -128, -128, 127, 127, 29, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -66, 18, -128, 127, -100, -128, 127, -128, -90, -128, -112, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -58, -124, 127, -128, -128, 127, -57, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -37, -128, 127, 127, -42, 127, -128, -128, 127, 127, -128, 127, 17, -106, -128, 127, 127, -128, -128, -128, -128, 52, 127, -128, -128, 127, 127, -128, -128, 127, 12, -128, -128, 127, -128, 127, -128, -128, 127, -22, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 65, 127, 18, 127, 127, -128, -128, 127, 127, -85, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -53, 124, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -18, -128, 127, 127, -128, -128, 127, 127, -92, -128, -128, 127, -128, 16, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -96, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -97, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 98, -128, -128, 127, -128, -128, -128, 127, -128, -112, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 24, 66, 127, -128, -128, -128, 127, -85, 96, 75, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -18, -128, 81, 127, 127, -128, 127, -128, 127, 127, -49, -128, -128, 127, -128, -128, 127, -128, 127, 127, 127, -128, 63, 127, 127, -128, -87, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, -119, 127, -92, -128, 127, -128, -128, 127, 127, 127, -63, -128, -128, -128, 127, -65, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 103, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 91, -128, 127, -128, 127, -128, -128, 127, 127, 127, 2, -103, -106, -52, -128, 127, 45, -128, 127, -85, -128, 127, -111, -128, 127, -80, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -111, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -87, 127, 127, -128, 127, -128, 66, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 37, -128, 127, 127, 127, -128, -128, 127, 127, -128, 16, 127, 127, -80, -128, -128, 127, 127, -128, -80, 127, 127, -128, 33, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 23, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -118, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 102, -128, 127, -128, 127, 127, -128, -128, -22, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -73, -128, -60, -128, 127, 54, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, 39, -128, -128, -63, 127, -114, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, 117, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -68, -128, 127, -128, -128, -31, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 18, 127, 127, -128, -128, -85, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 116, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 3, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -43, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, -58, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -81, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -80, 101, 127, -128, -128, 127, -128, -128, 57, 127, -128, -128, -128, -128, 127, 127, -128, -26, 22, -128, 127, -102, -128, 127, 127, -128, -128, 127, 127, -128, -128, 108, 127, 127, -128, -27, 127, 127, 127, 93, -128, 127, -128, 127, -128, -58, 127, 127, -128, -128, 65, 127, -128, 122, -128, 127, -128, 127, -128, -128, 127, 121, -128, -102, -128, 127, 127, -96, 127, -128, 127, -128, 127, -31, 80, -128, 127, -27, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -64, -128, -128, 127, -128, -128, 5, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -50, -43, -128, 127, 127, -128, 127, 127, -128, 3, 127, 127, 127, 127, -128, -128, -128, 127, 127, 54, 127, 127, -128, -128, 127, 127, -128, 127, 85, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -98, 127, 127, -112, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 123, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 68, 127, -128, -128, 127, 127, 118, -128, -128, 127, -102, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -109, 122, 127, -128, 39, -128, 55, 127, 127, -128, -122, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 5, 127, 127, -128, 127, 127, -128, -128, 127, 127, 47, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -121, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 55, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 18, 127, -128, 29, 127, -128, -128, 127, 127, -128, -128, -128, 66, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -12, -128, 127, -97, -128, 127, 127, 127, -128, -128, 127, -10, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 117, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -100, -128, 127, 127, 127, 127, -128, 74, -128, 127, -128, -128, 127, -128, 127, -80, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 79, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 44, 127, -128, 127, 127, 127, -128, 127, 98, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 102, 127, -128, -128, 127, 127, -128, 127, 18, 127, 127, 127, -128, -8, 27, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 66, -128, 127, -128, 127, 127, 5, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 55, -128, -128, 127, -128, -128, 127, 127, -128, 127, -106, -128, -128, 127, 127, -13, -128, -128, -128, 127, 127, -128, -128, 127, -128, -58, 127, -128, -128, 127, -128, 127, -128, 127, 127, 28, 127, -128, 23, -128, -128, -43, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 102, 127, 127, -128, 127, 127, -128, -128, 1, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 54, -128, -128, 127, -128, 127, 80, -128, -128, 127, -23, -17, -128, 127, 127, -128, -128, -128, 127, -128, -92, -128, 127, -128, -128, 127, 127, 127, -128, -24, -128, 127, 45, -128, 127, -128, 127, 127, -128, -128, -33, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -91, 127, 127, -128, -128, 127, 127, -128, -49, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -101, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -45, -128, 127, -128, -128, -81, 42, 127, -128, 101, -128, 127, 107, -128, 127, -113, 127, -128, 127, -128, 127, 127, 127, -113, -128, -128, 127, -128, -7, 127, -128, 127, 127, 127, -85, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -53, -64, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 0, 127, -128, -128, -128, 127, 106, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, 127, -3, -128, -58, -128, 127, -128, -128, 127, 127, 127, 60, -128, -103, 127, 127, -128, 127, 127, -128, -128, -76, 127, 127, -128, 127, 74, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -79, 127, -128, 127, 127, 42, -128, -128, -128, -128, 127, -128, -80, 127, 127, -128, -52, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -39, 127, 127, -128, -128, 127, 43, -128, 127, 127, -128, -128, -128, 127, -128, 127, -39, 127, 36, 127, -128, -128, -63, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -123, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -93, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 29, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -39, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -59, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -122, 127, -128, -7, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 66, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -48, -128, 127, -128, -55, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -11, 127, -128, -128, 54, -128, 127, 127, -128, -128, -128, -80, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -85, 127, -118, -128, 71, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 45, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -17, 127, -128, 127, 121, 127, -128, 127, -87, 117, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 58, 127, -95, 127, 127, 127, -128, -98, -128, -128, 28, 127, 81, -128, 127, -128, -128, -11, 127, 127, 117, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -88, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -36, 127, 127, 127, 102, -128, -128, -128, 127, 127, -128, -128, 114, 127, 127, 127, -128, -128, -128, 127, 127, 127, -44, -128, -128, -128, 127, 127, 127, -128, -54, 127, -128, -128, 127, 127, -106, -128, 44, -128, -66, -128, 127, 127, -128, -128, -116, 127, 127, 127, -128, -128, -128, 31, 127, 127, -119, -128, -128, 127, 127, 97, 127, -128, 127, 127, -11, -128, 127, 127, -128, -128, -8, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -101, -128, -128, 127, 127, -128, -128, 63, -128, 127, 127, -128, -128, 127, -128, 127, -128, -27, 127, 127, -128, -128, -128, 127, 127, 66, -128, 127, 127, 127, -128, -128, 127, -128, -107, -128, 127, 27, -39, -42, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 17, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 64, -128, 127, 127, 127, -128, -128, 127, -38, 36, -128, 127, -36, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -38, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 23, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 80, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -33, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 113, -8, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 37, 127, -128, -128, -128, 127, -128, 127, -128, 127, 33, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 111, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -124, -128, 127, -128, 127, 127, -75, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 73, 127, 127, 113, 95, -128, -128, -128, 127, -78, -48, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -6, -128, 127, -128, -128, 127, 42, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 57, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -73, -75, 127, -128, -90, 127, 127, -128, -128, -78, 127, 127, -128, -128, 127, 127, -128, -128, 79, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 22, -128, 127, 117, -128, -128, 127, 127, -47, -128, -128, 127, 127, -68, -128, 127, -128, -50, 127, -128, -128, 52, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, -54, 127, 127, -128, -128, 127, -128, -128, 53, 127, -128, -128, -128, 127, 127, 102, -128, -128, -23, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -96, 127, -128, 43, -128, -128, -128, 127, -128, 127, -15, 127, -128, 127, -128, -7, 118, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 101, 127, 127, 98, 127, -128, -128, 127, 127, 127, -74, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, 127, -117, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -76, -128, -33, 127, -128, -128, 127, 127, -50, -128, 127, 127, -128, 16, -128, -128, 127, 127, -128, 48, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -64, 127, -128, -128, 127, -128, -121, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 59, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -48, 127, 57, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -54, -128, -128, -124, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 63, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -3, -128, -128, 127, 127, -128, -128, 127, 127, 127, -122, -128, -128, 127, 47, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 102, 127, 29, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 70, 127, -128, -128, 127, 127, 127, -101, -128, -128, -128, 127, 127, -128, -128, 103, 127, -128, 127, 127, -128, -28, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 17, 127, 109, -128, -128, 127, 127, -128, 127, 112, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -96, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, 102, 127, -128, -128, 127, 127, -128, 127, -128, 2, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 21, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 5, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -114, -128, 127, 127, 127, -128, -47, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 106, -128, 18, 127, 127, -128, -128, 127, 127, -107, -128, -128, 127, 127, -128, -22, 127, -68, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -86, -128, -128, 127, -128, 127, -128, 127, 127, -128, 109, -128, 127, -58, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -101, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 24, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -108, 127, -128, 127, -128, -128, 127, -128, -128, 52, 127, -128, 127, -92, -128, 127, 127, -128, -128, 127, 52, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -123, -128, 127, 127, -128, -128, 21, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 52, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 71, -128, 127, -43, -128, -128, 127, 127, -128, -128, 127, 127, 44, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 81, 127, -128, 29, -128, 127, 127, -128, -128, -49, -114, 127, -128, -128, -128, 127, 127, -128, -128, 127, -81, -128, 127, 127, -128, -128, -17, 127, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, 103, -128, -128, 108, -128, -128, 127, -108, 127, -128, -128, 127, -128, -58, 127, 127, -128, 98, 127, -128, -128, 90, -128, 127, 127, -128, -128, 127, 127, 90, -128, -128, -128, -124, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -42, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 91, -128, 47, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -76, -128, 127, 127, -128, -90, 127, 127, -128, 127, -127, -128, -57, 127, 127, -128, 112, 127, -128, 98, -78, 5, 127, -93, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 97, -128, -128, 127, -100, -128, 127, -128, 114, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -13, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, 127, -71, -128, -3, 127, -119, 80, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -69, -128, -128, 127, -128, -128, 127, 17, 10, -128, 127, -128, -128, -128, 127, 127, -128, -128, -60, 57, -128, 127, -128, -128, 127, 60, -128, 127, 127, -128, -128, 17, 127, -23, -85, 38, -128, -128, -128, 127, 31, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -71, -128, 127, 103, 127, -128, 127, -128, 127, -128, -54, 127, 127, -128, -128, 127, 127, -128, 127, -128, 78, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -42, 127, 127, -128, 69, 127, 75, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -50, 127, -128, 127, 127, 127, -128, 42, -128, 127, 127, -128, 123, 127, -128, -128, -128, 90, 127, -96, 127, 127, -128, -128, 127, 127, -128, -128, -95, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, 49, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, -92, -128, -128, 127, 127, -128, -128, -128, 116, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -21, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, 60, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -103, -128, 127, -128, 127, 127, 18, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 22, -78, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -52, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 12, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -31, 127, 127, -128, -128, -128, -128, 127, -128, 127, 127, -128, -128, 10, -128, -128, 127, -42, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, 98, -128, -128, -69, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 64, -128, 127, 127, -5, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 81, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -121, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -97, 127, -128, -128, -128, 127, -50, -128, -128, 31, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 0, 127, -128, 73, -128, 127, -128, 127, -128, 7, 58, 119, -128, 109, -128, -128, 127, 127, -128, -128, 127, -63, -128, 108, 127, -106, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 75, -3, 127, -128, 127, 127, 59, -128, 127, 127, 127, -128, -128, -13, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -117, 127, -128, 113, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 58, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -79, 108, 127, -26, -128, -128, 127, 127, -128, 127, 127, -128, -128, 97, 127, -128, -128, -16, 26, 127, -54, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 49, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -66, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -10, -55, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 116, -109, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 0, -128, -43, 127, -11, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 0, 90, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 118, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 27, -128, 127, 127, -128, -128, 127, -98, 118, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 2, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 119, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 60, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -76, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 69, -128, -128, 127, 127, 127, 32, -128, 119, 127, -128, 127, 127, -80, 127, 17, -128, 127, 127, -128, -128, -128, -128, 127, 127, -36, 127, -128, -128, -128, 127, -34, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 76, 127, 42, 127, -128, -102, 127, 127, -128, 127, -128, -15, 113, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 26, -128, 127, 127, -128, -128, 127, 127, -128, -75, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 64, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -108, 127, -128, 127, -128, -128, 127, 127, -12, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 112, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 80, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -57, -128, 92, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -117, 127, -128, -128, -55, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 71, -128, 11, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 52, -128, 127, -128, -128, 127, -128, 71, 127, 127, -128, 127, -128, 81, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -116, -128, 127, -128, -128, -128, 127, 114, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 43, 127, 127, 127, -128, 114, -22, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -39, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 42, -6, 127, -122, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 70, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -34, 127, -128, -128, -54, 127, 127, -128, -128, -128, 127, 127, -96, -128, -128, -128, -128, 127, -118, 127, -128, -128, -128, 127, 6, -128, 127, -128, -128, 127, 127, -68, 127, -128, -13, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -1, -128, 127, 127, -128, -111, 119, -128, 127, 127, -128, -128, 127, 127, 127, -88, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -18, 127, -128, -128, 127, 127, -128, -128, 127, -128, 68, 127, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, -117, -128, 127, -128, 127, 127, -128, 127, 127, -128, 57, -128, -128, 127, -128, -128, -128, 127, -128, 127, 29, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -69, 127, 127, -128, 42, 127, 127, 127, -128, -29, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 22, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -96, -128, -92, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -8, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -114, -128, 127, -128, -128, -28, 127, -113, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 107, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -28, -128, 127, -128, 127, 127, -128, -128, 127, 127, -117, -128, -128, -128, 127, 127, -17, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -23, 127, -73, 127, 71, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, 95, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 17, 28, 127, -107, -128, 127, 127, -128, -92, 116, 127, 127, -128, -116, 127, -128, 127, 127, 127, -128, -128, -107, 127, 7, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -54, -128, 127, 127, 127, -128, -128, -128, 127, -33, 127, -18, -128, 127, 127, 127, -128, -128, -58, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -101, 127, -95, 127, 127, -128, -121, -98, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, -80, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -90, 127, -128, -118, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -101, -128, -128, 127, 127, -106, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -32, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 118, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 0, 127, 90, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -24, -128, 127, -128, 127, -128, 127, -128, 127, 127, 112, -128, 127, -128, -128, -22, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 5, -128, 111, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 38, 127, -128, 127, 127, -128, -128, 127, -128, 43, 127, -128, 127, -128, 127, 117, 127, 11, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, 26, -80, -128, -128, 127, 127, 86, -128, 103, 127, -128, -128, 127, -87, -128, 127, -128, 127, -124, -128, -128, -123, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 76, -50, -128, -128, 127, 127, -128, -79, 127, -128, -128, 127, -128, -128, -128, 127, 108, 127, -128, 127, -128, -128, 69, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 0, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -109, -128, -128, 124, 127, -128, -128, 127, 127, -128, 98, 29, -128, -128, 127, -100, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 49, -117, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -106, -128, -64, -128, 0, 127, -101, -128, 127, -60, 127, -128, -28, -128, 127, -49, -128, -10, -128, 127, 127, -36, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -102, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, 63, -128, 127, -128, 73, 127, 127, -106, 127, -128, -128, 127, 127, 127, -128, -100, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -13, 42, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 102, 127, -128, 127, -128, 127, -128, 127, 73, 127, -124, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -3, -128, 127, 127, 127, -128, -128, -128, 121, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 59, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -73, -128, 127, -128, -128, -128, 127, -128, 127, -128, 26, -128, 127, -128, -128, -128, 127, -128, 127, -22, -128, 127, 47, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 59, 127, 127, -128, 127, -128, -128, 96, 127, -128, -66, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -18, 127, 127, 127, -128, -128, 127, -128, 127, 127, 74, -128, 127, -128, 53, -128, -128, 127, 127, -128, -128, 127, 127, -23, -128, -128, -128, 127, 127, -128, -128, 127, 127, 34, -128, -128, 127, 127, -128, -70, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 15, -128, 127, 127, -128, -128, -128, -128, 111, 127, 127, 23, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 78, 127, -128, 127, 127, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -109, 127, -128, -128, -128, 127, 127, 101, 91, 127, -116, -128, 127, -128, 127, 127, -128, -128, 127, -128, -103, -128, 127, 127, -128, -128, -79, 127, 127, 127, -128, -128, 127, -128, -128, 127, -11, -98, -128, -128, -10, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -88, 127, -128, 127, 127, 102, -128, 127, -128, -128, 127, 127, -128, -128, 42, 127, 127, -119, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 32, -128, 127, 24, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -63, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 121, -128, -128, 127, -128, 127, -23, -128, -128, 127, 118, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 2, -128, -47, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -42, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, -21, -128, 93, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -65, 127, -128, -121, 127, 127, 127, -128, -128, 127, 127, 80, 127, -95, -128, 127, -128, 127, -128, 127, 127, 36, -128, -128, 127, 127, -128, -128, -128, 32, -128, 111, 127, -128, -10, 127, -128, -128, 15, 127, -128, 127, 127, -128, -128, -128, -59, 127, 121, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 5, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 11, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -90, 127, -128, -128, 127, -92, -128, 127, 127, -128, -128, 32, 127, -128, -128, -128, 127, -128, -128, 127, -66, 127, -128, -128, -128, 127, 127, -128, 127, 73, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 101, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 112, 44, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -52, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 23, 7, -128, -8, 127, -128, -55, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -116, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -48, 127, 127, -128, -128, -34, 127, -127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -44, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -22, 127, -128, -128, 127, 127, -87, 127, -128, -102, -128, 127, 127, 127, 127, -128, -128, 102, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 7, 76, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 32, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -12, -128, -128, 127, 127, -128, 127, 127, -128, -87, 127, -128, -128, 127, 127, 127, 127, -128, -128, -21, 127, -128, 48, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 58, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -79, -128, -128, 79, 127, -128, 127, -128, -128, -128, 127, 127, -128, -97, 127, -128, 127, 127, 127, -128, 88, -128, 127, 127, 60, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -96, -128, 127, -128, 88, 26, 127, -128, -128, 127, -128, -128, 81, 127, -128, -128, 127, -28, 127, -128, -128, -128, -128, 103, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -122, 127, -128, -58, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 29, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 124, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 70, 127, -128, -44, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -3, 127, -128, 127, 127, 78, -59, -128, -128, 127, -128, -128, 127, -128, -128, 127, 107, 127, 76, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -111, -128, 108, 127, -103, -128, -128, 127, 127, 127, -128, -128, 48, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 76, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -64, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -87, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 111, 109, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, -128, 111, -128, 78, -128, -128, 127, 127, -128, -128, -128, 127, -128, -80, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -6, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -38, 127, 1, -128, -128, 127, 127, -128, 127, -128, 127, -128, -124, 43, 127, 127, -128, 127, -128, -93, -128, 127, -128, -128, -65, 127, -54, -128, 49, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -65, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -92, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 13, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -39, -100, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 79, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -87, 127, -32, -128, 127, -128, -73, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -66, 75, 127, -128, -128, 127, -128, -128, 127, -11, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -80, -128, 127, 76, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 113, -128, 127, -128, 127, -128, 127, -128, 127, -78, -128, -128, 127, 102, -128, 127, -128, -128, 127, -128, -128, -75, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -122, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 10, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -119, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 97, 127, -128, -128, -39, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -34, -128, -128, 127, 71, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -16, 127, -128, -128, 38, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 118, 127, -128, -128, 127, -12, -128, 127, 127, 127, -128, -98, -128, -128, 127, 127, -128, -128, 127, -113, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 29, -128, -128, -128, 64, 127, 127, -128, 117, -128, -118, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 27, -128, 39, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 28, -65, 127, 127, 127, -128, -128, 127, 127, -95, -128, 127, -128, 127, 127, -128, -128, -128, 127, -52, 26, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 69, 127, 127, -96, -128, -128, 112, 127, -128, 127, -128, 127, -128, -128, 127, -128, -128, -128, -80, 127, 127, -128, -128, -128, -128, 116, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 60, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, 55, -128, 127, 127, -128, 127, -93, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -107, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 59, -128, -128, 127, 127, 127, 127, -128, -128, -50, 127, 127, 127, -128, -128, 127, 127, -128, 127, 109, 39, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -117, 127, -128, -128, 127, 47, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -36, 127, -128, -128, 127, -128, -128, 127, 53, -43, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 98, 127, -128, 127, 127, -128, -128, -128, 127, 127, 60, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 39, 44, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -106, 127, -113, -128, -59, 127, -128, -128, -114, 127, 127, -128, -128, 127, -128, -128, -107, 127, 127, -128, -128, 127, 127, -128, -128, 127, 70, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -69, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -80, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 22, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 81, 127, -128, -128, 127, 0, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -108, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 39, 127, -128, -128, 98, 127, -128, -128, 127, 127, -128, -128, 64, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -87, 127, 127, -128, 127, -128, 127, 127, 127, -6, -128, -128, -128, 127, 127, -128, -128, 54, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 106, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -44, 127, -128, 127, 127, 127, -128, -119, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -57, 127, -128, -128, 127, 127, 127, -128, 121, 127, 18, -128, -128, 127, 127, -128, -128, 127, 127, -128, 1, -122, -128, 127, 127, 127, -128, -128, 127, 127, -128, -31, 50, 127, 127, -128, -128, -128, 127, 127, 118, -128, -128, 127, 127, -128, -128, -28, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, -106, -13, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -109, 45, 127, 127, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 32, 127, -128, 127, 127, -128, 118, 127, -128, -128, 127, 127, -128, 127, 127, -119, -128, -65, -128, 127, 127, 127, -128, 2, 127, -128, -128, 127, 127, -128, -128, 109, 127, -128, -79, 127, -128, 127, 127, -128, -128, 127, 127, 127, 79, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, -128, -128, 113, 127, 122, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 23, -128, -128, 127, 127, 48, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -85, 127, 127, -128, 127, -31, -53, 127, -128, 127, 127, -128, 59, 127, -96, -128, -122, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, 127, 60, -128, 127, 127, -128, -128, 127, 127, -107, -128, 65, 127, -128, -128, -128, 22, 111, 127, -128, -128, 127, 127, -128, -128, -68, -12, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -50, 127, 127, -128, 127, 127, -22, 127, 127, -128, 100, 127, -96, -13, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 7, 86, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 36, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -101, -128, 127, -128, -128, -128, 127, 45, 127, 127, -128, 109, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 32, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -114, -128, -78, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 113, -128, 3, -128, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -92, 127, -128, 90, -128, 127, 127, 127, -128, 63, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 93, -68, 127, -128, -128, 127, 127, -128, -128, -18, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 36, -127, 127, -17, -128, 47, -128, -128, 127, -128, -70, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 13, -128, 127, 127, 127, -128, -128, 127, 127, -128, -122, 127, 127, -128, -128, 127, 127, -128, 16, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 100, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -97, 127, 127, -128, -128, 127, -88, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 55, -128, -128, 36, 127, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, -112, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, -53, 127, -36, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -57, 127, 127, -128, -128, -128, -22, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 90, -128, 127, -128, 23, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, -111, 127, 127, -128, -23, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 27, 127, 127, -128, 127, -128, -128, -11, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -124, -128, -128, 127, -75, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -102, 127, -128, -128, -70, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 66, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -86, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -93, 109, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -22, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 27, 127, -128, 127, -23, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 39, -128, 127, -128, -128, -128, 127, -75, -128, 127, 127, -128, -128, 127, -128, 79, 127, 123, -128, -128, 127, -36, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -118, 127, 127, -128, -128, 127, -27, 127, 127, 16, -128, -128, 127, 127, -71, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 10, -128, -55, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -90, 127, -128, -128, 39, 32, -128, 127, -128, 127, 127, 68, -128, -128, 127, 49, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -8, 127, 127, -128, -128, 114, 127, -128, -64, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -50, 127, 127, -128, -128, 127, 55, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 95, -128, -128, -128, 127, 127, -128, 127, -128, 127, -93, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 0, -128, -128, 127, -128, -119, -128, 127, -128, 127, 80, -128, -63, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 3, 127, 71, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 55, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -97, 127, 85, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -111, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 28, -17, 127, -128, 101, 127, 127, -86, -128, 127, -128, 18, 127, 127, -128, -128, 127, 127, -128, -58, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 8, -128, 127, -128, -128, 3, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, -26, 55, -101, 79, 127, 127, -128, 6, -128, 127, 127, -128, -128, 127, -93, 127, -73, -128, 127, 127, -128, -128, -128, -128, 17, 127, -128, -128, 127, -128, -128, 127, 127, -128, 26, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 87, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 17, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 38, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 57, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 28, -128, 127, 127, -128, -128, -118, 127, 29, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 91, 127, -22, 127, -128, -128, -128, 127, 80, 127, -128, 127, 127, -128, 78, -128, 127, 127, 117, -128, -128, 127, 127, 127, 81, 127, -128, -128, 127, -73, 127, -128, -128, 79, -128, -128, 127, 127, 127, -128, -128, -128, 127, 107, -128, 127, 58, -128, -128, 127, 127, 127, -128, 127, 127, -128, -91, 127, 127, -128, -39, -128, -13, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 44, 127, -128, 127, 12, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 37, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 2, 127, -128, -128, 0, 127, 8, -128, 127, -63, -128, -128, 127, 127, 28, -128, 127, -128, 127, -128, -128, -128, 127, 23, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 54, -128, 127, -128, -128, -128, 127, -87, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -53, -33, 127, -128, 76, 127, 127, -128, 127, -128, -59, 127, -128, -128, 127, -116, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, -128, -60, 127, 44, -128, -128, 127, 127, -128, -128, -12, -128, 127, 127, -128, -128, 127, 8, 127, -128, 47, -70, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 43, 127, -128, -128, 127, 43, 127, 127, -128, -128, 127, 109, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 86, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 42, 127, 127, -128, -128, 127, 127, -128, -128, -17, 118, 127, -128, 127, 127, -128, -128, 31, -128, 127, 127, -128, -128, 103, 127, -28, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -116, -118, 127, 127, -128, -128, 127, 127, 127, 127, -119, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 124, 127, 127, -128, 127, 57, 24, 127, -128, -128, 127, 127, -128, -128, 127, -128, 34, 127, 127, -128, -128, -128, 116, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -95, 127, 127, -44, -128, -128, 127, 127, -128, -128, 127, 113, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 93, -128, 127, 127, -128, -45, -128, 127, 127, 127, -128, 90, -128, -44, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 38, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, -128, -8, 127, -128, -128, 54, 127, -128, 127, -16, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, 64, -128, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -24, 127, 127, -128, 127, -128, 34, 127, 127, -128, 127, -128, 127, -87, 127, -128, -128, 127, 127, 127, 127, 65, -128, -12, 127, 127, -128, -128, 85, 127, 127, 127, -128, -128, 127, 127, 69, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 0, -128, 127, 127, 127, -128, 127, 10, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 106, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 8, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 33, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 98, 127, 127, -128, -119, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -13, -8, 127, -128, 127, -128, -112, -128, 54, 127, -36, 127, 60, -106, -128, -128, 127, 127, -36, -128, -128, 127, 127, -128, -128, -128, -28, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -6, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -28, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 97, -17, -128, 127, 127, 13, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, -39, 127, 127, 127, -128, 0, -128, 127, -128, 127, -128, 127, 10, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 48, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -112, 127, 127, -128, -74, 127, -128, -128, 108, 127, 45, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -18, -91, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 91, -128, 57, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -16, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 103, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 28, 127, -128, -128, 127, 127, 57, -128, 127, 127, 127, -128, 0, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -103, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -85, -128, 127, 127, -128, -128, 127, -128, 127, -128, 73, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 1, -15, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, -96, -128, 127, 127, -128, -128, -128, 127, 127, 122, 127, -128, -106, -128, -128, 127, 127, 127, 92, -128, -128, -128, -128, 127, -128, 127, -97, 127, 48, -128, -128, -128, 7, 127, -128, -22, -85, -58, -128, 127, 127, -128, -128, 127, -128, 24, 127, 127, -85, -128, 10, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, -11, -128, -128, -70, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -95, -121, 127, -128, -128, 70, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -66, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -68, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -107, 127, -128, 127, -128, 116, -128, -100, 127, 127, -128, 127, 127, 127, -128, -29, 32, 127, -128, -128, 127, 127, -128, 34, 127, 127, -90, -128, -128, 127, 127, -128, -128, -28, -128, 127, -128, -128, 127, 127, -128, -128, 116, 127, 127, -128, 119, -128, 127, 127, 63, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 119, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -38, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 42, -101, 127, -128, 127, -128, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 112, 127, -128, 127, 127, -75, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 11, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, -39, -128, -128, 127, -128, -128, 127, -124, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -64, -117, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, 116, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, 28, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, 29, 127, 2, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 31, 127, -128, -128, -128, 127, 127, -112, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, -128, 60, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, 127, -70, -128, 127, -128, 127, -128, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -47, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 73, 127, 127, -128, 34, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -106, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, -48, 127, -128, -86, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 121, -128, 127, -128, -128, 127, -128, -38, -128, 127, -128, 127, -128, -128, 100, -128, -42, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -64, -128, -128, 127, 28, 127, -128, 3, -128, 96, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -60, 127, -128, -128, 127, 127, -128, -106, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, -74, -128, 127, 88, -128, -128, 127, 127, -128, -38, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -49, -128, 127, -128, 127, -128, 2, -128, -128, 43, 127, -128, -128, 127, 97, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -7, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, 127, -128, -128, 66, 127, 127, -128, -128, 78, -128, 127, 127, -128, -128, -71, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -98, 127, -128, -128, -128, 48, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 23, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -47, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 127, -124, -128, 127, 127, -128, -128, 127, -112, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 47, 127, 127, -128, -128, 127, 127, -128, 13, 127, -128, -128, -123, 3, 127, 127, -128, -128, -128, 127, -122, 127, -128, 2, -128, 127, -128, 103, -128, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, 127, 100, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -18, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 114, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -102, 127, -128, -112, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 22, -128, 127, 127, -128, -128, 127, -38, -128, 127, -128, -128, -128, 127, -128, -108, 127, 38, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -34, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 117, 127, -128, 8, 127, -128, -128, -128, -116, 127, 127, 127, -128, 116, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 16, 127, 64, -128, -128, 127, -128, -128, -128, -59, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, 55, 127, -128, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 95, -128, -128, 127, -128, 127, 127, -22, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -74, -128, -128, 127, 127, -128, -128, 127, -54, -128, 127, -128, -128, 127, 127, -128, 10, 47, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, -128, 127, -80, -117, -128, 127, -128, -31, 127, 127, -26, -128, -128, 127, 127, -128, 32, 127, 127, -128, 127, -128, 127, 127, -128, -128, 73, 127, 127, -128, 127, 6, 127, -93, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 52, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 28, -64, -128, 127, -128, -128, 127, 127, -128, -128, 59, 127, 127, -128, 33, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -13, 127, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 42, 127, -100, -95, -93, -128, -128, -128, 127, 111, 127, -101, -128, -128, 127, 127, 127, -106, -127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 78, 127, -128, 127, -128, -128, 127, -128, -128, -128, 127, -128, -117, -128, -128, 127, 127, -128, -128, -127, 127, -128, -128, 80, 127, 127, 127, -128, 127, 127, -128, -128, 50, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -88, 13, 127, -128, 127, 127, -17, -128, -128, 73, 127, -123, 127, 127, 127, -128, 39, 127, -128, -128, 127, 127, -128, 127, -128, 127, -108, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 100, -54, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 71, -12, -128, -128, 127, 79, -128, 127, 127, -128, -128, 127, 127, -128, -128, -27, 127, -128, 127, 127, -128, -80, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -45, 127, -128, -128, -128, 127, 127, -122, -128, 127, 127, -128, -128, 127, 127, -128, -128, 47, 127, 114, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, 114, -112, -128, -128, 127, 127, -53, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 27, 80, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, -70, -128, 127, -128, -128, 42, 127, -128, -128, 127, -128, 127, -128, 127, -52, -128, 6, -39, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 1, 44, 127, 127, -128, -128, -128, 127, -73, -128, 127, 127, 127, -128, -16, -128, -128, -128, 127, 127, -128, 127, -128, -123, -128, 127, 127, -128, -5, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 121, -128, 127, -128, -128, 127, 127, 5, -128, -128, 127, 127, -128, -128, -36, 127, 127, -128, -128, -128, 127, 98, 127, -128, 127, 96, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -23, 127, -31, -128, -55, 127, 127, -128, -29, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 54, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, -128, 0, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -59, -128, -128, -128, 127, 6, -128, 127, -93, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -74, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 28, -128, -128, -128, 127, 127, 127, 127, -128, -128, -75, 127, 127, -128, -128, 127, 127, -128, 127, 21, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, 64, 127, -48, -128, 127, -128, -128, 22, 127, 127, 45, -128, -128, 127, -1, 127, 15, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, -45, 127, 127, -128, 127, -128, -128, -75, 127, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, -15, -128, -93, 127, -128, -128, 127, 127, 127, -128, 127, 87, 127, -128, -128, 127, 127, -128, 50, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -63, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -55, 127, -128, 127, 98, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -100, -63, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, 127, 21, 127, -128, 80, -128, 127, -128, 127, -128, 127, -128, -16, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -113, -128, -128, 127, 127, 127, -128, -128, -128, 88, 100, 127, 127, 127, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 13, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 107, 127, -128, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 29, 127, -128, -128, -114, 127, 76, 13, -128, 127, 127, -128, 127, 7, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, 33, -128, 127, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 127, -34, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, 127, -7, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, 88, 127, -54, 127, -112, -128, 23, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 39, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 12, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 21, -128, -128, 127, -128, 86, -128, 127, -128, 127, -128, -128, 111, 127, 127, -128, -86, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 28, -128, -128, 127, 127, 127, -128, -128, 0, 127, -128, 127, -128, 127, -128, -128, 127, 93, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -12, 127, -128, -128, 111, 121, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 127, 55, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -43, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 108, -128, 3, -128, -52, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 69, -128, -128, 127, -128, 127, -128, 127, 127, 78, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, 92, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 53, 127, -128, -128, 127, 127, -48, -128, 127, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -28, 127, -128, -128, 127, 127, -121, -128, -81, 127, -128, 127, 127, 127, -128, -128, -128, 127, 0, -128, 127, 16, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, 0, 113, 127, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -58, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 109, 127, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -23, -128, -128, 127, -128, -128, 127, 127, 116, 76, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 60, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, -128, 124, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 63, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 74, 123, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, -128, -128, 127, -28, -128, 127, 59, 127, -128, -57, 127, 127, -128, -128, -128, 5, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -91, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 103, 127, -128, 127, -128, -128, -74, 127, -128, 127, -128, -128, -128, 127, 127, -128, -29, -128, -36, -128, 33, 127, -91, -128, 127, 127, -128, -128, 127, 29, -128, 127, -128, -128, 127, 127, -128, 127, -124, -128, 127, 127, -128, -128, 16, 127, 127, -91, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 79, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 68, -128, -128, 127, -128, 127, 127, 38, -128, -100, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 54, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, -128, 60, 127, 127, 17, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -101, 127, 127, 49, -128, -128, 127, -128, 69, 127, 76, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -47, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -27, -128, -128, 127, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -63, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, -58, -128, -95, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -24, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 11, -128, 127, 127, 127, -128, -128, -44, 127, 70, 127, -128, -128, 127, 127, -128, 127, -108, -12, -34, 127, 127, -128, -128, 127, 127, -128, 53, 127, -128, -128, 127, 127, -79, -128, 127, 127, -128, 127, -128, 127, -128, -128, -127, 127, -128, -78, 127, 127, -128, -128, 127, 127, -128, -34, 127, 121, -128, -128, 127, 127, -128, -86, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, 127, -128, 3, 49, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, 26, 127, -12, -128, 27, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -87, 127, -128, -128, -53, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -43, 127, -128, 127, -86, 127, -128, -128, -128, -50, 127, 127, -128, 65, -128, -109, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 16, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 65, -128, 127, 127, -128, 127, 127, -128, -128, -21, 127, 127, -128, 127, 127, -128, -79, -128, 127, -128, 127, 127, 53, -128, 1, -128, 127, -128, -50, 127, -128, -117, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 58, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, 15, 127, -128, -128, -128, -128, -31, 127, 127, -128, -128, 127, 127, -128, -128, -114, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -42, -128, -128, 127, 127, 127, -6, -128, -128, 127, 127, -128, -128, 127, 127, 90, -128, -128, 127, -128, -128, 127, 127, 16, -70, 1, -128, 86, -128, 127, 90, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -100, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -43, -128, -24, 127, -64, -128, 127, 127, -128, -128, 127, 109, 127, -128, -128, 18, 127, -109, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, 33, -128, -128, 127, -128, 127, -6, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 80, -128, -128, 86, 127, -128, -128, -128, 127, -128, 127, 127, 127, -128, 127, -24, 127, -128, 73, -128, -44, 127, -87, -50, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 76, -128, -128, 127, -128, -128, -128, -128, -128, 127, 127, -96, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 45, 127, -108, -128, 127, 127, -128, 127, -128, 127, -128, -109, -128, -113, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, 127, -88, -128, -128, 88, -128, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 52, -128, 127, -128, -128, 127, 127, -128, -128, -113, 127, -128, -128, 127, 127, -128, -128, -34, 127, 127, -128, -128, 127, 127, -59, -128, 127, 21, -128, -128, 127, 12, 127, -128, -128, 127, 127, 127, -102, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, -128, 91, 127, -128, 127, 127, -128, -128, 127, -128, 127, -68, 127, -128, -128, 16, 127, -128, -128, 127, 127, -7, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -42, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 74, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -127, -128, 127, 127, 27, -128, -74, 127, 127, 127, 127, -128, -128, 127, -128, 12, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, 53, -128, 127, 78, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 102, 127, 127, -39, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 111, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -95, 127, 127, -128, -128, -3, 127, -96, -128, -128, 127, 127, -103, 127, -128, -128, 127, 127, -106, -42, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -27, 127, 127, -128, -128, 127, 127, -128, -50, -128, 127, 127, 73, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, 21, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 63, -128, 127, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -79, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 101, 127, -50, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -50, -128, 127, -128, 127, -128, 127, -128, 121, -107, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -102, 127, 127, 58, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -33, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 22, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 1, 127, -128, -128, 127, -123, 74, 127, 127, -128, -128, 127, 6, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 28, -28, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 75, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -97, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, 13, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, 112, -128, -128, 127, 127, -128, 127, -128, -128, 16, 127, 73, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, 0, 127, -128, 127, 127, 127, 23, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 52, 127, 127, -128, -128, 127, -128, 127, -128, -128, 127, 127, -128, 98, -128, 127, 127, 127, -128, -128, 127, -3, 127, 127, 127, -128, 21, -128, -128, 127, 127, -11, -128, 127, -128, 127, -64, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -12, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, -128, -128, -128, 127, 127, -128, 127, 47, -128, -128, -128, 8, 127, 127, -128, -128, 127, 127, -27, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 60, 127, -128, -16, 74, -5, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -88, -128, 23, 80, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 33, -128, -128, 127, -103, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 66, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, -52, 127, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 121, 127, 118, -128, -128, -128, -128, 127, 127, -128, 127, -128, 127, -128, 80, 127, 127, -128, -128, 37, -128, -128, 127, -73, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 118, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -102, -128, 127, 127, -128, -128, 127, 127, 80, -128, -128, 127, -128, -128, -128, 127, 127, -112, -128, 127, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -112, -128, 127, -128, 127, 127, -128, -128, 127, 127, -128, 37, 127, 127, 26, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, 37, 117, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -12, -128, -128, 127, 127, -128, -128, 127, 127, 100, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -117, -128, -128, 127, -128, 127, -128, -128, 127, 127, -2, -128, -128, 127, -128, -128, 127, 33, -128, 127, 127, -128, 127, -128, 97, -128, 127, 127, -128, -128, 26, 127, -128, -100, -128, -128, 127, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 65, 127, 127, -128, 122, 127, 80, -128, 127, -128, 127, 127, 127, -128, -128, 127, 64, -128, -128, 127, 127, 127, -128, -128, -128, -75, 127, 127, -128, -128, 127, -128, -128, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -86, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 95, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 0, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -5, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 15, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 76, 39, 127, -128, -128, 5, -128, -128, 127, 32, 127, -128, 127, 127, -128, -128, 127, 127, 47, -57, -128, -128, -128, 127, 127, -128, -128, -128, -7, -128, 127, -128, -128, 127, 127, -90, -128, 127, -128, -128, 127, 127, -128, 127, 26, 127, -128, 127, 127, -128, -128, -128, 127, -128, 0, 127, -128, -128, 127, -128, -128, -128, 127, -128, 127, -128, -128, -128, 127, 127, -128, 127, 127, -22, -128, -128, 127, 127, 64, 127, 80, -128, -128, 127, 45, 127, 127, 127, -128, -128, -13, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, 96, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 74, -128, 127, 6, -128, -32, 127, -111, -76, -128, 127, 127, -128, -128, 127, -128, 127, -93, 127, -128, -128, 27, 127, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 16, 127, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -86, -128, 127, 127, -128, -128, 127, 11, -128, -36, 127, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, 6, -128, 127, 127, -128, -128, -128, 127, 127, -128, -101, -128, 127, 127, -128, 79, 75, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 70, 127, -128, 127, -128, -128, -80, 127, 88, -128, -128, 127, 127, 127, -128, -60, 127, -128, -39, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 31, -128, -128, -128, 127, 127, -128, -128, -33, -128, 127, -128, 127, -116, 127, -128, 79, 127, -128, -128, -128, -128, 127, 107, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -39, 127, -2, 127, -128, -128, 127, -128, 127, 74, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -48, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -128, -128, 109, 127, 127, -128, -128, 127, 127, 81, -128, -128, 127, 127, -128, -128, 127, -128, 87, 127, -128, -128, 127, -128, 0, 127, 49, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, 122, 127, -128, 127, 127, -128, 127, -128, 127, 127, -128, -128, -54, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 109, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 33, 127, -128, -128, 127, 127, -69, -128, -98, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 97, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 54, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -10, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 50, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, -128, -75, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, 127, -128, -90, -128, 127, 127, 127, -128, -128, 127, 127, 73, -128, 127, 127, -122, -22, 109, 127, -128, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 121, -128, 127, -128, 127, 108, 127, -128, 127, 127, 127, -128, -92, -128, 127, -128, -128, 11, 127, 127, 127, -128, -128, -128, 127, -43, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 7, -107, -128, 127, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -38, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 43, 127, -128, -128, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -100, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, -128, 127, -128, 127, -60, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 2, 78, -128, -128, 127, 127, 127, -8, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -27, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, 114, -128, -128, 127, 127, 127, 114, -128, -128, -128, 127, 127, -128, -128, 127, 16, -128, 127, 127, -128, -128, -128, 96, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 108, 127, -128, 22, 127, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 92, -128, -128, 127, 127, -128, -128, 127, -128, 127, -79, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -109, 127, 127, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, -63, -128, -128, 127, 127, 127, -128, -128, -60, 127, 127, 127, -128, -128, 127, 127, -128, -128, -127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, -128, 48, 127, 127, -128, 127, 127, -128, 54, 127, 127, -128, 127, -128, -60, 44, 127, -128, 127, 127, 127, -128, -128, 127, 127, -91, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -38, 127, -128, -128, 127, 127, -128, 66, 127, -128, 127, 116, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 80, -128, 107, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 81, 127, -128, 127, 127, -128, 127, 127, 127, -128, 127, -128, 127, 60, 127, -128, 127, -128, 36, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, -128, -128, 127, -128, -128, 127, -50, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, -128, 58, 127, -128, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, 127, -16, -106, 127, 58, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, -57, -128, 127, 127, -87, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, -128, 127, 68, 127, -128, -128, 116, -128, -128, 127, -128, -128, -70, 127, 127, 127, -128, 127, 127, 127, -128, 127, 66, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -34, 127, -128, -128, 127, 127, -128, 127, -74, -128, 127, 127, -128, 127, 127, -128, -128, -66, -128, 127, 127, -128, 127, 127, -119, 127, -128, 28, -44, 127, -128, -128, 119, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, 127, 127, 111, -128, 108, 127, 127, -128, 73, -128, 127, 127, -128, -128, 119, 127, 127, -118, -128, -47, 127, -128, 127, 127, 127, -128, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, -128, -128, -36, 127, -128, 127, -128, 127, -128, 127, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 36, 127, 122, 127, -128, 127, -128, 127, 127, -128, 127, 127, 127, -128, -128, 127, 127, -128, 21, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 114, -128, -128, 127, 127, -128, -128, -128, -15, 127, 127, -128, -33, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 127, 127, -128, -128, 127, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 3, -128, 127, 127, -128, -128, 127, -128, 18, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, 38, -128, -76, 127, -128, 127, 116, -128, -128, 127, -128, -128, -128, 127, 127, -10, -128, 127, 127, 127, -128, 64, -128, 127, -128, 127, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -128, 127, -128, 127, 63, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 127, 127, -128, -128, 101, 127, -118, 127, -128, 127, 127, 127, -128, 127, -128, 127, -128, -128, 81, 127, 127, -128, 31, 127, 127, -128, -128, 127, -128, 127, -128, -33, -128, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 64, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, 113, 127, -39, -128, -128, 127, 127, 50, -128, -128, 127, -90, 127, -128, -128, -128, 127, -114, -128, -128, 127, 127, -128, -128, -128, -52, -86, -29, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, 27, -128, 127, 127, -32, -128, 101, -128, 127, 127, 127, -128, 127, -128, -128, 127, -128, -128, 127, 127, -128, -128, 127, 127, -116, -128, 127, 127, -128, -128, 127, -128, 127, 127, -128, -92, 127, -128, -128, 127, 127, -128, -28, -128, 127, -128, 127, 22, 127, -128, -128, -128, -128, 127, 127, -128, -128, 127, -128, -38, 127, -128, -128, 127, 127, 127, -128, -128, 127, 127, 127, -74, -6, -128, 127, 127, -128, -98, 2, 85, -128, 127, 127, -128, -128, 127, -128, -18, -128, 127, -128, 127, -128, -128, 127, -128, 54, 127, -128, 37, 127, -128, 85, 127, -128, -128, 127, 127, -128, 127, -128, 127, -128, 127, -128, 127, 127, 127, -128, -128, 127, -128, 112, 127, -128, -128, 127, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, -128, -128, 85, 127, -128, -128, 127, 127, -128, -128, 127, 92, -128, -128, -128, 127, -122, 127, -128, 127, -128, 45, 55, 127, -128, -128, 70, 127, 127, -128, 127, 127, 127, -128, 24, -128, 127, -128, 107, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, 127, -128, 127, 127, -128, -128, 127, 127, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, -128, 81, 127, 127, -128, -128, 24, 127, -128, 127, -128, 87, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, -128, 127, 127, 109, -128, 127, 127, -128, -128, 127, -128, 127, 127, 127, -128, 127, 127, 59, -128, 127, -128, -128, 127, 127, 127, 127, -122, -128, -128, 127, 127, -128, 127, -128, -128, -128, 127, 127, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, -128, 127, -128, -128, 127, 127, -128, -128, 52, -128, 127, -128, -128, -52, 127, -29, 127, 127, -128, -128, 127, 127, -128, -128, 127, 117, -128, 127, -128, 127, 127, -128, -38, -128, 127, -128, -48, -128, 127, -128, 127, 127, -128, 117, 127, 127, 127, -128, -128, 127, 127, -6, -128, 127, 117, 127, -128, 127, 32, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, 127, -128, -128, -128, 127, -128, -128, -128, 127, -128, -128, -128, -128, 127, 127, 127, -128, -128, 127, -24, -128, -128, 127, 127, -128, -128, 127, 127, 127, 33, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 16, 112, -128, -128, 127, 127, -128, 127, -128, 127, -128, -128, -128, 127, 127, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, 127, -27, -128, 127, -128, 127, 127, 127, -128, 127, 127, -96, -128, -128, -128, 127, 127, 127, 127, -128, 23, -128, 127, 127, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, 22, 127, 39, -100, -128, 127, -118, -128, -128, 127, 127, -128, 127, 127, -128, -128, 55, 127, -128, -128, 127, 127, -109, -128, 127, -128, -128, 127, 127, -128, 127, 127, -128, -128, -128, 127, 127, 127, -22, -128, -128, 127, -128, -128, 127, 127, 31, 127, -63, -128, 127, -128, -128, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, -71, 127, -128, -128, 127, -128, -128, 127, -128, 127, -128, -128, -85, 127, -128, -128, -128, 127, 127, -128, -65, -128, -128, 59, 127, -128, 127, -128, -60, 127, 127, -128, -128, -128, 127, 127, -128, -128, 127, -128, -128, 87, 127, 127, -128, -128, 127, -128, -128, 127, 127, -128, 127, -128, 127, 38, 127, 127, -128, -128, 127, 127, -128, -128, 127, 127, 127, 11, 127, -128, -128, 127, 127, -128, 127, 127, -128, 127, 127, 127, 127, -128, 127, 127, -128, -128, 127, 127, -128, -128, -28, 127, -6, -128, 127, -128, -107, 127, 127, -128, -128, 127, 73, -128, 127, -128, -128, 127, 127, 127, -21, -128, 127, 127, 127, -128, -128, 127, 127, -128, -80, 34, 127, -128, -128, 127, 127, 109, 0 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
