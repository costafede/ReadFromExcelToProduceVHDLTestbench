-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
            1, 17, 11, 12, 18, -16, 1, 10, -13, -1, 0, 4, -19, 14     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -7, -21, 102, -124, -77, 22, 10, 45, -41, 22, -82, 122, -34, 7, 94, -99, 48, 32, -38, 13, -81, -84, -8, -18, 95, 113, -67, 44, 60, -84, 20, -45, 77, 124, -51, 15, -110, -47, -60, -55, 19, 107, 32, 74, -69, -99, -79, -4, -25, -36, 61, -85, -79, 101, -81, -58, -32, -117, -54, -43, 85, -85, 109, -50, -59, -27, 30, 90, 87, -76, 1, 98, -2, 117, -109, 10, -86, -55, -83, 40, 31, -18, 108, -123, -69, 105, -126, 126, -60, 93, -47, -23, 14, -104, -14, 124, -54, 60, 46, 103, -100, 13, -59, -24, -54, 38, 31, 33, -13, -67, 20, -2, -42, -47, -7, -11, -60, 82, 35, 63, 109, 68, 96, -89, 19, -90, 52, 99, -70, 4, 7, -86, 125, 111, -102, -122, -41, 112, 81, 64, 83, 2, 106, -67, 25, -86, 78, 93, 68, -17, 41, 60, 7, -81, -115, 79, 19, -14, -5, -56, -9, -57, 4, -70, -18, 1, 14, -51, 11, -73, 29, 118, 62, 113, 72, -105, 81, -7, 98, -105, 12, 100, -117, 112, -70, 6, 28, 49, 113, 122, -48, -17, 43, 83, 119, -50, -121, 10, 89, -117, -12, 80, -11, -98, 82, -102, -127, 23, -40, 2, 61, 107, 106, -26, -15, -89, 27, -83, 22, 14, 121, 117, 86, -102, 108, -82, 77, -9, 86, 29, 99, -56, 44, 22, 108, 72, 58, 29, -24, -107, -7, 94, 83, -117, -103, -83, 14, -42, 50, 123, -117, -56, 82, 63, -107, 95, 66, -124, -93, -72, -93, 0, 81, -40, 48, 59, 104, -7, 21, 69, -70, -101, 39, 23, -62, 52, -15, -56, 82, -22, -36, 15, -65, -95, -123, 22, 15, -128, 27, 88, 62, 9, 113, 70, -70, -74, 90, -107, -3, 8, 13, -96, 18, -12, 69, 21, 97, -29, 67, 33, -12, -99, -123, -30, -42, -86, -121, 47, 64, -46, 6, 78, 54, 68, 21, -81, 20, 31, 45, -59, 65, 102, 85, -16, -40, 96, -96, 27, 3, -72, 18, 51, 50, 21, 63, 112, -29, 103, -85, -25, 118, -99, 32, 13, -11, -71, 98, 37, -44, -117, -79, -119, -38, 106, 21, 101, -57, 65, 51, -41, -33, -115, -37, -118, 79, 84, 2, -83, 113, -39, 41, -104, -128, -106, 117, -68, 36, -46, 109, -124, -28, -16, 22, -57, -83, -38, 92, -101, 95, 116, -106, 38, 100, -26, 118, -68, 34, 123, -24, -61, 67, -87, 89, -34, -64, 26, -60, -14, -14, -6, 90, -90, -113, 88, 9, -72, -10, 54, 78, 50, 95, 37, -10, -120, 66, -9, 120, 17, 74, -98, 1, -70, -57, -47, -1, -120, 117, 91, 122, 99, -111, -73, -74, -17, -88, -40, 30, -63, -87, -68, -77, -38, 112, -115, 41, -107, -91, -94, -36, -72, -46, -25, -15, 10, -56, 110, -79, -7, -35, -65, -29, -106, -22, 89, -90, -82, -12, 116, -73, -51, -87, -7, -119, 95, 71, 116, 91, 111, -109, -6, -85, -82, 78, -76, 33, 87, 106, 29, 7, -11, 6, 48, -59, 90, -76, 50, 90, 56, -45, 16, 31, -105, -106, 69, -81, 99, 29, -49, -100, -111, 100, 93, -97, 27, 88, 93, -8, -66, -122, -42, -112, 11, -79, -108, 99, -59, -42, 90, 110, 52, 29, 7, -71, 28, -83, 11, 56, 103, -4, 32, 81, -16, 43, 53, -4, 51, 103, -84, -11, 68, -117, 57, 118, -75, -38, 74, 25, 20, 13, -58, -10, -100, 59, 24, 125, 89, 113, 35, -56, -107, 60, -79, -65, -38, 23, -124, -127, 120, -95, -123, -123, 93, -61, 62, 101, -83, 122, -89, -85, 55, 63, 32, 86, 25, 83, -80, 119, -118, 21, -42, -64, -14, -110, 84, 84, 16, 45, 54, 93, 10, -100, 54, -95, -15, 110, 64, 37, -95, 41, -127, -123, -127, -119, 64, -26, -75, -72, -15, -20, 123, 45, -6, 24, -127, 74, 126, -2, 99, -112, -91, -25, -18, 119, -49, -70, -12, 122, -118, -46, 104, 51, -113, -16, 74, -62, -39, 92, -99, -69, 96, 103, 123, -123, -16, 104, 123, 77, 88, -67, -97, 40, -42, 124, 44, -87, -128, 122, -44, 69, 64, -113, -64, 104, -90, -57, 40, 13, 21, -7, -104, 55, -34, 98, 66, 20, 74, 85, 18, -35, 73, -26, 16, 0, 26, 102, -89, -60, -119, -119, 85, -94, -62, -73, 54, -64, 30, 112, -113, 85, -60, -125, 44, 119, -34, 23, 2, 58, -36, 56, 8, 33, 50, -93, -73, 42, 87, 2, 122, 34, -39, 84, -70, 14, 66, 82, 78, 125, 76, -88, 33, -110, -117, -98, -26, 31, 66, -55, 24, 27, -108, 44, 38, -47, -102, 5, -86, -79, 26, -58, -51, -54, 118, -70, -4, -90, 69, 33, -70, -101, -30, 98, 27, -122, -113, -127, -123, 55, 62, 38, 34, -46, -121, 28, -27, -94, 5, -69, 89, -72, -59, -8, -97, -77, 78, 42, -64, -63, 5, -82, -3, 108, -64, 14, -92, -72, 31, -59, 32, 111, 9, -54, 124, 21, 0, -33, 123, 77, 11, 101, 82, -53, 95, -68, 66, 7, -58, -125, 8, -1, 119, -42, -6, -123, -121, 76, 6, 33, 38, -126, -104, -60, 28, -55, -80, 102, -115, -79, -81, -41, 24, 43, -72, 48, 36, -6, 113, -65, -49, 106, -119, -86, 67, -74, 124, -10, 36, -113, 57, -74, 13, -88, 30, -96, 117, 16, 96, 16, 111, 91, 98, 112, 53, -23, -99, -63, -87, 126, -116, 47, -97, -54, 56, 32, -70, -37, -90, 76, -46, 120, 91, -121, -116, -99, -101, 83, -33, 72, -88, 127, 1, 64, 35, -56, 116, 110, 30, 43, -82, 37, -95, -31, -15, 57, 19, 125, -70, 113, -8, -79, 65, -93, -71, 33, 54, -79, 119, 112, -64, 116, 99, 91, 37, 35, -114, 43, -111, 28, -96, -47, 45, -33, 95, -126, 22, 66, 54, 2, 116, 69, -63, 58, 82, -80, 103, -65, -39, 104, -29, 108, -32, 116, -94, -101, 63, 118, 116, 118, 42, 42, 26, 26, 81, -67, -68, 6, -35, -53, 38, -104, 54, -21, -30, -90, 68, -29, -105, -71, 67, -93, 103, 24, 25, -44, 61, -97, 96, -28, 108, 126, 37, 63, 117, -37, -112, -33, -96, -104, 53, -23, 43, 76, -14, -82, -46, -106, -29, -74, 24, -109, 24, -65, 46, 122, 36, 105, 53, 8, -94, 104, -50, 99, 15, 1, -55, -123, -19, 48, 19, 8, 76, -12, 38, -117, 23, -105, 118, 39, 109, 63, -85, -9, 53, -50, -50, -55, -62, -68, 42, 95, -27, 26, -10, 115, -72, 0, 41, 72, -27, -86, 34, -2, 112, -121, 84, 59, 35, -44, -67, -30, 119, -12, -39, 15, -78, 21, 23, -3, -1, -106, -73, -8, 92, 11, -66, 111, -98, -10, 53, 50, -64, 78, 73, 94, -107, 25, -33, 27, -51, 42, -26, -21, -11, -49, 105, -63, 15, -54, 56, -119, 70, -115, -123, -111, 118, 47, -26, 97, -97, -4, 18, 84, -43, 8, -72, -17, -96, 109, 3, -27, 3, -65, 74, 106, -18, -2, -126, 103, 83, 73, -125, -102, 46, 40, 13, 60, -110, -88, -74, 49, 94, 95, 42, -7, -118, -113, -61, -123, -74, 103, 89, -116, 92, 44, -41, -22, -33, 61, 28, 25, -87, -18, 59, 45, -9, 97, -19, -97, 21, 65, 95, -18, -66, -109, 7, -47, -89, 78, -92, -91, 4, -35, -85, -15, -6, -46, 21, -10, 23, 22, 85, 15, 82, 73, -29, -48, -106, 118, 87, 85, -52, 94, -55, -3, -78, 13, 47, -17, 125, 110, 92, -56, -60, -15, 84, -90, 43, -69, -45, 114, 40, 31, 28, -5, -70, 19, -10, 87, 119, -25, 91, 52, 93, 64, 17, 48, 62, -91, 127, 113, 38, 55, -118, -26, 24, -63, -19, -92, 111, 59, 42, -30, 97, 29, 17, -2, 44, -115, -9, -102, -55, -104, 100, -98, -70, -42, 27, 127, 85, 4, -76, 6, -7, 7, -124, 76, -4, -99, 61, 97, -32, -105, -4, 71, 11, -70, 63, -110, -87, 15, -30, -17, 106, 124, -55, -83, 109, 78, -93, -94, -98, 9, -98, 10, -122, 71, -33, -90, 63, -114, 13, 82, 59, 0, 116, -63, 30, 78, 73, -109, 29, -28, 59, 105, -13, 99, -82, -77, 119, -2, 99, 120, 47, -84, -82, -118, 115, 126, -84, 81, 30, 97, 98, 127, -51, 77, 55, -96, 95, -23, -125, -116, -44, 7, 83, -123, -121, -94, -109, 115, -7, -114, 75, -99, -52, 57, 57, -72, -22, 75, 59, 74, 108, -29, -120, -11, 109, 120, -3, -34, 118, -100, 88, 65, 109, -31, -42, -123, -69, -27, -23, 83, -99, 62, 96, -121, 61, 66, -24, -100, 34, 107, 67, -15, 120, 30, -42, -65, -53, -85, -78, 81, 70, 33, -31, -60, 15, -102, 15, -111, -19, 37, 9, 67, -83, 47, -72, 127, -3, -22, -20, -98, -113, -69, -88, 77, 56, 80, 44, 22, 24, 55, 85, 14, 16, 47, 25, -95, -54, -120, 21, -100, -10, 87, -39, 106, 97, 36, -49, -101, 35, -4, 124, -112, 74, -7, 125, 126, 102, -2, -80, 22, 100, -65, -123, -31, 21, 91, -85, 63, 55, 13, 111, -19, -109, 32, 80, -45, -100, -70, -29, 97, 68, 58, -90, -81, -76, -35, -101, -120, -37, -75, 102, -9, -101, -104, 98, 57, -73, 124, -81, -52, 33, 3, 126, -8, -68, -49, -26, -109, 39, 99, -8, -118, -93, -5, -34, 66, -22, -109, -55, 72, -55, 84, -90, 122, 107, -122, -109, 38, 65, -104, 106, 11, 5, 43, -14, 93, 75, -84, -35, 20, -116, 60, 83, 77, -70, -83, 122, 10, -73, 100, 123, 104, -114, -55, 27, 24, 77, 20, 110, 23, 56, -50, -91, -82, -116, -126, -83, 81, 120, -48, 104, -32, -65, 111, -10, -101, 58, -127, 51, 119, -44, -15, -77, 85, -105, 101, -19, 12, 19, -67, 24, 48, 5, 2, 55, -30, 58, 58, 57, 27, -121, 85, 2, -25, 42, 116, -41, 28, 120, -55, 103, 60, 33, -68, -32, -91, 17, 31, -3, -9, -79, 84, 11, 29, -95, 18, -7, 44, 102, -85, 30, 65, 48, -27, -62, 18, -96, -49, -106, 44, 31, 124, -27, -124, 90, -53, 61, -120, 127, 5, 92, 118, 36, -49, 4, -128, -12, 41, 86, 59, 67, -113, 120, -96, -1, 122, 22, -86, -116, -119, 92, 81, 101, 110, 37, -30, 127, -88, 99, -22, -121, -88, -58, 66, -32, 15, -2, -124, 72, 18, 101, -128, 62, 41, 47, 108, -101, 20, -66, -125, -85, 12, 9, 64, 68, 28, 14, 83, -65, 81, -62, -58, -73, -112, -55, -81, -29, 57, 29, -105, 74, -29, -88, 124, 93, 127, -25, 31, -119, 1, -2, 90, -75, -110, 50, 90, 94, 92, 27, -120, -66, 111, 24, -101, -124, 107, -115, -120, -63, 106, -51, -103, 21, 46, 1, -94, -89, 81, -82, 96, 75, 113, -3, -99, 42, 18, 73, -3, -84, 107, 94, 71, -66, 19, 91, 57, 18, -21, -83, -118, 22, -69, -77, 14, 64, -10, -33, 53, 77, -40, 77, -27, 3, -76, 100, 45, 40, 39, 97, 14, 65, 125, 21, 118, -10, -101, 33, -22, 79, 39, 66, 86, -21, -60, -47, 73, 62, 93, 13, 53, -60, 107, -104, 119, -20, -74, 28, 4, -117, 116, 30, -60, -53, -43, 87, 16, -97, -43, 39, -35, -96, -91, -81, 98, 117, -17, -100, -107, 87, 91, 59, -21, 73, -20, 27, -87, -125, 50, 38, -51, 92, 46, 19, 57, 25, 73, 106, -73, 28, 98, -105, 57, 0, -57, 15, -19, 107, 50, 35, 48, -64, -33, 73, 6, -26, 30, -14, 98, -91, 48, -80, 52, 109, -106, -29, -112, 54, 45, 64, 16, 40, 96, 118, -58, 79, 89, 42, 53, 97, 24, -34, 75, -89, 121, 0, -73, -8, 74, -29, -10, -83, 49, -58, -38, -17, -44, -34, 6, -84, -106, -86, -65, 76, 59, 22, -57, 109, 4, -16, 45, -20, -37, 46, 64, -19, 42, 4, -77, -42, -118, -102, 92, 52, -40, 27, -85, -117, 70, 109, -21, -75, 96, -48, -84, 12, -39, 81, 40, -11, 2, 93, 117, 33, 52, -90, 92, 47, 60, -110, -4, -87, -51, -64, -82, 74, -38, 11, -28, -26, -54, -17, -108, -33, -35, -86, -120, 68, 6, -35, 91, -2, -52, -88, 90, -3, 69, -19, -34, -24, -33, 98, -17, 55, 70, 83, 19, 98, 55, 45, -27, -25, 52, -33, 94, -89, 117, 118, 126, -98, 96, -16, 0, 70, 107, 119, -128, 65, 8, 59, 31, 94, 25, -37, 97, 103, -120, 60, 107, 98, -95, -101, -77, -107, 66, -110, -22, 19, 27, -80, -50, -44, -8, 125, 44, 39, 119, 82, -52, 88, 1, 124, 87, 107, -93, 92, -91, -10, -11, -67, -56, -17, -101, 92, -76, 110, -71, -116, -93, -108, -69, 93, 72, -8, 46, -91, 120, 45, 79, 97, 63, 52, 95, -104, 68, -57, -54, 4, -103, 111, 121, 13, -27, 23, 52, 113, 15, 38, 66, -20, 62, -68, 1, 62, 73, 39, -67, 70, 44, 70, -121, -79, -45, -58, 116, -12, 44, 19, 22, 61, 43, -8, -22, -31, 110, 103, 90, 56, 73, 16, 92, -70, 59, 71, -32, -71, -91, 8, 19, 57, 29, -77, -28, 112, -24, -7, -92, 28, -75, -4, -92, 61, 63, 10, -102, -82, 103, 45, 127, -70, -97, 74, -23, -101, -60, 12, -113, 69, -61, 127, 100, -53, -48, 9, -28, -87, 100, -40, 7, 54, -101, -94, -76, 109, -26, -124, 96, -3, 7, -61, -30, 53, 100, 17, -44, -16, 24, 86, 63, -6, 89, -98, -50, 108, -17, -128, 76, -57, 8, 50, -29, -101, 46, 34, 41, 90, 15, 34, 25, -34, -45, 119, -104, 52, 53, -80, 118, 60, -22, 72, 2, -66, -36, 42, 123, 9, 65, -118, 51, -43, -85, 35, -72, 6, -124, -6, -80, -7, 76, 55, 25, -6, -35, -103, 108, -3, -39, -57, -93, -67, 25, -128, -128, -24, -3, -117, -77, 53, -96, 99, -52, -5, -3, 73, 8, 96, 53, -45, 2, -83, 46, -21, 60, -92, -68, 38, 96, -76, 99, -37, -96, 22, 90, -109, -80, -80, 127, -90, -26, -64, -16, -64, -123, -77, 19, 20, 53, -26, 111, -29, -1, 93, -89, 4, 126, 122, 0, 53, -40, -118, -25, 45, 30, -114, 7, 14, -80, -17, -120, 11, -113, 71, -127, -26, -96, 106, 64, -61, -44, -24, 89, 84, 123, -4, -108, -58, -87, -62, 121, 19, 96, -79, -121, -123, 96, -123, -113, 101, 28, 46, -35, 81, 75, -59, 32, 28, -22, 46, 62, 43, 24, 89, -21, -83, -91, -99, 111, 88, 41, -55, -123, 125, 0, -60, 108, 61, 88, 14, -63, 35, 69, -88, -89, 41, 74, -108, 66, 27, 80, -67, 76, 119, -18, 48, -60, 40, -24, 110, -79, -121, 111, 95, 80, 15, 71, 29, -116, -106, -32, 89, 7, 2, -52, -69, -95, 63, -54, 109, -81, 26, -74, 58, 57, -10, 72, 97, 22, 31, 75, -29, 44, -4, -83, -17, -125, 25, 18, 45, 92, 55, 98, -23, -32, -21, 104, -27, -34, 119, 2, 74, -112, 104, 68, -11, 31, -103, -102, 123, 94, -49, 49, 116, 107, 71, 72, 82, -8, -26, 80, -91, 88, -103, 79, -12, 69, 55, -97, -124, -114, -32, -55, -13, -66, -66, 112, -16, -48, 39, -44, 77, -51, 104, 33, 127, 51, 60, 20, 116, 35, -42, 111, 9, 95, 64, 7, -72, 108, 103, -50, 80, -110, 59, -55, 27, 95, 51, -71, -24, -105, 72, -39, 81, -2, -69, -89, -69, -84, 36, -72, -22, 13, -120, -86, 85, 70, 111, -21, -100, 88, -40, -68, -60, 123, -78, -47, 106, -92, -22, 108, -110, -56, -108, 47, -81, 38, 82, 34, -31, 49, 103, -122, 95, -69, 59, 54, 0, 16, -41, -97, -17, -101, 102, 44, -73, 87, 97, -101, -8, 36, 112, -47, -79, 49, 103, -42, 35, 37, -14, -105, 43, 110, 35, 69, -72, -55, -57, 42, 91, 113, 76, 117, 23, 20, 75, -120, 0, -47, 40, 17, 89, 28, -104, -101, -14, -51, -66, 36, -69, 19, -19, -10, 32, -104, -102, -38, -49, 79, 28, 61, -68, -87, -30, 6, 119, 0, 31, 51, 35, 21, 93, -55, -67, 30, 75, -42, 127, 27, 70, -80, -32, 11, 47, -46, 32, 34, 117, 121, -128, -88, 61, 22, -2, 1, -127, 62, -82, 73, 47, 85, 33, -85, -94, -53, -120, 125, -48, -100, -56, -113, -105, 14, -88, -16, 85, 17, -99, -68, -28, 59, -37, 63, 18, 17, -11, -1, 40, 115, -121, -86, -93, -71, 21, -88, -44, -87, 83, 26, 69, -61, 41, 94, -43, -11, 68, -27, -104, -89, -14, 33, -2, -91, -88, -47, 95, 9, 110, 122, -79, -63, 103, 94, 82, -95, -111, 127, -82, -120, -120, -89, -33, -69, 21, 73, 68, 53, 111, -106, 103, 115, 80, -52, -101, 47, 56, 27, -97, 25, -102, -51, -113, -92, 80, 7, -64, 30, 99, 67, 37, -5, -67, 89, -31, 119, -76, 36, -128, 121, 103, 1, -75, -71, -41, -105, -126, -25, -30, 17, -79, -107, 25, -110, -109, 68, 121, 111, 110, -74, -85, -27, -99, 72, -5, -77, -81, -93, 96, -102, 74, 115, -57, 32, -113, 0, 54, 108, -23, 117, -16, -124, -78, 84, -53, -78, 12, 2, -113, -6, 7, 19, 0, 65, -17, -34, 11, -22, -110, -48, 117, 54, -87, 13, 30, -118, -100, 44, -4, -1, 56, -77, 78, -124, 90, 26, -31, 0, -22, 79, 81, 51, -97, -116, -85, 38, -3, -113, -105, 102, -123, 85, 39, 0, 15, 7, -105, 34, 47, -9, 25, 67, 12, 3, -56, -50, 2, -85, 27, -88, 119, 97, 87, -78, -105, 20, -63, -12, 127, -120, 54, -119, 97, -113, -43, -74, -28, -21, 17, 67, 90, 24, -94, -69, 104, -18, -8, 126, 121, 72, -67, -44, 2, 52, -22, 113, -24, -94, 87, -104, 40, 62, -72, 5, -81, 115, 12, 54, 48, 113, -21, 56, -103, -24, -8, -59, -16, -94, 10, -32, -40, -55, -101, 19, 84, 45, 109, -119, -95, -82, 125, -60, -4, 57, -36, 103, -17, 110, -43, 29, -123, -35, 28, 85, 5, 71, 110, -81, -75, 112, 69, 80, -121, -15, -82, 49, -82, -72, 106, -12, 47, -118, -78, -95, 90, -6, 103, 5, 6, -63, -78, 30, 65, 12, -21, -43, 13, 9, 2, 99, -124, -77, -85, 21, 86, -9, -74, 4, 120, 47, -111, 26, 37, -102, 72, 70, 12, 11, -75, 88, -109, -108, -24, -56, 71, -96, -92, 110, 8, -114, -18, 49, 33, 99, 123, 76, 125, -53, -92, 87, -92, 120, -16, 64, -13, -5, 69, 66, 41, 1, 48, 109, -1, -67, 68, 7, 72, -47, 62, 49, 16, 85, -40, 3, 16, 95, 107, 29, -57, 67, 126, -106, 26, 9, 60, -80, 33, 66, 19, 65, -23, -127, 30, -74, 49, -94, 31, 106, -28, -75, 102, 50, 45, -75, -5, -94, -67, -103, 110, 121, -56, -105, -52, 46, -8, 80, 80, -35, 68, 16, 23, 109, -49, 85, -74, -9, 63, -10, -104, 2, -102, 97, 61, -81, 104, 99, -125, 102, 0, 86, -67, 32, -18, -24, -72, 102, 29, -64, -50, 82, 84, -89, -18, -89, -64, -124, -1, 54, -89, 107, 125, -25, 35, 85, 53, 75, 61, 11, -44, -4, -72, -81, 115, 114, -38, -40, 1, -118, -19, -101, -12, 47, 16, -55, -35, -19, -22, 45, 37, 107, -122, 92, -39, -53, 5, -16, -33, 94, -50, 24, -82, -85, 41, 12, -1, -100, 46, 90, -33, 4, 119, -19, 23, -28, 21, -74, 70, -40, 92, 68, -37, -9, 50, -128, -35, 113, 28, 42, -19, -51, 6, -27, 24, 104, -96, 111, 63, 115, -51, 36, -74, 42, 126, 70, 17, 87, -122, 113, -3, 11, 33, 121, -87, -7, -27, -51, 123, -24, -2, 68, 95, -40, 109, 4, 67, -12, 111, 28, 1, -52, -2, 39, 80, 91, 31, 22, -49, -64, -10, 20, 50, 13, 1, 109, -32, 58, 24, -13, -26, -99, -107, 123, 2, 11, -2, 8, 60, -2, -104, 18, -121, 125, -35, 96, -1, -31, 10, -121, -103, -119, 49, 12, -24, 48, -2, -60, 29, 100, 11, 108, -123, -8, -36, 1, -119, 49, 0, 10, -85, 98, 84, -67, 27, -71, -124, 104, -36, 41, 127, 125, 127, -112, -87, 79, -73, -66, 23, -70, 116, -70, 49, -63, -78, -60, 81, 10, -124, -9, -77, -26, 113, -7, -33, 16, -104, 10, 93, -100, -117, -57, -71, 111, -20, -49, 123, -56, -128, -84, 110, -127, -79, -61, 115, 113, 10, -101, 66, -100, 101, -50, -40, -24, -50, 66, 25, 118, -44, 28, -84, 67, -114, -83, -122, 50, 115, -119, 26, -58, -75, 60, 93, 86, 109, -23, -38, -107, 2, 101, -58, -128, -29, 66, -104, -8, -100, -112, 85, -13, -59, 88, 117, -25, -55, -92, -114, 116, 12, 28, -23, 49, 62, -9, 103, -112, -78, 116, 86, -77, 44, 35, 26, 15, 97, 87, 54, -125, 31, -65, -93, -85, 34, -101, -93, -6, 99, 109, 21, -8, 13, 70, -52, -124, 100, -55, 76, 119, 110, -25, -93, 14, 68, -12, -127, -47, -70, 9, 39, 74, -18, -84, 42, 3, 116, -48, 37, 79, -126, -40, 115, 70, 56, -96, -110, 74, 44, -68, 13, -25, -127, 52, 72, 96, 99, 19, 1, 10, -96, 9, 52, 15, -70, 30, -10, -91, -35, -52, 66, -51, 67, -9, 39, -78, -102, -95, 14, -8, 85, 97, 64, 93, -78, -54, 69, -52, -66, 13, -98, 72, -101, 84, 103, -125, -21, -122, -87, -71, 2, 72, -95, -23, 124, -91, 83, 116, 68, 115, 46, 94, 125, -96, 116, 75, -68, 60, -78, 105, 83, 96, 32, 58, 89, 90, 99, -63, 3, -51, 120, 103, 13, -123, 126, -1, -73, -24, 75, -66, -44, -77, -47, 25, -19, -105, -121, 57, -100, -75, 46, 82, -28, 15, 12, -54, 82, -88, 10, -106, 120, -122, -67, -24, -89, 92, 27, -27, 115, -9, 28, 54, -61, 125, -120, -83, -57, -51, -124, 90, -30, 23, 94, 108, -70, 20, 75, -62, -76, 70, -115, 27, 64, -72, -19, -12, 4, -48, -79, 67, -3, 114, 72, 98, 22, 39, -107, 104, 30, 96, 79, -115, -48, 62, 61, 19, -120, 24, 110, 6, 58, -8, -58, 34, -128, 110, 97, -102, 42, 106, 30, -30, 109, -29, -113, 8, 91, -102, 19, 63, -5, -27, 115, 32, -29, -124, -62, -24, 117, -15, 106, -45, 47, 46, 13, 28, 71, -96, -79, -9, -41, 86, 52, -4, -46, -115, 70, 126, -93, -75, -70, -51, 8, -78, 116, 85, -26, 118, 82, 109, -51, -30, -10, -49, -126, -111, -20, -111, -121, 69, -39, 5, 27, -21, 85, 53, -30, 29, 99, 13, -49, 23, -19, -16, -108, 56, -16, -123, -3, 125, 45, -37, -55, 37, -79, 60, 6, 35, -23, 88, 42, 47, 119, -75, -8, -62, -75, -83, 45, -75, -58, -21, -94, -99, 105, 67, 95, -82, -95, 105, -94, 92, -10, -29, -60, 1, -48, 21, -31, 36, 82, 0, -34, -96, 0, 43, -41, -35, -30, -51, 83, 93, -127, 46, 9, -128, -32, 12, -45, -96, -95, -15, 11, 43, -98, 33, 78, -29, 105, 112, -8, -34, -86, -30, 23, -12, 39, 8, 71, 45, 124, 27, 88, 54, -56, 87, -99, 37, 88, 121, -9, 51, -13, -60, 65, -45, 53, -86, -35, 114, -59, -34, -97, 76, -5, -115, -57, 24, -104, 111, 45, -29, -64, 29, -124, -8, -111, 119, 102, 49, 34, -30, -16, 39, -76, -109, -66, -106, 57, 16, 85, -26, -92, -25, -63, -19, -56, 28, 95, -68, -15, 47, -57, -34, 93, -88, 112, -75, -128, -99, 105, -29, -69, 90, -58, 41, 80, 48, -92, 41, 24, 77, -74, 51, 116, 53, 26, 48, -107, 3, 51, -21, 40, 41, 96, -62, -16, 126, 86, -76, -21, 31, -53, -23, 67, -45, 69, 96, -63, 90, 33, -92, -92, -66, -87, -91, -82, 38, 42, -64, -81, 48, -64, -88, -122, -52, -26, -110, -127, -25, -24, 96, -27, 51, 14, -50, -111, 95, -40, 85, 119, -105, 34, -27, 52, -35, -108, 36, 21, 22, 89, 11, 15, -37, -125, 68, 109, 13, -47, -75, -64, -58, -45, 67, 105, 121, -12, 23, -15, -79, -96, -81, -80, -86, -70, 81, -66, 107, 44, 115, -71, 0, -17, 112, 121, -56, -43, -79, 55, -12, 92, -83, 90, 124, -114, 51, -128, 31, -72, -22, -124, -43, -81, 69, -81, -91, 87, 92, 5, 110, 20, 40, -30, 86, 17, -47, 66, -92, -98, -84, -47, -96, 120, -40, 34, -56, 9, -13, 27, 36, -22, -110, 122, 33, -49, 22, -47, -39, -12, -124, 15, 25, 85, -110, -71, -13, 94, -109, -121, -81, -117, 40, -26, -127, 126, 86, 49, 64, -22, -122, -40, -79, -30, -9, -21, -124, -119, 71, -10, 88, -85, 3, -61, -104, 127, -61, 67, -89, 102, -36, -92, -7, -60, -48, -96, -64, 49, 114, 122, -46, 28, -94, 31, -85, 75, 72, -109, -83, 28, -9, -24, 7, 25, 63, 84, 74, 98, -71, -37, 50, 56, 14, 110, 44, 117, -23, 27, 61, 32, -90, 40, -96, 33, -103, 75, 55, 82, 85, 73, 14, -54, -108, -120, -57, 43, -9, -35, -9, 80, 74, -126, 52, -24, -60, 64, -100, -31, -59, 117, 48, 7, 23, 85, 32, -20, 113, 49, -119, 97, -6, -70, -101, -87, -3, 34, -114, -4, 123, 30, -96, 70, 105, 59, 19, 113, 110, 20, -94, 111, -67, 57, -126, -106, -52, -29, 25, 81, -53, 35, 43, -111, -12, -63, 124, -78, 42, -118, -72, -25, 79, -24, 51, 120, 36, -73, 95, 38, 18, -56, -119, -124, 116, -54, -21, -18, 32, -95, 9, -10, 27, 89, 63, 80, 50, -12, 45, 88, -44, -23, -93, 53, -111, -112, -80, 124, -125, 85, 52, -101, -49, 29, 18, 17, 77, -90, 112, -25, 65, 25, 53, -82, 54, 98, -124, 6, 45, 41, -77, -72, -8, -6, -100, -114, 127, 85, 90, 33, 70, -108, -111, -121, 76, 31, -86, 41, -114, 0, 112, -73, -11, 15, 95, 85, -15, 55, 46, -119, 116, 7, 126, 62, -31, 81, -49, -46, 70, -80, 113, -87, 8, -72, -78, -17, -46, 17, 73, 109, 101, 25, 17, -84, 45, -70, -89, -84, 64, 122, 47, 64, -15, 3, 25, -58, -81, 56, 35, 3, 38, 44, -83, -119, 81, -76, -44, -51, -8, -59, -49, 52, -31, -101, -19, -94, -125, -83, 51, -28, -80, -33, 33, 17, -95, -79, -106, -88, -61, 104, 32, -93, 43, -46, 31, -62, -3, 119, -73, 8, -106, -61, 62, 92, -35, 72, 78, 70, 49, -41, 60, 49, -13, -88, 111, -105, -15, -51, 113, -78, 54, 89, 32, -127, -61, -23, -103, -127, -78, 27, -55, -9, 107, -21, 106, -104, -36, -3, -20, -11, -88, -36, 60, -90, -75, -29, -33, -88, -18, -15, 41, -39, 0, 16, -115, 114, 88, -79, 116, 91, -57, -121, -118, -109, -14, -37, -66, -108, -70, -16, -66, -87, -70, -11, 53, -126, -40, 45, -107, 109, 70, 108, -121, -22, 123, 36, -124, 94, -62, -52, -57, -1, 23, 52, 107, 68, 92, 123, -35, 52, -79, -107, 68, 69, -47, -51, 56, 46, -36, 119, -94, 16, -115, -3, -124, 86, 115, -8, -30, 38, -103, 65, 114, 81, -12, 6, -68, -78, 117, -37, 113, 97, -107, -36, 54, 45, -124, 35, -77, 16, 56, -29, 100, 66, -111, 38, 16, -24, 93, -30, -122, 27, -106, -78, 23, 49, 43, -105, -11, -66, 85, -114, -73, -37, 118, 107, 41, 38, 3, -6, -24, -109, 92, 27, 37, 37, 31, 6, 126, 71, -20, 29, 75, 96, 127, 67, 46, 120, -29, -39, -10, -64, -108, 60, 80, -99, 21, -43, 36, 92, 55, -91, -10, 119, -49, 24, -32, -112, 48, 11, -110, -43, -101, 101, -107, -65, 17, 90, -3, 43, -90, -54, -9, -92, 46, -23, -69, -124, -18, -17, 33, 39, 86, -91, -113, 127, -89, -85, 122, -98, -19, 96, -37, 64, -80, -66, 94, 52, -22, -98, 21, 68, 20, -81, -79, -29, 56, -120, -46, -14, 49, -116, 55, -51, -27, 110, -34, 39, 118, -36, 16, 125, -87, -121, -18, -71, 72, -67, 67, -67, -119, -44, -40, 69, 62, 18, -83, -10, -36, -80, -41, 107, 108, -117, -78, -126, 48, 69, 45, -55, 110, -91, 0, 52, -111, 6, -74, -16, 60, 29, 88, -79, -71, -56, 33, -126, -94, 47, 40, -113, 66, -18, 50, 126, 40, 70, 64, 96, 106, 41, -27, -33, -77, 27, -74, -102, 46, -5, 76, 124, 12, 21, 72, 43, -78, 3, -63, 69, -127, 43, 48, 104, 49, -126, 125, 118, -17, -71, -77, -72, 70, 4, 104, 54, -115, 23, -91, -64, 125, -64, -117, 36, 28, 9, -106, 103, -39, 16, -47, 45, 60, -24, -20, 22, 56, -98, -10, 69, 93, -104, 5, 125, -90, -107, 75, -4, -37, -90, 117, -57, 116, -46, -58, -105, -91, 114, -44, -42, 115, -91, -65, -125, 19, -45, 78, -83, 90, -63, 58, 52, 53, -86, -3, -115, -92, -111, -102, -81, -52, -97, -62, -59, 29, 59, -61, 9, -17, 30, -18, 106, -53, 42, 35, 96, 25, -123, 16, -91, -107, 33, 118, -94, 55, -76, -49, -79, 8, 33, -18, 49, 8, 90, 108, 44, -69, -101, 78, 98, -24, 69, 9, -45, 84, 45, -52, 55, -20, 84, 59, 69, -84, 5, 67, 78, 124, -52, -32, 6, 13, 28, 122, -80, 98, -70, 50, -64, 80, -46, 91, -16, 70, 121, 23, -43, -87, -86, 23, 126, -88, 0, 41, -29, 69, 8, -81, -65, 93, 52, 81, 76, 121, -116, 34, -85, 27, 67, -76, -17, -29, 6, 103, -62, -79, -104, -87, -41, -14, -49, -83, -75, -126, -30, 90, -52, 108, -123, 5, -63, -8, -50, -54, -105, -112, -27, -77, 61, 28, 42, -47, 119, -97, 88, -94, 8, -29, 77, 85, -128, 92, 42, -43, -74, -75, 86, 123, -128, 13, 22, 88, 91, 3, 17, -78, 10, 29, 8, 29, -123, 66, -39, 60, -5, -64, 27, -58, -49, 98, 81, -63, -121, -82, 85, -27, -120, 96, 68, -39, -65, 1, -7, 78, 106, 1, 15, 48, 66, 108, 100, 113, 85, 113, 17, -52, 45, 0, -60, 53, 117, -15, -117, -98, -35, 117, 33, 81, -94, -57, -31, -61, 82, 36, -53, -102, 28, 62, -80, -123, -41, 32, 4, -57, -112, -127, -7, 93, -87, 91, -46, -45, -43, -99, 74, 5, 127, -13, 29, -53, -55, 32, 11, -15, -79, 118, -18, -11, -28, 68, -86, -18, -10, -103, -49, 58, -55, -26, 103, -64, -81, 37, 74, -84, 36, 66, 46, -84, -75, 19, -33, 22, 72, -73, -2, -127, 17, 53, -117, -110, -22, -30, 113, 65, 60, 45, -89, -46, 47, -55, 73, 71, -57, -62, -122, 124, 40, -55, -65, 0, 80, 46, 112, 15, -15, 112, -94, 46, -54, -120, -34, 122, -44, -95, 4, -14, -124, 101, 76, 108, -70, 0, -126, 29, -1, -2, 39, 120, 13, 73, 46, -101, -31, -34, 28, -74, -117, -21, 46, 28, -74, 84, -45, 32, 94, -113, -109, 103, 121, -93, -78, 107, 42, -4, 71, -118, -54, -73, -18, -98, 1, -116, 87, 6, -50, -59, 93, -1, 15, 4, -110, -68, 124, -60, 125, -4, -18, -35, -42, -86, 13, -115, 107, 105, 51, -100, 59, 16, -118, -127, -44, 103, 108, -30, 13, -23, -72, 43, 99, 89, -1, 17, 2, -14, -64, 43, -118, -69, 39, 41, -44, -2, -86, 18, -9, 73, -3, -89, -102, -5, 27, 91, 21, -7, 91, 80, 41, 95, -79, -53, -2, 74, 109, 54, -63, -52, 92, -61, -89, -108, -108, 17, -85, -4, 111, -51, 64, 86, -111, -55, 80, 7, -122, -51, 61, -98, -24, 1, -74, -49, -49, -25, 0, -32, -106, 53, -68, -44, 90, -123, -35, 10, -61, -46, -46, -45, -86, -39, 86, 5, -72, -53, 69, -93, 103, 64, -49, 14, -15, 34, -44, -115, -28, -101, -99, -30, 39, -31, -44, 13, 58, -2, -119, 75, 86, 113, -121, -65, 120, 109, 49, 36, 29, 97, 11, 79, -120, -17, -8, -65, -38, 42, -98, 107, 73, -55, -50, 4, -114, 112, 61, 100, -75, 84, -53, 78, -48, 68, 47, -71, 33, 59, -23, 45, 86, 115, -50, -20, -48, 3, 89, -94, -87, -30, 66, -125, 91, -54, -119, -44, -34, 92, 65, 61, -83, -77, 38, -97, 98, -26, 113, 127, -60, 118, 113, 58, 24, -102, -31, -65, -43, -48, 9, 66, 92, 7, 44, 54, 45, -83, 1, -79, -123, 73, 51, 80, 94, -96, -106, 126, 119, 126, -102, -79, 96, -126, -53, -13, -53, 9, 1, -109, 25, -99, -106, -46, 100, -28, -29, -92, -15, -56, -91, 24, 14, 112, 13, 122, 82, -96, 63, -66, -53, 31, 21, 113, 47, 14, 85, -109, 53, -110, 125, -44, 2, 81, -106, -23, 110, -51, 86, -42, 67, -93, -30, -8, -2, -7, 3, -73, -113, 64, -119, 1, 64, -42, -74, -124, -80, -40, -32, 95, 24, -56, 16, 80, 102, 19, -106, 94, 110, -128, 65, -20, 19, -84, 0, -119, -95, -78, 78, -54, -116, -46, -39, 88, 23, 49, -69, -65, -50, 4, -121, 66, 95, -15, -25, -45, -48, 72, -22, -103, 60, -20, 16, -86, -23, -13, -57, -6, -34, -45, 57, -13, -40, 55, -57, -30, -59, -5, -47, -47, 19, -30, 10, 32, -1, -70, -92, -13, -6, -99, -103, -114, -45, 22, 102, -107, -75, 115, -52, -56, -44, -86, -75, -124, -75, -31, 29, -92, 86, 53, 115, 104, -100, 104, -94, -68, 96, -39, -69, 84, 55, -123, 49, 70, 43, 117, 98, -15, 74, -20, 88, -113, 82, -67, 62, 92, -78, 1, 12, 34, 34, -3, -80, 6, 28, 59, 49, 80, -100, -128, 8, 35, 3, -56, 72, -65, 62, -30, 94, -30, -124, -78, -102, 95, 17, 34, 16, 80, -46, 88, 78, 111, -94, -21, 71, -24, 101, 105, -30, -116, 80, -127, -91, -126, 97, -25, 95, -35, 2, -115, 2, 82, 89, -78, -92, 122, -68, 97, 78, 96, 109, 125, -44, 32, 65, -98, -88, -45, -111, 24, 36, 67, 126, -92, -6, -123, 125, -80, 74, -38, -97, 20, -102, 13, 71, 123, 84, 18, -69, -81, -127, 114, 124, -102, 37, -53, -118, -121, 72, 7, 28, 104, -70, -14, -53, -47, 116, -81, 34, -117, 48, 0, -52, 104, -33, -39, 115, -41, -10, 58, -31, -33, -41, -68, -38, -119, -39, -24, 96, -18, 78, -55, -119, 111, 118, -124, 65, 71, 18, 92, -125, -89, -67, 33, -40, -68, -112, -113, 96, -8, 49, -27, -22, -21, -26, 24, 126, 40, 69, 9, 44, -83, -63, 43, 99, 32, 81, -89, 88, 90, -57, -18, 87, -33, -63, 81, 117, -10, 82, -124, -95, 70, 54, 104, 42, 102, -38, 55, -79, -2, 89, -76, -4, 85, 125, -38, -68, 56, 93, -78, 120, 10, -29, 100, -110, 102, -40, -16, 86, 84, -85, -85, -104, -40, 49, -61, 9, -94, -117, -117, -58, -4, -70, -115, 57, -53, -52, 72, -6, 104, -47, -34, 97, 102, -90, -113, 35, -13, 23, 3, -41, 22, 51, 10, 15, -20, -74, 22, 79, -43, 45, -125, -97, 42, 3, -59, 28, 65, 28, -121, -27, -57, -84, 63, -54, -10, -70, 55, -88, -89, 106, -49, -49, 53, -49, -117, 33, 62, -38, 5, 70, -16, -108, -114, -10, 22, -95, 100, -30, -110, -65, -64, 79, 43, -10, -96, 105, 84, -79, 38, -15, 68, 106, -43, 122, -64, -99, 115, -123, 85, -110, 58, 14, -44, 31, 108, 36, -91, 45, -79, -22, 106, -98, 102, -9, -74, 6, 64, 97, -8, -70, -61, -109, 126, 116, 28, 37, 86, -57, 53, -92, -110, -30, 101, 97, 4, -47, 85, -110, 115, 68, 31, -20, -10, -57, 80, -118, 10, -54, -27, 122, -125, 4, 41, 36, -116, 71, -21, -124, 86, -104, 34, -45, -32, -102, -20, -56, 26, -9, 71, 47, -99, -95, -86, 36, -43, 8, 121, -127, -59, -3, -79, 43, -67, -42, 22, 116, -45, 20, 53, -65, -56, 73, 53, 35, -102, -47, 94, 64, 76, 66, -124, 97, 124, -87, -105, -91, -37, -90, -117, -106, -42, -12, -48, 46, 37, -108, 80, 44, -21, -36, 81, -83, -64, 23, -65, -107, 9, 107, 36, 43, 81, 66, 95, -91, 121, -70, -92, -5, -114, 116, -83, -106, 24, -70, 23, 110, 86, -34, 76, 41, 42, 98, -43, -84, -80, -8, 7, -99, -33, -77, 36, -88, 8, -29, 3, 94, -61, -26, 20, 17, 6, -38, 38, 126, 22, -83, 14, -42, 51, -66, 82, 22, -47, 21, -99, -97, 114, -88, 1, 121, -127, 104, -115, 114, -41, 111, 61, -115, 106, 15, -118, 80, -50, 70, 23, 84, 28, -75, -115, 105, -90, 48, -92, -119, 106, -12, -9, -56, -34, -63, 45, 120, 3, 6, 4, -104, -24, -41, 68, 103, -65, -25, -99, 64, -43, 47, 88, -37, 80, -36, -69, 121, -60, 95, -125, 22, -85, -118, 23, 43, -11, -51, 29, -19, 75, 37, -83, 53, -2, 98, -18, 127, -73, -52, -83, -108, -67, -23, 57, 45, -8, 113, -85, -61, -41, -92, 41, -120, -118, 39, -63, -22, -10, 95, -2, 22, -54, 109, 52, -29, -88, 85, 83, -78, -10, -53, 95, -30, 106, -4, -34, 108, -16, 25, 94, -32, -71, 103, 38, -114, -71, -53, 82, -59, 112, -93, -19, -1, -25, 11, -82, -101, -1, 55, 110, 99, 106, 14, -101, 45, 63, 80, 91, -32, -91, -22, -56, 107, -104, 113, -89, -86, 45, -80, -20, 88, -5, 96, -99, -38, -2, 108, -126, 85, 109, -90, 124, 55, -98, 88, 40, -105, -42, 64, -39, 84, 43, -122, -36, -40, -26, -75, 56, 54, -14, 43, -84, 103, -110, 43, 44, -76, -50, 62, 75, -7, 109, -126, 12, -23, -51, 54, 22, -46, -85, -107, 44, -76, 80, -4, 47, 52, -67, -69, 54, -45, -81, 64, -1, 47, -40, 49, 67, -51, -33, -62, -82, 104, 120, -94, 35, -79, 13, -103, 4, 71, -57, -78, 98, -99, -106, -81, 80, 113, 19, 29, -48, 29, 40, -40, 123, -12, 110, -41, -38, -31, -34, -104, 112, -54, -40, -8, 8, -69, 80, 125, 120, 93, 95, 91, 18, -109, 114, -69, 102, -89, 127, -89, 8, -73, 103, 31, -47, -116, -44, 90, 5, 88, -2, -21, 121, -42, -75, -72, -9, -102, -64, 19, 68, -2, -5, -75, 110, -121, 11, 96, -86, 126, 119, -28, 20, -49, -121, -110, -110, 102, -128, -9, -120, -104, 88, -115, 46, 33, -83, -58, -104, -17, -120, 94, 115, 42, 78, -70, -72, 90, 72, 83, 12, -26, 77, 115, 41, -41, -109, -86, -84, -62, -17, -68, -56, 69, -100, -15, 101, 78, -53, -124, 95, 121, 89, -93, -21, -98, 40, -53, -81, 95, 5, 120, -86, -98, 108, -27, 54, 95, -115, 3, 88, -4, -84, -97, -119, -77, -100, -128, -32, -118, -6, -86, 102, 79, 121, -124, 121, -20, 39, -37, 126, -21, 2, 30, 2, 118, -80, -101, -11, 96, -93, 111, -88, -82, 19, 24, -98, -125, -125, 12, 75, 57, 109, 74, -14, -41, -71, -106, 67, -47, 67, 27, -109, 10, 13, 93, 49, 63, -1, -48, -74, 79, -123, -79, 87, 47, -112, 62, 7, 89, 62, -9, 30, 119, 39, 13, -85, -41, -8, 82, -116, 45, 104, -64, -112, -33, 106, -71, 21, -69, -120, -123, 80, -103, 8, -5, -121, 75, 37, 36, 109, 20, 49, 19, -40, -63, 124, -39, -96, -23, 126, -2, -97, 113, 7, 42, 73, 98, 3, 23, 66, -117, 111, -22, 37, 34, -18, -57, 11, -121, 106, 95, -21, -46, 26, -113, 116, -63, -24, 112, -123, -3, -30, 96, 93, -33, -85, 110, -1, -123, 31, -61, 127, 83, 81, -12, -32, -89, 91, 23, -12, 123, -112, 83, 127, -110, 123, 63, -72, 0, -6, 6, 11, -67, -42, 112, 31, -93, -91, -2, -27, 42, 13, 98, -82, -31, -116, 67, 127, 101, -31, 73, -112, -119, -77, -62, -11, 12, 35, 56, -6, 127, -57, 70, -91, 103, -128, 56, -59, -89, 13, 82, -71, 10, -40, -102, -128, 118, -15, 122, -55, 18, 50, 29, 66, 99, 33, -125, 46, 48, 111, -86, 101, -43, -61, 106, -123, -53, 118, 73, 42, -84, -29, 124, 92, -89, 91, -18, 2, -55, 39, -103, -57, 77, -73, 120, 70, 96, -9, -102, -25, 35, -81, -72, -12, -6, -92, -61, 41, -41, -99, -22, 102, 98, 108, -97, -32, 44, -108, -37, -45, 37, -95, -100, -73, -61, -114, -58, 90, -111, -54, 68, 81, -67, -46, 78, -103, 54, 41, 107, -82, -65, 2, 82, -113, 57, -10, 85, 70, -113, 104, 23, -30, 46, -63, 41, -3, -72, 78, 77, -119, -107, 48, -4, -6, -19, 119, -39, 123, 4, 113, -15, -24, 120, -48, 52, -79, -107, -58, -106, -51, 46, 49, -71, -29, 104, -127, 78, -60, -26, -16, -42, -110, 16, -97, -118, 50, -106, -47, -28, -91, 75, 117, 94, -62, 1, -56, 53, -88, -15, 101, 24, -96, 50, -20, 123, -31, 113, 74, 4, 84, 110, 3, -128, 51, 59, 13, -8, -107, -47, 121, 2, -108, -85, -16, 18, -57, 65, 121, -62, 85, 93, 71, 118, -57, -111, -101, 116, 113, -71, -69, -112, -126, -39, -59, 118, -56, -19, 75, 55, 78, -72, -3, 87, 86, -32, -126, 15, -102, 62, 72, 80, 20, 110, 76, -32, 48, -113, -29, -32, 84, 23, -37, -38, 71, 111, 25, -50, 59, -109, 103, -77, -128, -83, -25, -102, -107, -109, -13, -61, -47, -1, 21, 105, -17, -92, -52, -109, -71, -8, 126, 90, -8, -91, -110, 64, -95, 109, 82, 100, 19, -68, 126, 37, 11, -12, 90, -16, -37, -119, 38, -57, 31, -100, -60, 5, 59, -31, -90, 33, 118, -109, -84, 89, -26, 55, -45, -81, -37, 35, 13, -106, -66, -73, -73, 55, -122, -83, -85, 123, -112, 93, 81, 61, 93, -43, 104, 110, -52, -110, -54, 60, -73, 67, 29, 72, -17, -91, -37, -65, -117, -98, 76, -56, 39, -76, 9, -70, 67, -2, 6, -60, 125, 8, -104, 45, 16, -116, 91, -105, 117, 99, 40, -19, -110, 60, 12, -65, 119, 6, -112, 122, 16, -85, 47, -22, -93, -86, 44, 78, -59, 65, 48, -96, 67, -75, 38, 41, -15, 98, 41, 30, -107, -40, -35, -92, 66, 95, -122, -118, 67, 6, 70, 125, 41, -31, 53, -77, -124, 70, -6, 4, -41, -58, 89, 76, -9, 12, -17, 36, 34, -12, 80, 22, 42, 118, 32, -33, 20, -127, 58, 49, -106, 104, 114, -44, -75, -26, -54, 30, 102, 64, -27, 108, -64, 74, -74, -92, 30, 126, 2, 49, 47, 3, 42, 57, 61, 49, -34, 14, -93, -102, -4, 82, -103, -54, -58, -26, -26, 62, -23, 49, -123, -108, -9, 92, -92, 4, 116, -59, 93, 13, 105, 11, -92, 58, -71, 23, 84, 101, 82, -56, -94, 19, -110, 48, 120, -50, -78, 106, 43, 28, -19, 36, 111, 35, -15, -3, 62, -49, 32, 15, 10, 77, -55, 11, -116, -35, -112, -25, 26, 35, -59, -9, 22, 68, 123, -113, 122, 47, 98, -95, 111, -54, 39, -96, 113, 109, -66, -21, 87, 120, 19, 19, -85, 60, 107, -128, 19, 104, -53, 122, -61, -53, 89, -1, -122, -21, 7, -20, 37, 90, 77, 35, 121, 110, -108, -65, -2, 58, -19, -75, -29, -25, 82, 43, 105, 49, 40, 19, -89, -59, -46, 55, 56, 54, 17, -128, 89, -109, 77, 4, 47, -59, -121, 36, -124, -97, -4, 116, -41, 53, 16, 82, -126, -2, -16, -40, -7, -78, -30, -26, -57, 40, -80, 125, -104, 114, -44, -103, -49, -97, -118, 74, 105, -91, 11, -93, -63, -86, 8, 114, -7, 118, -11, 72, 57, -78, -92, 118, -29, 58, 69, 73, 116, -61, 6, -48, 43, -116, 37, -3, 4, 80, 99, -75, -31, 122, -63, 5, 84, 115, 1, 5, 97, -117, -73, 94, 119, 80, -42, 96, -114, 5, 34, -102, -72, -47, 109, 124, -49, 14, -113, -97, -62, 93, -115, 32, 21, -123, 103, -3, 38, -26, 18, 109, -100, -9, -73, -9, -40, -95, 55, 12, -34, -2, -62, -16, 102, -31, -122, -18, 15, 14, -2, 13, 60, 52, 99, -89, 72, -126, -71, 76, -53, 55, 46, 75, -107, -107, -32, 82, -48, 45, -56, 29, 121, 33, 127, 111, -71, 52, 35, -121, 7, -14, -89, -109, 97, -98, 60, 66, -21, -119, -121, 38, -63, -12, -37, 0, -100, 18, -40, -26, -103, -56, -14, -57, 69, -118, -54, -67, 120, -5, 91, 4, 116, -116, -16, -94, 87, 4, -31, -35, -85, -42, 84, -60, 67, -41, 87, 70, -27, -76, 89, -44, 77, 125, -39, 39, 38, -93, -89, -59, -97, 66, -125, -99, 112, -77, -117, -112, -28, 88, 121, -124, -73, -72, -32, -46, 86, -115, -75, -43, -22, -61, 18, -87, 97, 52, 98, 45, 95, -20, 41, 50, -8, -95, -42, 69, 53, 90, -59, -126, 56, 85, -85, -111, 66, 36, -49, 75, -54, 75, 39, 34, -94, -88, -86, 73, -74, 48, 113, -124, 80, 51, 89, 51, -70, -37, -56, 27, -88, -28, -50, 28, 14, -50, -88, 102, 48, -41, -25, -93, 102, -2, 126, 66, 1, 75, 114, 46, -98, -56, 65, -37, 116, 113, 107, -96, -24, 79, 90, 78, 13, 76, -71, -24, 125, -8, 83, -41, 12, -18, -89, -61, -64, -17, -85, -107, 26, -39, 63, -110, 65, -123, -51, 54, 111, 56, -2, 68, 30, -45, 2, 126, -88, -122, -63, 86, -5, -125, 75, 47, -80, -49, -24, 64, -42, 79, -17, -82, -62, 0, -77, -29, 67, 100, -75, -67, -44, -120, 4, -100, -53, -51, -37, 17, 118, -28, 70, 22, 98, 125, -89, -53, 82, -78, 44, -74, 95, 4, -79, 100, 55, 124, 121, -122, 97, -111, 55, 10, 34, 29, -91, 63, 123, -17, 0, -37, -72, -58, -123, 101, -51, 74, 18, -47, -116, 57, 56, -12, 1, 73, -93, 14, -8, 63, 1, 20, -112, -81, 69, 116, -108, -61, -64, 25, 49, -80, -102, 42, -101, -7, 100, -90, -48, 125, 21, -69, 29, -105, 125, -99, -88, -62, -40, -16, -112, -49, -73, 38, -127, 2, -29, 70, -103, -122, -93, 36, 28, -47, -26, -63, 103, -122, 66, -119, -85, 53, 69, 42, -86, -54, -78, -86, -8, -45, 75, -127, 46, -51, 57, 52, -121, 21, 4, 53, -118, 54, -113, -103, 22, 106, 38, 43, -75, 101, 14, 60, -39, -50, 75, 19, 126, -88, 86, -41, 47, 22, -101, 120, 47, -119, -46, 60, -74, -125, 84, 38, -61, -107, -98, 125, 92, 37, -83, 44, -50, 48, -52, 114, 34, -58, -99, 78, 112, -116, 119, -29, 44, -115, -60, -78, -52, -73, -72, -122, -31, 57, -75, 123, 102, -76, 126, -77, 4, 90, -115, -57, 89, 20, 91, 52, -24, 49, 53, -47, -83, 91, 53, 60, 91, 23, 74, -39, -73, 5, -64, 37, -105, 91, 114, -9, 94, 75, -30, -8, -61, -103, 16, -108, -52, 24, -97, -122, -37, 91, -119, -93, -13, 62, 46, -68, -126, -83, 49, 21, 51, 119, 58, 59, -3, 82, 82, 13, 9, -10, 99, -36, -76, -99, 94, -125, 117, -124, 48, -126, 48, 112, 62, -50, -104, 40, 46, 75, -13, -22, -33, 111, -50, 51, 75, 19, -75, -42, 73, 56, -97, 90, -10, 84, 47, -68, -85, -70, -14, 46, 7, -81, 56, -28, -11, -12, -67, 2, 61, -125, -126, 88, 115, -2, 106, 38, 125, 78, -3, 36, 22, 101, -88, -4, -94, -5, -2, -54, -11, -35, -16, 74, 26, -127, 86, 90, 124, 19, -57, 20, 111, 62, 43, -104, -109, 31, -59, 113, 26, 57, 45, -8, 115, 125, 104, -12, 24, 122, 126, 59, 60, -96, 121, -12, -44, -32, -94, -6, -11, -75, 52, -49, 80, 47, -62, -96, -88, 114, -92, -126, -81, -74, -100, 89, 40, 97, -43, -47, 22, -114, 59, 123, -76, 11, 25, 83, -21, -6, -76, 126, 61, -9, -76, -40, -49, 38, -119, -1, -53, -127, 3, -85, -111, 94, -1, -44, 90, -125, -39, 30, 25, -70, 40, -79, 95, 93, -95, -3, 96, -78, 83, 18, -104, -99, -19, 24, -94, 45, -88, 104, -13, 100, -106, 30, -126, 12, 81, 31, 118, -24, -80, -75, 101, -67, -49, -6, 89, -23, 122, -105, -109, -50, 103, -126, -11, -59, 117, -22, 101, 39, 14, 20, 50, -84, -72, -99, -115, 102, 85, -92, 41, 95, 99, -28, -73, -44, -26, 0, 100, 127, 54, 37, 67, 100, -43, -3, -54, -98, -21, 43, -35, -87, -62, -25, 47, -48, 87, 7, 64, 55, -101, -93, -19, -73, -49, 102, -21, 59, -13, -3, 31, -7, -116, 68, 57, -36, -4, 95, -79, 6, -23, 102, -61, -60, -70, -118, 87, 75, 2, -46, 22, 109, 67, -24, -60, 64, -40, -120, 73, 87, -41, -8, 9, 92, -84, -17, 44, -113, 117, 84, -49, -37, -52, 78, 31, -18, 82, -11, 123, -24, -17, 47, 49, 97, 62, 124, 55, -93, -18, 78, 117, -72, -127, -72, -103, 125, -110, -111, 83, -105, 87, 103, 67, -97, 112, -64, -122, 47, 48, -120, 82, 62, -97, 71, 82, -96, 111, -68, -9, -42, 7, 26, -40, 102, 57, 68, 84, 108, 5, -2, -5, -35, -116, -12, -63, -9, 107, 29, -84, -28, -32, 92, -115, 50, -107, 102, 58, -4, 99, 82, -66, 84, -22, 67, -35, 126, -55, -53, -62, -38, -93, -24, -103, -26, 50, 46, -61, -66, 104, -39, 33, -120, 62, -59, 36, 73, 121, -91, -50, -44, -85, 20, -87, 51, -127, 55, -68, -4, -67, 104, -103, 113, 111, 109, 110, -76, -43, -59, 32, -7, -14, -117, -128, 100, -128, 22, -92, 59, -85, 119, 2, -19, -21, 7, -54, 5, -93, 80, 19, -67, 88, -22, -79, -87, -103, 50, 86, 40, -11, 99, -78, 106, 11, 108, 6, 6, -104, 37, -50, 99, 124, -45, 104, 69, 102, 97, 32, 80, 54, 27, 90, 66, -33, 37, 50, -29, 90, 82, 62, -87, 121, -120, 83, 33, 30, 59, -28, -18, -116, -4, -73, -65, -28, -16, 99, 26, -23, 116, 109, -108, 90, 77, -58, 123, 99, -81, 54, -80, -87, 33, 101, 91, -22, 8, 4, -23, -92, 45, 63, -73, 37, -105, -115, -75, -93, 113, 12, -63, -90, -45, -70, -100, 119, 105, 27, 64, 40, -6, 74, -11, 93, 105, 58, -117, 25, 69, 96, -72, 9, 60, 47, -79, -12, -100, 96, 43, 55, 99, 15, 119, -68, 113, 35, 44, -10, 27, 91, -66, 89, -63, 81, -62, 34, -10, 33, 21, 74, 111, 88, 3, 121, -90, -89, 21, -1, 83, 12, -43, -91, 99, -94, 124, -122, -19, 46, -102, 27, -64, -74, -91, -39, -110, -118, -117, 48, 121, -43, 71, -29, 106, 49, 31, 18, 86, 116, 43, -109, -78, 21, -103, 68, 56, 111, -60, -57, -29, 19, 13, -55, 65, 4, -58, -82, 20, -35, -43, -30, 121, 10, -60, 118, 58, 76, 82, 32, 70, -127, 98, -55, -93, -81, 108, 79, 13, 60, -68, 83, -21, 46, -55, -2, 41, 96, 68, 127, -102, 6, -105, 104, -110, -5, -71, -83, 101, -84, -111, 39, 33, -107, -55, -78, 114, 68, 106, 20, -118, 66, -46, -121, 77, -92, 2, 115, 2, -116, 80, -13, 21, -73, 101, -121, -126, -7, 24, 71, 103, 27, 23, -83, 47, -5, 125, 5, 123, 72, -18, -106, 57, 44, -51, 100, 118, -115, 71, -35, 98, -33, 71, -9, 52, -19, 20, 107, 6, 52, -60, 8, -25, -11, 118, 117, 83, 92, -34, -52, 91, -18, -84, 120, -4, 7, 10, 99, 95, 43, -120, -109, 119, 88, -40, 19, -21, 38, -42, -112, 10, 6, -17, -8, -82, 50, 113, -3, 68, -98, 92, -109, -9, 115, 112, -105, 24, 102, -47, -4, -96, -124, 120, -43, -57, -85, 71, -26, 112, -14, -105, -70, 5, 36, -7, -108, -91, 52, -118, -116, -127, -13, 55, -36, -107, -111, 118, -111, -55, -50, -33, -111, -110, 24, 91, -122, -94, 10, -128, 84, -26, 65, -72, 93, -116, 26, 7, -53, 64, 66, -71, -85, -8, 42, -108, -62, 1, 19, -94, 105, -92, 91, 119, -61, -74, -122, 122, -32, 52, 101, 59, -24, -66, 103, 21, -114, 124, 17, -9, 93, -123, -88, 1, 69, 124, 13, -60, 91, -90, 53, -36, 23, -51, 126, 92, 109, -50, 65, 32, -68, -66, 86, 111, -126, 92, 33, -68, -94, -116, 25, -42, -120, 80, -48, -50, -1, 87, -19, -114, -18, 2, -67, -45, -97, 56, 32, -1, -78, 86, -113, 23, 73, -29, -40, -102, -110, 101, 12, -55, 38, 4, 85, -88, -112, -98, 119, -3, -65, 42, 23, 2, 8, 13, 3, 57, 6, 85, 21, 108, 84, -110, 48, -90, 98, -70, 54, 42, 69, 125, -13, -42, -109, -7, -98, 31, 77, 39, 71, -40, 30, 3, 53, 39, -116, 106, 76, -44, -95, -11, 85, 13, 4, 25, 52, -88, -96, -113, 69, 121, -5, 99, 114, -96, -58, -111, 91, 71, 95, 78, -100, 67, 93, -99, -88, 0, 41, 75, 107, -126, 20, 89, -11, 100, -120, 82, -80, -30, 117, 116, -41, -2, 95, 64, 16, 103, 68, -53, -17, -122, 93, 25, -19, 78, 78, -96, -45, -95, 117, 107, -41, 36, 22, 18, 49, 98, -79, -74, 61, 11, 79, -104, 21, -79, 64, -71, 40, 107, 17, 118, -97, 36, 108, -109, -30, -91, 32, -6, -122, 30, 53, -65, 53, -111, -115, 115, -83, 76, 99, 62, -63, 68, 1, 34, 80, 36, -78, -43, -60, -59, 69, -94, 32, 67, -2, -43, -2, -51, 1, -42, -48, 123, 54, 114, -31, 30, -31, 24, -29, -43, -61, 12, 93, -49, 55, 12, -121, 59, -114, -72, 110, -102, 66, -3, 48, -98, 65, 100, 43, 92, 22, -87, 6, 70, 83, 98, 77, 111, -73, -79, -14, 107, 40, 80, 90, 44, -56, 65, -93, -120, -34, -22, 114, -7, 94, 103, 121, 94, 104, -94, 97, 34, 74, -27, -111, -68, -91, -2, 82, 105, -34, 54, 114, 102, -18, 10, -100, -81, 106, 61, 7, 49, 93, -94, 113, -36, -25, -126, 87, -104, -36, 80, -46, -76, 86, 41, -105, -43, 34, 68, -72, 105, 110, -17, 21, -60, 72, -40, -96, 53, 73, -26, -1, 13, 121, -24, -12, 8, -89, -34, 94, -6, 79, -126, 82, -13, 58, 110, 44, -101, -41, 25, -96, -91, 42, 110, 3, -56, -25, -53, 114, -4, 51, 70, 0, 16, 22, 16, -10, 48, 123, 2, 51, -113, 36, -79, 52, -32, -7, 47, -93, 49, 44, -21, -55, 95, -95, -108, 40, 58, -96, -97, -79, 12, -80, -107, -97, 74, 76, 38, -43, 116, -105, 96, 32, 26, 73, -93, 112, 2, -128, 24, 66, 105, -16, 88, 40, 25, -26, -11, -86, -60, 112, -50, -75, 34, -40, 52, -45, 13, -122, 118, 2, -123, 108, 88, 77, 114, -124, -104, -19, -39, -121, -74, -88, -4, -44, 85, -85, -36, 114, 34, -94, 121, -1, -54, 99, 108, 70, 56, -46, 85, -86, 104, 4, -95, 119, 95, -24, 90, 77, 127, 20, 98, -53, 70, -47, -115, 44, -3, -43, -21, 33, -128, -38, 48, 1, -66, 122, -94, 50, -86, -25, 83, -16, -74, -19, 17, -74, 46, -45, 17, 121, -46, -62, 9, -94, -26, 0, -42, -77, 17, -80, -11, 112, 43, 91, -110, 23, 87, 20, 108, -37, -58, -58, 69, 105, 90, 17, 19, -40, 2, -3, 3, -48, 87, -127, -43, -8, 57, -48, 50, 115, 0, -63, 11, -5, 5, 38, 118, 69, -14, -99, -66, -27, -43, -14, 48, -116, 35, 5, -90, -63, -78, 15, -80, -36, -100, 47, 112, -48, -76, 28, -77, 96, -28, -46, 14, -57, 3, -39, 101, 89, 81, -80, 114, -20, 35, -35, 64, -120, -118, -22, -31, 112, -43, 101, 109, 88, 22, 65, 107, 107, 11, 31, 65, -127, -99, -107, 36, 8, 30, -45, 58, 41, 23, 78, -107, 24, -12, 88, -93, 98, 100, -37, 122, -77, 24, 104, 74, 14, -86, -73, -38, -27, -2, 38, -61, 14, -10, -48, -8, 32, -70, -116, 22, 83, -64, 2, 31, -128, 26, -1, -42, -9, -86, -87, -113, -42, -47, -15, -96, -42, 70, -74, -8, -11, 30, 34, -15, -70, -86, 121, -56, -114, -83, 117, 85, 97, -33, 76, 46, 57, 57, -68, -25, -122, -59, -127, 91, 17, 115, 0, 66, 119, -11, 115, 66, 1, -20, -51, -82, -16, 13, 18, 72, 66, 120, -69, 49, -34, -52, -78, 9, -77, 41, -91, 101, -69, -76, -43, -105, 87, 36, -35, -93, 111, 105, -36, 6, 47, -65, 124, 65, -48, -54, -76, 21, 105, 0, -23, -71, 73, -68, 28, -1, 78, 5, 116, -114, 59, 54, 15, -62, -83, -73, -58, 125, 32, -41, 79, 9, 45, -51, -37, 123, -92, 44, 125, 57, -9, -13, 64, 52, -21, -37, -3, 114, -25, -16, 58, -86, 76, -80, -70, -88, -6, 75, 120, 123, -88, 117, -127, -107, 1, -110, -25, 92, 105, 17, -28, 9, -2, -80, 121, -83, 112, -38, 10, 77, -80, 35, 123, -65, 95, 8, 39, -42, 114, 95, 82, 34, -115, -14, 85, 95, -34, 99, 75, -106, 47, -84, 15, 67, 11, -4, 80, -68, 80, 37, 3, 89, 49, -27, 72, -105, 104, 114, -72, -83, -98, -22, 28, 119, -98, -40, -68, 51, 52, 25, 89, -72, -6, -25, 53, 102, -85, 121, 3, -1, 94, 22, 21, -3, -1, 35, 1, 126, 74, 17, 120, -82, -72, -114, -45, -17, 2, 73, -17, -38, -32, 14, -45, 79, -14, -100, 120, 72, -52, -8, 90, -61, 64, -116, 92, -82, 35, -96, 25, -89, -11, 44, -72, -81, 46, 14, 13, -51, 85, -2, 33, 0, 108, 111, -60, 107, -108, 27, -67, 118, -123, 66, -60, -4, 76, 112, 0, -5, -55, -25, -57, -95, -77, 93, 73, -67, -61, 24, 26, -94, 118, -120, 66, 53, 98, 52, 33, 25, 71, -87, 19, 10, 80, 60, 75, -1, 21, -10, 89, 7, 90, 78, -36, -102, 41, -91, 78, -69, -81, 25, 49, -100, -48, -114, 106, 40, -114, -79, 67, 11, 116, 48, 4, -71, 28, 60, -125, -12, -127, 6, 112, -75, -14, -100, 6, -67, 68, -77, 2, 32, -28, -96, -90, 92, -92, 74, -58, 113, -18, -75, 125, -78, -52, -18, -26, -2, -89, -51, 103, -18, 111, 1, -11, -112, -72, -91, -43, 61, 81, -86, 98, -50, -70, 28, -127, -34, 114, -67, -123, 9, -108, 4, -43, 75, -81, 118, 21, 78, -42, -82, -35, 54, -125, -112, 50, -35, 126, -79, 86, -89, 0, 15, -111, 121, 28, -88, 105, -88, 46, -36, 106, 17, -74, -1, -26, 119, 124, -56, -42, 7, -122, -33, -84, 37, 119, -72, 7, 61, -16, 115, -19, -108, -36, -91, 74, 61, -30, -19, 16, 40, 119, 28, 91, -77, -100, 90, 26, -67, -66, 9, -69, -57, 98, 63, 47, -89, 110, 18, 32, -96, -91, 37, 113, 51, 117, 66, -115, 95, 30, -34, 95, -126, 60, 92, -79, 119, -128, 77, -73, 79, 8, 90, 0, 87, -17, -68, 95, -73, 34, 103, -102, -84, -73, 90, 114, 59, 114, 26, 79, 41, -89, -68, 102, -122, -1, 27, 103, -29, 30, -13, 121, -97, -103, 78, 35, 52, 51, 12, -90, 17, -102, -96, 110, -63, 73, 74, 88, 114, 97, 5, 90, 0, -23, -43, -12, -71, -46, -20, 38, 101, -84, 104, -78, -71, -23, 82, -94, 119, 58, 75, 10, 13, -120, 60, -112, -68, -93, -38, 3, -66, 13, 50, 124, -13, 84, 4, -101, -91, 75, -70, 53, -40, 81, 69, -70, -9, -97, 114, -99, -20, 41, -60, -42, 21, -105, -79, -64, -67, -105, 116, -109, 73, -16, -29, -44, -67, -119, -47, 46, -6, -113, -74, 80, 3, 75, 24, -85, 63, 100, 104, 21, -4, -1, 77, 83, -120, -65, -101, 21, 34, -19, 81, 55, 19, -29, 66, 15, -40, -11, 107, -122, -87, -29, 26, -89, -69, 61, -5, -49, 87, 83, 79, 92, -67, 25, 118, 74, 1, -93, -122, -92, -118, 110, 29, 125, -25, 11, 84, 102, 94, -87, -83, 87, 47, -16, -93, 56, 0, 37, -42, 124, -112, 81, 46, -122, 127, -109, -53, 127, -53, 57, -125, -20, 27, 92, 36, -78, 69, -45, -99, 77, -88, 99, -113, 68, -57, 49, 31, -102, 47, -31, -112, -60, 70, 110, 14, 74, -2, -116, -69, 26, -76, 88, -106, 116, -9, -71, 88, 36, 126, 51, 34, -82, 64, -7, -33, 114, 41, -94, -55, 58, -57, 72, 124, -6, -52, 98, -67, -47, 65, 112, 72, 74, 89, 65, -110, -82, 57, 104, 27, -3, 99, 87, -56, 23, -104, -27, -26, 75, 107, 71, 99, -57, -20, -125, -68, 19, 91, -93, 113, -93, 60, -19, 28, 31, -16, 109, -108, 87, 12, -15, -44, 0, 97, 85, -122, -104, 25, 56, 121, -10, -25, 111, 78, 84, 45, 70, 4, -18, 118, 63, -51, -116, 91, -19, 62, -73, -106, 84, 76, -93, -93, 22, 83, 95, -61, -57, 44, -67, -88, -98, 11, -72, -74, 104, 11, -70, 65, -63, -124, 57, -54, 87, -27, 80, 126, -81, 56, -97, 120, -102, -104, 126, -34, 24, -13, -89, -22, 113, -79, 97, -92, -80, 115, 121, -126, 59, 1, -68, 81, 50, 47, -112, 125, -68, -59, 17, 44, -3, -67, 71, 88, -104, 35, 92, -64, 109, 126, 112, -59, 94, -84, -89, 105, -98, 51, -72, 45, 1, 55, 3, 96, 125, -2, 72, -22, 122, 114, -48, -2, -115, 41, -100, 39, 65, -86, -20, -89, -91, 30, -21, 122, -16, -89, 15, -121, -66, 83, 108, 112, 60, -28, 1, 26, -108, -13, 95, 123, 18, 39, -104, 49, -27, -24, -39, -45, 85, 72, 73, 26, -45, -44, -61, 49, -32, 6, 15, 0, 30, -110, -116, -63, -23, 42, -91, 86, -120, 9, 43, 47, 32, 76, 110, -51, -116, 19, -73, -42, 24, -16, 5, -89, -112, 20, 126, -1, 46, 90, -13, -120, -116, 26, -122, 53, 84, -43, -23, -80, 9, 122, 119, -112, -34, -37, -90, 41, -113, -75, 31, -8, -39, 40, -24, -3, 71, -9, 119, -42, -33, 68, 82, 83, 33, 36, -39, -53, 53, 113, 97, -128, -35, -122, 97, 113, 71, -85, -81, -1, 93, 105, 65, -126, -96, 84, 25, 105, -4, -9, -26, 101, -99, -55, 55, -10, -104, 119, -4, 102, -8, -121, 70, -109, -96, -22, -68, -8, -48, -20, -51, 122, -11, -117, -65, 117, -8, -55, -2, 78, 27, 25, 108, -19, 56, 13, -106, -128, 90, 47, -126, 89, 115, -26, 4, 63, 73, 25, 53, -58, -118, -38, -53, -76, 31, -32, 65, 62, -34, 17, 39, -21, 19, 77, 109, -19, 124, 68, -103, -49, -78, -30, -3, 22, -118, 67, 20, 14, 115, -42, -123, 57, -126, -110, -71, 83, 83, 88, -36, 127, -70, -62, -19, -14, 35, 91, -103, 116, 31, -19, 116, -20, -49, -25, 78, -71, 119, 51, 52, 101, -34, 76, -80, 88, 17, 9, -118, -110, -7, -115, 89, 96, -70, 88, 81, -116, -89, -2, -15, 124, 11, 103, -39, -72, 31, 60, -83, 118, 114, 14, -59, -2, 19, -7, -29, -75, 127, 49, -56, -77, -39, 49, 18, 96, -67, 79, 69, -32, 9, -88, 92, -121, -88, 50, -97, -1, -43, 13, -8, 114, -28, 97, 14, -33, -87, 69, -85, -58, -45, -30, -61, 75, 74, 31, -4, 68, 122, 108, 107, -25, -20, -98, -76, 118, -49, -5, -72, 89, -113, -41, 2, -40, -39, -79, 23, 90, -26, -116, 95, 51, 0, -55, -56, 88, 124, -66, 34, -80, 94, -14, 51, 5, -30, -84, 123, -116, 115, 67, -83, 111, 108, 124, 38, 18, -65, 84, -103, 81, -38, 68, 1, 72, 35, 45, 27, -103, -109, -74, 10, 1, -95, -127, -115, -124, -18, 94, -33, -46, 14, 107, -65, 44, 5, -45, -123, -52, -81, -30, 33, 43, -60, 15, -81, -97, 22, 14, -16, 91, -99, 25, -91, -35, -127, -95, 87, 23, -27, -69, -37, -64, -83, 83, 56, -41, -122, 85, -57, -15, -69, 114, 87, -21, 100, 67, 7, -25, 69, 122, 111, 42, 45, -97, -118, -38, -74, 93, 7, -53, 59, -105, -113, 30, -25, 124, -111, 38, -121, -22, -45, -91, 122, -87, -29, -7, 27, 116, -68, 99, 93, 8, 19, -110, 12, 87, 93, 2, -23, -54, 101, 125, -69, 52, 15, -125, -52, 52, -97, -121, -102, 106, -124, 36, -20, -24, -61, 93, 74, -58, -47, 95, -70, 122, -104, -41, -127, -115, 51, 102, 78, 66, -113, -27, 126, 87, -91, 103, 125, -102, 5, 85, 37, 59, 83, -21, -95, 100, 96, -75, -22, -90, 44, -102, -20, 72, 1, 4, 127, -42, -33, 103, -87, 28, 89, 38, -40, 120, 124, -82, 78, 61, -20, -125, -60, -32, 23, 95, 106, -26, -90, -72, -124, -11, 67, 40, 122, -36, 60, 94, -73, 64, 110, -37, -82, 56, -112, 28, -35, 106, -44, 94, 116, 93, -79, -123, 114, -61, 16, 2, 75, 77, -67, -49, 75, -114, 110, 99, 123, 101, 79, 67, 9, 2, -51, 124, -115, 75, 12, -127, -93, -46, -34, -104, -111, 54, 44, 111, -12, 94, 99, 43, 91, -65, -50, 54, -96, 76, -11, 25, -31, -91, -117, -36, 56, 61, -112, 7, 57, 77, -20, -89, -124, -100, -66, -30, 2, 99, 5, -63, -111, -82, -44, 113, -97, -12, -21, -55, -74, -60, -119, 29, 22, -60, -96, -41, -2, 29, -22, -25, 22, 75, 52, -62, -76, 3, -31, 73, 111, 9, 85, 24, 25, -128, -59, 23, 75, 20, -9, 111, -23, 43, 53, -75, 99, 41, 95, -93, -68, -76, -78, -50, -95, 2, 106, 51, 94, -117, -35, -115, 81, 43, -128, -9, 108, -89, -52, 42, -18, -81, -9, 87, 19, -95, -110, -124, -5, -19, 28, -58, 67, -123, -83, 42, 15, -53, -49, 55, 3, 34, 44, 114, 100, -81, 104, 2, 9, 88, 80, 95, -68, -31, -95, 27, 94, 8, -62, -89, -94, -73, -57, -8, -27, -25, -26, -37, -97, 24, 78, -21, 102, -74, 83, -95, -113, -41, -59, -15, 17, 53, 56, -33, -6, -118, 117, 98, -115, 82, -20, -100, -64, 109, 28, -99, 119, -114, -114, 20, 58, 88, -46, -33, 110, 32, 70, 126, 127, -54, 58, 46, 107, -107, 109, -34, -106, 76, 64, 84, 103, -48, -86, -40, 66, -125, -91, 36, 6, -96, 66, 66, -44, 109, -31, 78, 125, -114, -69, -40, 125, 117, -110, 114, -108, -97, 27, 4, 33, -23, 84, 61, 40, 58, 24, 9, 8, 67, -79, 99, -47, 56, -113, -58, 104, 59, -14, -19, 127, 41, -91, 45, -121, -111, -19, -33, 24, 91, -86, 91, 11, 89, 61, -58, 106, -48, -56, -34, 102, -86, 82, 6, 57, -73, 61, -77, -54, -13, 20, 102, -87, 55, -23, -49, -60, 23, 108, 27, -44, 48, 21, 127, -64, 12, -79, 72, -78, -88, 96, -85, -29, -77, -20, 112, -30, 17, -37, -40, 111, -95, -6, 108, 105, -85, 119, 122, -94, -117, 35, 37, -8, 46, 47, 13, -28, -4, -104, -109, -34, 114, -7, -80, 90, -67, 33, 31, 99, 80, 92, 95, -116, 117, -90, 68, -82, 6, 64, 17, -87, 9, 12, -12, -120, -35, -119, -52, -37, 103, -74, 29, -115, -78, -17, 13, 14, 84, -2, 102, 95, 120, -122, -23, -59, -42, -3, -68, -32, -51, 57, -39, 124, 11, 48, 32, -74, -71, -13, -91, 115, 19, 50, 28, -127, -86, -60, 96, 40, -80, 97, -115, 6, 86, 36, -117, 126, 94, -66, -56, 85, 38, 22, -86, 111, 88, 59, 40, -53, -16, -30, -87, -39, 80, 57, -75, 85, 61, 13, 70, 39, -69, 115, 92, -80, -3, -23, 37, 70, -111, 96, 31, -27, -56, 34, 72, 41, -67, -96, 46, -1, 23, -53, 121, 14, 84, -103, 20, 79, -34, -123, 115, 58, 13, 34, -107, 88, 105, -56, 115, -114, 10, 127, 87, 81, -106, 103, -80, -86, 127, 90, 115, 98, -22, -34, -30, -102, 26, 71, -90, 88, 17, -81, 48, 57, 60, 84, 22, -63, 39, -19, -5, 50, -92, -7, -20, 127, -58, 113, -128, -71, 83, -110, 92, -71, -21, -21, -112, -36, 33, 79, -73, -8, -124, -97, -41, 0, 71, -88, 23, 122, -46, 116, -61, -52, -117, -123, -93, -49, 113, 58, -45, 79, -122, 72, -73, 105, 117, -5, -121, 55, 19, 24, 5, 17, 9, 8, -117, 75, -118, 76, 3, 15, 62, 116, 39, 46, -104, 122, -94, 2, 75, 68, -21, -51, -18, -5, -15, 126, -100, -65, -11, 70, 123, 60, 21, 125, -48, 46, -68, -11, 43, 125, 51, 18, -127, 59, -27, -73, -67, 54, -122, 95, -73, 47, 110, 48, -28, 109, -107, 49, -25, -57, 83, 54, -92, 75, 124, -19, -115, -99, -82, -31, 67, 127, 55, -10, -71, 27, -1, 23, 86, 67, -107, 104, -70, 52, 50, 109, 66, 79, -71, -51, 101, 59, 24, 81, -23, -34, -58, -62, -56, -38, -127, 81, -23, 95, -103, 127, -68, -28, -96, -15, -35, 9, -124, -88, 73, 91, -122, -73, -66, 93, 122, 47, -100, -36, -53, 79, 112, -24, 22, 85, -36, 118, -46, -43, 109, -46, 75, 108, 55, 97, 125, -100, 25, 76, 53, 116, 50, 37, -22, 25, 54, -35, -11, -100, 59, 51, 45, -44, -125, -95, 39, 21, 18, -61, -110, -80, 2, -67, 112, -16, 1, -109, -118, 42, 50, -107, -115, -35, -110, -1, -121, -98, -42, -60, -90, -34, -71, -42, 102, -104, -55, -12, -65, 93, 39, -59, -18, 49, 24, 104, -118, -108, -95, -38, -14, 67, -11, -22, -75, 64, 125, 29, 25, 52, 31, 112, -122, 86, 114, -46, -13, 65, 62, -7, -103, 62, -112, -25, -114, 38, 88, -93, 59, 101, 3, -107, -99, 54, -22, 109, -86, 77, 114, -101, -30, -128, 82, -69, -79, 17, -69, -67, 90, -28, 34, 19, 43, 50, -36, -10, 122, -40, -25, 16, -14, 88, 96, -89, -60, 95, -99, -19, 59, 51, -43, -110, -17, 57, -28, 93, 3, 102, 37, 46, 69, 103, 110, 6, -116, -101, 106, 103, -15, 66, 19, -112, -38, -35, -46, 24, 73, -106, 53, 38, 35, 109, -71, 119, 15, 22, 71, 15, -106, 63, -43, 25, -60, 109, -84, -99, -17, -46, 122, 117, -43, -48, -10, 25, -102, -119, -12, -11, -51, 66, 103, 72, -14, -119, 51, -89, 47, 93, -81, -75, 14, 75, 80, -115, 34, 98, 23, -38, 89, 47, 47, 118, 101, -112, -89, 73, 34, -42, -23, -59, 35, 60, 67, 66, -110, 127, -11, -101, 77, -65, -30, -127, 95, 42, 58, -22, 90, 39, 9, -30, 72, -95, 81, -67, 33, -53, -9, -17, 112, -95, 8, -18, 75, 34, -81, 95, 96, 57, -53, 12, 50, 50, 111, 41, -126, -34, 71, -1, -29, -99, -95, -128, 12, -110, 113, 122, 80, 104, 15, 96, 13, 104, -119, 77, 0, 125, 95, -54, 31, 3, -29, -61, 72, -113, 11, -53, -100, 94, 30, 14, -42, -20, -78, 23, 83, 90, -63, 113, -32, 50, -91, 120, 19, -104, 88, -51, -61, 74, -79, 93, -74, 113, 15, -80, -119, -58, -87, 86, 54, -66, -79, 50, -13, -100, -128, -93, 61, -73, 88, -59, 108, 111, -7, 68, 52, -34, 45, -113, -9, -69, 13, 41, -62, 1, 77, -80, 103, 58, 23, 112, -69, 22, 101, 60, 5, -44, -71, -85, 49, 60, -115, -28, -23, -83, -93, 23, -76, 121, 45, 24, 84, -91, -15, -125, 102, -72, 105, -126, -103, -18, 107, -119, -98, -19, -64, 72, -26, -104, -28, 4, 4, 41, 108, 127, 82, -91, -23, 116, 71, -67, 112, 114, 47, 32, 105, -15, 98, -106, 101, -67, 11, 11, 6, 10, -126, -72, -74, -108, 68, 28, -41, -84, 35, 103, -102, -1, -110, -104, -24, -71, 0, 16, -40, 85, 33, 108, -32, -80, -51, 79, 85, 115, -53, 20, -66, -68, -105, 69, 119, 37, 9, 116, -45, 12, 38, -99, -121, -17, -3, -63, -74, -50, -59, 50, -88, -16, -63, 98, -112, -120, 83, 63, 37, -42, -97, -77, -67, -83, -5, -56, -94, -49, -16, 98, 72, 21, -11, 118, -79, 97, 87, -40, 43, -121, -26, 60, 7, -24, 60, -97, 41, 113, -127, -25, 79, -125, -94, -5, -119, -39, 66, 118, 124, -23, -39, -116, 63, -76, 127, 85, 93, 61, 111, 53, 18, -84, 108, -86, -61, 105, 47, 102, -14, 3, -39, -110, -117, -43, -27, -78, 30, -88, -76, -126, -88, 15, 93, 48, -58, 44, 110, -86, 85, 45, 117, -24, 82, 28, 118, 66, 100, 83, -67, 24, 92, -122, -60, 96, 4, 60, 88, 88, -83, 90, 76, -53, -79, -4, 88, -63, -22, -65, -66, 40, 91, 101, 90, -54, 85, -30, 92, -51, -38, -83, -110, -67, 2, 116, -120, -55, 21, -78, -87, -61, -58, -42, -56, 17, 22, 77, 26, -90, -32, 89, 58, 95, -2, 85, -103, -120, 88, -15, 32, -110, 60, 75, -15, -2, -2, 117, 48, -41, -78, -4, 95, 113, -41, 30, -122, 117, 73, 4, 63, -49, -79, -67, -115, -96, 33, 65, -59, 6, 65, -121, 95, -7, -120, -61, 101, -83, 12, 47, 48, -113, -115, 8, -72, -80, 32, 80, -83, 101, -59, -97, 116, -32, -100, 123, 86, -18, 20, 20, 91, -33, 72, -40, 14, 48, -108, 15, -92, 63, -41, -9, 30, -80, -22, 2, 60, -120, 25, -50, 38, 79, 11, -28, -103, -53, 84, 98, 121, 119, -22, 112, -119, 44, -19, -121, -2, 33, 23, 47, 107, -71, 38, 86, -51, -62, -36, -73, -71, 19, 85, -42, -66, -34, -100, -71, 82, 24, 67, -9, 94, 51, 77, 77, 0, -108, 11, -50, -36, -20, 21, 8, 69, -45, 106, 18, -118, -75, -57, -41, -25, 62, 65, -12, -79, -21, 44, 45, -31, -16, 8, -75, 51, 61, -51, -52, -9, 75, 116, -106, -127, -56, -81, 36, -49, 36, -59, -108, -99, 46, 45, -54, -60, -15, -83, -128, -120, -25, -120, 126, -86, -16, 115, -46, 31, 51, -36, -88, -62, -78, -9, 26, -56, 111, -6, -72, 72, -12, 72, -126, -93, -111, 63, 80, 117, -126, 54, -123, 37, -92, -10, 34, 13, 69, -53, 104, 71, -94, -21, 55, 1, -33, 48, 71, 79, 95, 52, -35, -114, -107, 22, -125, 22, -97, 39, -28, -58, -88, -22, -29, 63, -58, 89, 103, 28, -22, -89, -119, -124, -109, -113, -40, -90, 105, 66, -44, 86, -76, -116, 39, 106, 42, 2, 59, 49, -48, -46, -41, -65, 43, 59, -98, 2, -52, 21, 108, 35, 89, -11, 102, 45, 83, 47, 48, 14, 60, -97, -39, 24, 57, -65, -76, 24, 51, -65, -106, -40, 68, 56, -8, -9, -62, 60, 94, 40, -5, 106, 60, -90, -13, -29, 2, 79, -76, -18, -74, -39, 98, -62, 67, -38, -71, -120, 69, -15, 5, -85, 5, 103, 25, -18, -39, 78, -93, 56, 24, -68, -93, -18, -116, -91, -3, 54, 38, 91, 94, 29, -99, 65, -4, -12, 17, 40, 75, 126, -55, 87, -20, 38, -95, 26, -91, 3, 91, -55, -77, -104, 115, -54, -34, -115, 66, 71, 123, -83, 84, -73, -53, 86, -104, -98, -54, -60, 25, -69, 27, -24, 107, 57, 49, -30, 6, -82, -108, -19, 26, 61, 86, 120, -114, -80, 99, -76, 4, 70, 29, 37, -123, -38, -68, -49, 21, 86, -104, -122, 106, -9, -55, -82, 39, 105, -13, -66, 72, -107, -120, 56, 121, 34, 67, 73, -24, 48, -24, -89, 15, 75, 51, -92, -81, 29, -100, -59, 44, -69, -42, -68, 46, -98, -77, 2, 126, 105, 70, 10, -63, -5, -40, -32, 63, -120, 94, -61, -5, 69, -123, 70, 13, -60, 54, 126, 31, -66, -70, -81, 126, -92, -5, -43, -8, -126, -25, -6, -115, 44, 116, -50, -50, -91, 98, -81, 3, 46, -3, -79, 120, 35, -56, 71, -94, -67, -56, -22, 87, -122, 0, 62, 117, 54, 71, -116, -36, -40, -71, -125, -24, 82, 69, -122, -113, -51, 15, 118, 13, 66, 17, 88, -7, -32, 80, 113, -90, -91, 88, -57, -87, 32, -100, -47, 9, 20, 68, 36, 93, 56, -117, -32, -81, 111, -127, 84, -31, -46, 56, 81, 94, 36, 77, 92, -110, 118, -77, -70, 90, -32, 123, -21, 83, -115, -113, -115, 54, 85, -74, 70, 60, -20, 77, 75, 91, -25, 20, -83, -121, -25, 39, -119, -42, -22, 53, -70, -86, -92, 97, 14, 67, 78, -118, 52, -4, 98, -117, 67, -17, -88, -47, 99, -47, -7, 6, -126, 77, -104, -46, -66, 77, -1, -126, 94, -14, 45, -2, 60, 79, 119, -9, -83, 66, 60, -34, -32, 61, 2, -127, -126, -8, 66, 114, 28, 87, 72, -127, 56, -107, -5, -37, -79, 20, -49, 57, -5, 17, -24, -126, 54, 80, 114, 18, -105, 27, -77, 26, -14, -61, -80, 123, -37, 23, -51, -21, 5, 7, 27, 34, -80, -83, 126, -23, 55, -107, 46, -86, -7, -72, -2, 40, 85, -83, 2, -55, -52, 38, 98, 44, -18, -17, 56, -25, 2, -50, -10, -59, 68, -105, -128, 45, -50, -23, -95, 78, 121, -111, 27, 103, 13, -2, 126, -71, 31, -36, 59, -28, 73, 3, -26, 73, 112, 96, -23, -23, -83, 18, -35, -54, -41, -53, 122, 13, 51, 82, -28, 49, 121, 59, -98, 110, 3, 25, -86, -31, -20, 56, 58, 74, 1, -88, 64, -24, 75, 48, 124, 112, 44, -21, 20, -1, 97, 15, -41, 94, -60, -60, 123, -61, 64, -24, 98, 90, 61, -109, 48, -61, -35, -126, -29, -128, -69, -51, 93, 25, 46, -61, 39, -80, -36, -69, 33, -79, 93, -4, -82, -107, 29, -102, 123, -108, 126, -42, -103, -70, -111, -4, -84, -21, 71, -108, 78, -13, -95, -71, 51, 73, 39, 70, -100, -21, 27, 125, 113, -125, -110, 109, 112, 86, 53, 91, 9, 36, 97, 53, 83, -81, -2, -101, 8, 13, 13, 77, -32, 45, -105, -68, -76, 4, -71, -82, 92, 8, 55, -37, -109, -19, 29, 77, 88, 16, 48, 19, -27, -111, -40, 67, -99, 44, 26, 53, -122, 40, 113, 57, -120, 87, 109, -41, 114, -9, 46, 58, -59, 19, -112, -73, 118, 74, -80, 10, 75, 15, 1, -120, -14, 117, 73, -77, -3, -104, 51, 119, 58, -31, -110, 12, -101, 95, 66, -20, 46, -9, -30, 12, -36, -22, 21, 0, 75, -101, 86, -107, 73, 45, 94, 21, -27, -3, 60, -71, -110, 14, 70, 42, -70, -20, -53, -128, 85, 31, 60, -105, 117, -92, -101, -120, 87, -39, 34, 20, 125, -1, 13, -13, 118, -105, 26, 76, -30, 89, -86, -122, -46, -16, 87, -46, 16, 86, -23, -105, 125, -52, -73, 35, -72, -26, 24, 48, 116, -59, 97, 107, -60, 14, 41, -110, 51, -61, -10, 7, -106, 67, -26, 70, 72, 73, 53, 29, -76, -108, 52, 61, 9, 6, 116, -26, 114, -8, 53, -71, 1, -56, -15, 44, 94, 87, 42, 98, -73, -17, 127, 29, -48, 2, 54, 123, 118, 41, -46, 31, 93, -107, 79, 105, 59, 5, -95, -53, 45, -19, -90, 13, 124, -51, -79, 60, -78, 63, -90, -118, -45, 28, -76, 95, 81, 110, 8, -120, -59, -122, 108, -29, -112, 25, -35, 64, -93, -33, -27, -5, -81, 123, 120, -10, 8, -102, -2, 120, 19, -32, -50, -3, 119, -4, -98, -34, -21, -65, -15, 71, -23, 45, -25, 0, 73, -52, -27, 13, -78, 53, -99, 46, 89, -49, -18, -25, -13, -76, 76, -14, 122, 57, 25, 90, -9, -21, 11, 21, -86, -71, -2, 111, -60, 49, -83, 2, -93, -31, -45, -107, 107, -2, -23, 12, 87, -35, 110, 114, 11, 49, 100, 122, 66, 39, 84, 16, 51, 123, -16, -47, -88, 17, 68, 83, -112, 102, -30, -112, -107, 39, -37, -96, -121, 0, -93, -82, 68, 13, -99, -64, -6, -30, -80, 116, 57, -105, 121, 57, 11, 71, -112, 33, 16, -65, -58, -44, 56, 125, 47, 27, -107, -3, -14, -27, 1, -13, -95, 76, -57, 110, 72, 23, 42, -12, -3, 98, -26, 93, 98, -9, -79, 17, -90, -33, 108, -25, 27, 66, -107, 76, -14, 113, 86, 47, 77, 61, -79, 89, -78, 104, 67, 72, 14, 73, 16, 16, -39, 73, 54, 83, -54, -87, 46, 29, -90, -95, 94, 81, 81, 51, 8, 116, -59, 21, -94, -33, -102, -66, -53, -51, -36, 1, -75, -12, -63, -15, -14, -128, 78, -36, 57, -73, -16, -84, -105, 54, 5, -51, 104, 73, -52, 70, -17, 53, 66, -91, -67, 27, -61, -118, 26, -46, 40, -35, 119, 31, -29, -118, -45, -11, -32, -73, 37, 112, 15, 19, -123, -59, -61, 32, 29, -77, -29, 127, 32, 27, 121, -109, 62, 113, 23, 119, -53, -110, -1, -44, -9, 50, 30, 10, -52, -84, -105, 12, -57, 73, 125, -113, 127, -120, 118, 92, -11, 79, 20, 117, -51, -106, 110, -35, 125, 85, 55, 72, 42, -86, -122, 9, 106, 123, 37, 87, 27, -83, 12, -103, 68, 105, 61, -76, -123, -67, 84, -81, 59, -35, -109, 76, 19, -26, -97, 122, -109, -46, -119, -104, -106, -17, 99, 64, 49, 101, 18, -17, -50, 63, 112, -11, -21, -121, 12, -116, 106, 65, 126, 72, -9, 15, 46, -78, 122, -114, 8, -38, -94, -93, -45, -23, 85, 1, 113, 111, -99, 69, -110, -61, -128, -20, 106, 106, -22, -105, -53, -32, 21, 119, 98, 64, 95, 82, -123, -2, -64, 0, 68, 67, -31, -72, -16, 42, 73, -19, -21, 4, 7, -127, -92, 102, -20, -125, 113, 30, 89, 80, -91, 49, -39, 35, -55, -41, -21, -83, -58, 14, -114, 85, -5, 9, -60, -120, 113, 117, 89, 103, -33, 65, 113, 94, 60, -84, 30, -80, -101, 61, 102, -35, 117, -92, -21, -103, -11, -120, -107, 81, 72, 101, 21, 22, 113, -101, 93, 55, 95, 0, -17, 37, -112, 72, -71, 92, 17, -113, -9, 50, -66, -58, -95, -122, -1, -107, 22, 17, -86, -119, 28, -79, 23, 90, 47, 33, 126, -30, 120, 124, 124, -73, -55, 25, -88, 69, -95, -102, -34, 111, -40, 42, -24, -39, 18, -44, 61, -56, 52, -11, 45, 73, -71, 73, -119, -12, -84, 32, -105, -53, -74, -25, 86, -87, -66, 88, -12, 70, -37, 24, 40, 112, 58, -85, 65, -101, 98, 17, -72, -73, 57, 89, -34, 105, -58, 3, -92, 52, -79, 60, 15, 57, -116, -102, 62, 48, -40, 14, -55, -51, 113, -116, 64, 97, 54, -35, -94, 35, -73, 99, -24, -84, -42, -44, 11, 17, -9, -22, 73, 7, 47, -92, 73, -102, -1, 55, -31, 100, -97, -69, 30, 87, 85, -25, -1, 117, -34, -117, -62, -58, 48, -56, 1, 27, -125, -119, -39, 61, 70, -106, 96, 84, 16, 43, -56, -64, -10, -85, 61, 93, 88, 56, 20, 15, 73, 26, -112, 31, 4, -75, -88, 69, -97, -62, -30, -77, -82, 79, -122, -104, -81, 59, 25, -102, -48, 80, -94, -65, -75, -13, -13, -125, 48, -86, -67, -21, -10, -67, 54, 5, 27, 95, 4, 49, -42, 125, -93, 29, 109, -80, 75, -72, 110, -102, 33, 17, 64, 13, -116, 27, 46, 44, -66, -117, -40, -72, -45, 86, 23, -103, 38, -73, -61, -88, -74, 122, -36, 50, -84, -1, -83, -32, 63, 119, -39, 120, 34, -55, 39, -106, 54, 102, -48, -47, 78, 122, 79, -60, -44, -97, 116, -124, 71, -3, 17, 47, 65, 116, 101, -1, -107, 61, -67, -71, -32, 12, 58, 25, -39, -34, 99, -68, -16, 23, 17, -14, 126, 97, -38, 38, 87, -37, 86, 44, -98, -44, -19, 11, -5, -71, -98, 70, -84, 38, -63, 107, 91, 116, 49, 59, -92, -61, 83, -82, -61, -86, -111, -27, 17, 46, -43, -45, 60, -88, -11, -31, 53, 126, 18, 47, -58, 30, 32, -111, 32, -117, 57, 103, 9, 121, -43, -75, -70, -15, 43, -56, -95, -110, 14, 72, -31, 65, 51, -44, -19, 108, 59, -54, -38, -80, -73, 53, 92, 16, -2, 107, 97, -44, -82, -71, 75, -59, -1, -104, -101, -77, 80, -4, -124, -49, -79, -45, 121, 127, 44, 39, 29, -67, -102, -106, -88, 111, 1, 92, -53, 66, -114, -82, -86, -128, -75, -86, -3, 48, -78, -88, -109, -32, 41, -74, 1, -28, -120, 92, 31, -65, 114, 114, -102, 121, -123, 28, 62, 72, 98, 50, 126, 91, -6, -17, -24, 8, 51, 66, -36, 126, -123, 107, -65, 82, -95, -85, 81, 53, 110, 117, 99, 0, -12, 1, 102, 48, 77, 124, -22, 28, -42, 43, 117, 7, 39, -64, -78, 35, 87, -43, -68, -122, -31, -101, 13, 73, 54, -18, 49, -52, -78, -53, 73, 92, -23, 51, -53, -14, -78, 124, -68, -35, -123, 119, -119, -15, 109, -44, -99, -6, 104, 79, -44, 36, -12, -11, -63, 22, 58, 56, 85, -86, 64, -51, -85, 86, -14, -65, -118, -112, 51, -119, -25, -86, 87, -25, 105, -2, 79, -40, 100, 99, 58, 36, -114, -29, 114, 77, -84, 88, 13, -27, 38, 124, 31, -27, 46, -91, -27, 124, 37, 15, 116, 118, -30, 43, 16, -73, 56, -96, -14, -56, -119, -3, -39, 15, 100, 45, -97, -7, 112, 53, -24, -8, -20, -71, -67, 97, -32, -62, 98, -37, 69, 109, -83, -39, 18, -71, 122, 9, -93, -9, -34, 93, -36, 107, 13, 20, -32, -23, -75, 55, -81, -78, -119, 93, -127, 21, 94, 4, -45, 45, -58, -44, -30, 42, 49, 40, 89, -107, 73, 117, 100, -32, -92, 105, -92, 43, -9, 109, -35, 61, 79, -29, 30, 76, -14, 56, 73, -97, -53, -68, -75, -17, 25, 37, 78, -102, -39, 79, -13, -65, 100, -12, -110, 93, -59, -88, -74, -117, 114, 53, 99, 59, -125, 23, -108, -26, 80, -74, -39, -72, 50, 87, -10, -109, 40, 34, 84, 60, -102, -53, -34, -19, -45, 69, -29, -70, -3, 84, -100, 34, 19, 27, -109, 1, 102, 114, 107, -121, -43, 34, -71, -91, 4, 81, 64, -54, -34, -61, 57, -3, 47, 42, 77, -77, 101, -22, 39, 34, -93, -32, -82, -68, 54, 50, -10, 4, -116, 79, 125, -41, -104, -5, -75, 121, -100, 83, 81, -70, 72, -48, 48, 48, -33, 94, -90, 44, -94, -100, -71, -23, 118, -88, 79, -44, 46, 93, -2, 22, 107, -34, 127, 73, -108, 111, -100, -111, 42, -116, 37, -81, -58, -34, 44, -2, 2, -32, 119, -71, 10, -72, 125, 112, -77, -53, 20, -122, 54, -88, -30, -56, 23, 60, -111, 81, -69, 28, 114, -31, 53, 117, 30, 46, 117, -39, -61, 46, -57, -112, 97, -27, -100, 118, -18, 55, 92, -7, 22, 41, -88, 57, -64, -10, 77, -55, -70, -47, 82, -89, 32, 119, 3, -7, -13, -112, -34, 72, -112, 58, 56, 126, -115, 61, -77, 105, -122, 93, -111, 116, 117, 93, 4, 88, 29, -29, 71, -100, 57, 43, -60, -22, 25, 73, 96, -125, -69, -35, -44, 61, 107, -41, -53, -128, -47, 104, 25, -7, -104, 43, 57, -27, -112, -63, -42, 50, 62, 38, 119, 88, -67, -125, -122, 41, 63, 108, -28, 16, -19, -94, 10, 75, 56, 50, -13, -86, 46, -3, 97, 18, 74, 52, 127, -8, -20, -61, 72, 68, 47, -112, 85, 29, 74, -111, 116, -34, 109, -32, -71, -81, 118, -105, 31, -32, -28, -73, -53, 61, -33, -88, 0, 61, -44, -84, -83, -64, -15, 16, -121, 40, 37, 93, -58, -16, -30, -92, -111, -68, 83, 79, -70, -108, 87, -32, -120, 14, 96, 91, -4, 8, -40, 122, -108, 27, 95, -54, 0, 103, 65, 7, -121, -26, 99, -55, 68, -71, 119, 91, 77, -119, -11, 84, 100, 63, -108, 111, -77, 50, 20, -38, -33, -68, 22, 75, 38, -112, 64, -82, -81, 10, -19, 86, -64, 127, 50, 9, 116, 53, -42, -35, -6, 13, -40, 77, 65, 25, -21, 3, 77, 90, 103, -98, 12, -1, -115, -62, -83, -53, -55, 80, -95, 33, 58, -84, 8, -69, 74, -18, 8, -18, -94, 61, 18, -84, -68, -56, -120, 65, 72, -17, -58, 7, -112, -56, 74, 105, -43, -41, 3, 16, 86, -75, 74, -17, 85, -124, 98, -8, -81, 60, -61, 29, -28, -34, 38, -124, -72, 26, -57, 29, 35, 36, 52, -14, -34, 50, 25, -121, 87, -72, -118, 54, -57, -104, -15, 124, 81, -105, 28, 16, -65, 11, 78, -128, 81, 111, 42, 26, -119, -113, -102, 73, 105, 19, -26, 98, -40, 40, 97, 59, 111, -85, 125, -85, -52, -48, -29, -35, 78, -89, 102, -104, 61, 105, -16, 122, 61, 101, 17, -37, -9, -90, 123, 91, -9, 1, -121, 53, 40, 2, 53, 74, 45, -65, -127, -15, -117, -30, -10, -9, -48, -91, 21, 45, 87, 31, 95, 110, -96, -124, 86, 29, 118, 47, -26, -12, -89, 19, 124, -13, -26, 120, 116, 72, 119, -34, -41, -78, 114, 91, 73, -21, -37, -56, 30, 111, -125, -35, 88, 89, 100, -87, 71, -34, 54, -54, -17, 84, 4, -8, -67, 73, -90, -38, 34, -81, -42, 110, -20, -109, -66, -113, 89, -80, 46, -126, -68, 103, 63, -58, -27, -80, -6, 44, 30, 115, 122, 7, 122, -17, 71, -35, 15, -1, 44, 89, 125, 98, 46, 36, 29, -105, -117, 39, 88, 5, -127, -92, -80, 2, 94, 79, 39, -33, 42, 0, 34, -57, -43, -8, -83, 3, 113, 48, -120, 15, -94, 92, -34, 9, 29, -112, -97, -126, 60, -49, 121, 81, 68, 101, -62, 127, -24, -74, -113, 11, -64, 12, -81, -98, -63, 72, 68, 26, -104, -93, -73, -93, -14, 103, 41, 81, -91, 78, 35, 15, -54, 12, -97, -90, 43, -96, -59, -76, -8, 64, -64, 43, 54, -127, -17, -58, -10, -9, -117, 84, -105, -126, 41, 76, 35, 34, -110, 4, 11, -6, -53, -112, -73, -62, -12, -55, 65, 99, -86, 80, 80, -115, 9, -67, 10, -27, -6, 123, 105, -103, 90, -55, -72, 2, -28, 15, 76, -116, 120, -10, 88, 126, -45, 103, 32, 112, 1, -11, 72, -58, -116, 107, -115, -116, -55, 75, 28, 25, -39, 3, 62, -44, 38, -95, 124, -59, 75, 115, 77, -13, -32, -106, 15, -60, -38, 68, 116, -93, 101, -79, -84, -56, 96, 90, -18, 48, 43, 112, 86, -81, -114, -24, 86, 81, 9, -101, -108, -116, -18, -17, 120, 114, -36, 98, 126, -39, -49, -24, -2, 95, 116, 103, 117, -18, -73, 72, 61, -98, 39, -106, 53, -32, 45, -56, 24, -63, -30, -27, -95, 25, -112, 10, 24, 5, -15, -77, -36, 53, 48, -121, 115, -1, -63, -114, 80, -59, -74, -122, 65, 76, 66, 64, -117, 109, -124, 40, 64, 91, -118, 34, -104, -48, 6, 2, -50, 72, 110, 97, 51, 69, 48, 82, -5, -44, 80, -118, 16, 60, 124, 5, -84, 51, 91, 13, -45, 62, -101, -99, 127, 106, -2, -15, 62, 19, 124, 75, 79, 43, 114, -51, -34, -111, 113, -39, -28, -84, 83, -46, -14, 91, 51, -25, 38, -21, -23, -93, -33, 114, 2, -12, -31, 32, 24, 6, 38, -104, 90, -78, 94, -108, 16, -6, -17, -118, 52, -109, -121, -37, 13, 21, -62, 72, 50, 105, 20, 4, -16, -65, 107, -107, 11, 123, 49, -34, -59, 108, -33, 90, 72, 120, -58, 73, 118, 15, 53, -108, 67, -2, -114, 4, -58, 49, -50, -84, -4, -114, 73, -94, -9, 69, -80, -99, -1, -53, -41, 87, 66, 77, -125, 64, 59, -6, 39, 41, 60, 64, 106, 17, -48, -66, -2, 31, 107, 36, -92, 48, -90, 101, -21, 40, 43, 38, -14, -128, -62, 10, -11, -21, -73, 119, -109, 42, 93, 100, 54, -68, 100, -53, -127, -19, 108, -71, 90, 36, 64, 75, 50, -17, 55, -57, -63, -79, -112, -3, 123, 70, 57, -80, 8, -49, -112, 68, -34, -34, -126, 34, 80, 109, 111, -37, 19, -20, -57, 17, 62, -26, 108, -86, -99, -107, -52, -15, 40, -35, -24, 90, -40, 13, -31, 24, -98, 106, -59, -108, -47, -24, -48, -76, 99, 39, -71, -97, -50, 87, 59, -122, -119, -123, 16, 11, 2, -101, 2, 96, -52, -64, 76, -55, 25, -57, -75, -15, 55, 113, -3, -36, 93, -93, 127, 71, 14, -48, 67, 77, -62, 50, 83, 82, 70, 53, 45, 21, -90, -35, -108, 117, -121, 9, 62, -60, 113, 15, -10, 78, 30, 31, 58, 115, 86, -76, -73, 93, -123, 20, 31, -110, -101, -6, -52, -85, 85, -112, 27, 26, -18, 96, 123, -51, 45, -71, 1, -78, 34, -35, 46, -67, 104, 83, 22, 63, 58, 82, -82, 32, -117, -9, 23, 11, 67, -5, 21, -54, -49, -27, -127, 9, 50, -80, 23, -92, -97, -123, -7, 19, -71, -91, -113, -99, 105, 90, -48, -32, -17, -41, 56, 16, -98, -121, -30, -88, 14, 12, 43, 125, -118, -105, -78, 121, -52, 65, -6, -12, 2, 23, -20, 65, 30, 101, 118, 14, -115, 47, -68, 52, 62, 31, 105, 67, -8, 30, 89, 7, -63, -4, -68, -66, -114, -20, 62, -38, -4, 99, -40, 52, -100, 1, 89, -5, -4, 66, -62, 14, 67, 49, -74, -119, 109, 98, -57, 57, 43, 14, -105, -80, -119, -58, 13, 107, 100, -103, -42, -35, 123, -67, 102, -5, -35, 1, -103, -59, 97, 44, 44, -3, 80, -127, 103, -124, -105, -27, 33, -74, -102, -35, 16, -33, 80, 62, -78, 24, 42, -33, -13, -60, -112, -19, -49, 55, -120, 14, -106, -98, -112, -55, -8, -100, 94, 50, -121, -18, 61, 5, 34, -112, -88, -104, 85, 32, -85, 6, 53, -104, -14, -34, -104, 81, -74, -105, 28, 72, 11, 111, -25, -32, -63, 84, 104, 51, -5, -6, -65, -76, -53, -128, -22, 40, -65, 21, -92, -111, 125, 28, 63, 16, -52, -119, -30, -5, -17, 123, -95, -63, -105, -108, -23, -46, -24, 53, -94, 116, -126, 43, -82, -81, 58, 45, 20, -65, 45, -125, -60, 13, 0, 16, 49, -64, -72, -114, -107, 12, -31, 59, -108, 92, 34, 89, 9, 87, 74, -31, -47, -80, -47, -37, -13, 74, 105, 42, -84, 26, 21, 35, 92, -100, 62, -104, -24, 95, -38, 0, 119, 21, 17, -21, -44, 105, -34, 118, -124, 84, -14, 103, 92, -40, -51, 80, -121, 7, -38, -21, 86, 62, -75, 22, 31, 66, -98, -37, 111, -29, -124, -46, 12, -51, -30, -91, -103, -78, 86, -43, -35, 15, -101, -88, 2, -123, 90, -57, 7, 120, -10, -16, -119, 14, -123, 14, -14, -74, -98, -7, 75, -4, 115, -101, 60, 54, -45, 59, -94, 93, -49, 79, -62, 111, -63, -115, -60, -33, 36, 127, 91, 1, -36, -60, -112, 24, 7, 9, -97, 110, 94, 123, -42, -17, -72, 50, -95, 37, 72, -96, -102, -96, 90, -41, 124, -41, 85, -39, -37, -34, -3, -27, 52, 103, -37, 102, -20, 37, 120, -19, -128, -44, -81, 74, 23, -4, -72, -66, 44, -26, -50, -4, 39, -92, 109, 31, -103, -83, -98, 99, 63, 103, 109, 22, -120, -53, 124, -35, -92, 62, -125, 43, 58, -103, -120, 66, 70, -78, -34, 41, -21, 2, -114, 5, 71, 45, 61, -116, 112, 35, 43, -55, -118, -67, -14, 92, -39, -50, 18, 69, 108, 89, 120, 54, -26, -31, -124, 20, 49, -118, 20, -42, -113, -111, -89, 96, 68, -2, 18, 71, -47, -32, -13, -26, -4, -17, -26, -22, -60, 110, -34, 112, 11, -22, 93, 20, -27, -121, 97, 108, 55, -110, 106, 54, -54, -96, -61, 29, -90, -98, -102, 56, -80, -92, 126, -11, 118, 29, -77, -64, -119, -106, -77, -43, 127, -124, -23, 120, 36, -102, 83, 41, 48, -99, 20, -96, 42, -102, -124, -62, 127, -19, -31, -117, -32, -85, 124, -92, -92, -45, -122, 42, -3, -99, 40, 123, 78, -69, -35, -33, -43, 103, -71, -23, 127, 89, -16, -7, -32, 62, 13, 118, -8, 1, -108, 108, 13, -84, -45, -20, 121, 108, -38, -51, 57, -84, 32, -115, 13, 117, 33, -66, 76, 15, 71, 119, -38, -39, -31, 0, 16, 1, -84, 94, -61, -15, -55, 98, -15, 82, -58, 120, 95, -35, 118, -10, -82, 48, 97, 10, -51, -2, 101, -127, -26, 107, -66, 72, 44, -7, -75, -108, -121, -4, 102, 20, -29, -69, 34, -122, 72, 44, -61, -2, 42, 113, 79, -98, -109, 34, -69, -36, -16, -62, -78, -115, 9, -63, -98, 83, 17, -72, -33, -72, -33, -52, -68, 31, -39, -47, 4, 63, -49, -84, 49, 72, 77, 105, -63, 65, 13, 22, 18, 15, -1, 64, 60, -113, -116, 113, 2, -104, 24, -118, 90, -117, -23, 7, -48, -6, -51, -69, -68, -88, 0, -75, -72, -83, 50, 44, 51, -40, -65, -2, -80, -100, -10, -90, -108, 34, 98, -125, 3, -119, -43, 80, 77, -65, 111, 91, 53, -22, 101, -92, 3, -30, -15, 113, -29, -42, 93, -13, -93, 99, 17, -124, -108, 10, -106, -26, 96, 50, -105, -4, -64, -41, -24, 39, -90, 3, -66, -21, -46, 92, 94, 74, -41, -45, -65, -16, 24, -39, -59, -126, -12, 87, 76, 118, -63, -25, 83, -78, 8, 95, 96, -106, -69, -83, 57, 61, -86, 54, -93, 56, -122, -95, 20, -67, 113, 82, -81, -5, -39, -113, 55, 116, 11, -108, 3, -71, 66, -121, 21, 40, -113, -36, 97, -111, 127, 83, -79, 84, 59, -126, -72, -18, 43, 52, -29, -94, -44, 50, -16, 46, -61, -114, -90, 78, -94, 74, 77, -23, 94, 56, 56, -70, 52, -96, -76, -73, -109, -7, -81, -22, 10, 35, 29, 112, 62, 104, 114, -30, -3, 66, 18, 110, -22, 44, 79, -115, 21, -127, -127, 71, 39, -115, -14, -91, -96, 82, 97, -57, -100, 43, -86, -22, -96, 38, 84, 68, -96, 63, 53, -24, 71, 113, 48, -2, 0, 108, 106, -39, 32, -81, 67, 84, 103, 111, 98, 12, 25, -69, -118, 75, -36, 4, 79, -93, 107, -3, -101, -79, -30, -108, 87, 27, 23, -89, -113, 112, 42, 50, -118, 37, 66, -89, 3, -95, -105, 83, -118, -47, 29, -54, 118, 8, -10, 14, -49, 120, -23, 69, -65, -35, 69, 63, 118, -86, 127, -73, -34, 6, -55, 45, -55, 27, 73, -87, 15, 113, 100, -16, -107, 116, -95, 4, -57, 78, 49, 112, -117, 42, -41, 56, -8, -45, -108, -92, 93, 1, 36, -58, 101, 79, 73, -64, 57, -111, -24, -41, -108, -123, -15, 69, -29, 38, 74, 32, 108, 107, 54, 67, -27, 84, 97, 75, 37, -61, -19, -101, 40, 79, -5, 24, -69, 30, 33, -61, -31, -37, -33, 50, 15, -69, -86, -14, 116, -78, 12, -31, -75, -95, 55, 77, 102, 76, 50, -13, 7, -10, -22, -38, -98, 62, -99, 94, 8, -32, 101, -110, -128, -80, -20, -105, 2, 43, 16, 57, -8, -95, 123, 121, -125, -63, -25, 97, -41, 91, 48, 27, 108, 102, 32, -48, -12, -31, 57, 106, 30, -127, 114, -78, -103, -65, -113, -93, -80, 115, -40, 103, 93, -17, -107, 124, 101, 36, -65, -25, 125, -106, -23, 115, -31, 89, -122, -89, -48, 44, 37, -48, -21, -100, -89, -114, -4, 44, -121, -71, 41, -19, 39, -4, -119, -39, 101, 11, 69, -57, -60, 91, 108, -1, -62, 109, 119, 95, -91, -119, 37, 125, 8, 84, -84, 121, 125, -83, 69, -37, 3, -91, 11, -107, 21, -91, -81, 74, 25, -18, -44, -4, -110, 16, 20, 69, -81, -26, 121, 87, -112, 57, 91, -40, 87, 15, 29, 37, 18, -60, 99, 79, 117, 79, 116, 106, -35, 43, 100, -45, -123, 109, -6, 16, 104, 52, 11, -37, 109, -17, -112, -38, -27, -98, -107, 121, -92, 90, -73, 50, 110, -31, 108, 99, 22, -59, -22, 5, 109, 82, 111, 88, 118, -112, 17, 80, 116, 39, -109, -52, 25, 117, 107, -96, -124, -78, -92, 85, 89, -105, -63, -53, 89, -12, 5, 122, -48, -5, 110, -88, 81, -72, 114, 102, -5, 91, 27, 22, -100, -106, -13, -113, -114, -20, 91, 91, -11, -21, -83, -69, 118, -13, 84, 55, -24, -79, 60, -23, -23, 0, -30, -107, 118, -79, -82, 89, -104, -50, 25, -50, -7, 95, -92, 104, 118, 45, 0, 52, -93, -124, -74, 126, -117, -41, 34, 33, 97, 115, -3, 11, 46, -33, -37, 48, 53, -65, -33, 115, 69, 16, -29, -43, 122, -25, -111, -90, -92, 127, 38, 110, 125, 35, 40, -106, 92, -21, 95, 17, -26, 59, 12, 23, -50, -123, 92, 113, 109, -2, -114, -127, -65, 52, 57, 42, 71, -15, -90, 47, 104, 91, -70, 38, -78, -112, -52, -61, -45, -87, 26, -49, 119, -113, -71, -19, -2, -74, -84, -98, -33, -19, 5, 35, 16, 101, -79, 1, -82, -56, 65, 66, 7, 101, -121, 66, -101, -51, 68, -108, -79, 92, 81, 104, 66, -79, 108, 102, 63, 12, -66, 100, -24, -101, -88, -104, -115, 89, 16, 21, 57, 117, -107, 9, -106, 46, 109, -94, 67, 47, 51, 94, -13, 114, 98, 11, -75, 69, -122, -23, -36, 103, 90, 13, -101, 14, -89, 55, 5, -99, -13, -67, 69, 101, 47, 20, -79, -127, 94, -73, -113, 25, 25, -35, 71, -49, 49, -10, 102, 14, 10, -80, -85, 52, 53, 26, -12, -69, 87, 81, 123, 72, 44, 0, 50, 72, 78, 31, 124, -117, 126, 79, -105, -117, 109, 67, -93, 45, -86, -24, 36, -69, 77, -55, -102, -106, 4, 106, -11, -57, -49, -51, -6, 107, -112, -87, 114, -56, 119, 102, 82, 109, -111, -53, -63, -121, -55, -15, 25, -8, -103, -44, 65, 62, 46, 123, -116, 55, -42, -89, 80, 33, 99, 10, -26, 100, 26, 63, 118, -69, 8, -35, -98, 45, -104, 18, 16, -6, -121, 21, -50, 57, -67, 76, -63, -123, 10, 42, 41, 48, -58, -91, -32, -37, 78, -50, 29, 124, -126, 16, 55, 8, 124, -111, 69, 32, -28, 17, -47, 100, 74, -126, 96, -109, 60, 50, -128, -105, 2, -63, -13, 81, 79, 64, -9, 48, 1, 22, -23, 15, -10, 88, -43, -73, -23, 112, 93, 8, 65, -26, 69, 29, -52, -14, -122, 54, -30, 89, -95, -43, 24, -98, 74, -37, -106, 40, 87, 119, 55, -24, 123, 85, -115, -110, -57, 64, 27, 18, 13, 6, -36, -75, -30, 126, 42, -98, -43, 112, -18, -3, -111, -37, -70, 89, -1, 6, 46, 46, 69, -6, -85, 90, -100, 69, -16, 93, -18, 57, -40, -71, 45, -114, -94, 119, 64, -44, -90, -33, 91, -5, 67, -106, 50, 97, -114, 33, -10, 73, 78, -113, -91, 97, -47, -74, -69, -34, 58, -55, -66, -124, -86, -128, 2, -50, 122, 34, 16, -33, 98, 9, 108, -80, 110, -26, -40, 93, -4, -78, -117, 88, -97, 72, -82, 17, 81, -25, -120, -99, -6, -117, 27, -128, 54, 118, -83, -11, -115, -25, 103, -48, 78, -54, -96, -38, -33, 54, 85, 80, -32, -8, -120, 28, -65, -58, 99, -53, 71, -14, 90, 45, 45, -2, 96, -75, 28, 113, -77, 0, 70, -53, 9, 121, 105, 93, -117, 35, 75, -34, 85, 36, 44, -57, 77, -93, 115, -2, -79, 33, -94, 101, 48, -21, -36, 97, -104, -21, 81, 98, -11, -5, -89, -113, -37, 94, -83, 87, 19, 115, 103, 35, 118, 0, 102, 4, -46, -67, -55, 50, -47, 19, 11, -127, -42, -84, 52, 77, 110, 51, 60, -29, 110, 26, 22, -41, 63, -64, 104, -69, 66, -37, 38, 9, -72, -8, -3, 21, -93, -115, -79, -15, 115, -69, -59, -41, 24, -27, 57, 104, -31, -116, -12, 47, -78, 118, -83, 70, -57, -1, 3, 68, -116, 55, -7, -34, 14, 21, 119, -90, 114, -12, -78, -96, 86, -106, -3, -80, -99, -48, 19, -45, 124, 80, -120, 46, 32, -57, -124, -98, 119, -81, 10, -71, -7, 123, 125, -72, -66, -126, 123, 93, -79, 50, 32, 100, 27, 50, 123, 76, 0, -11, 95, 1, 108, -118, -58, 57, -79, -102, -115, 45, 6, -107, 106, 91, 88, -103, -92, 10, 63, -52, 56, 108, -24, -125, 42, -36, 14, 35, 82, -81, -26, 8, -62, 112, -31, -2, 119, 123, -90, -103, -33, -46, -10, -16, 111, 65, -3, 75, -95, -118, -12, 73, -85, -26, -65, -82, 84, 43, 56, -119, 120, 105, -127, 105, 49, 25, -69, -83, -9, 15, -37, -120, 83, 53, -116, 117, 102, 1, 8, -72, 42, 106, -19, 47, -112, -87, 89, -26, -52, -101, 65, -99, -120, 99, -24, 71, -86, -105, 105, -9, -112, 90, 12, -83, -89, 12, -29, -77, 37, -85, -88, -6, 54, -109, 37, 18, -52, 75, 107, 44, -14, -57, -86, -116, 87, 125, 13, 30, 46, 81, 27, 38, 118, -31, -72, -30, -92, -55, -40, 103, -2, -34, 126, -109, -97, -90, -101, 29, -60, -107, -120, -5, 70, 120, -78, -116, 118, -79, -65, -58, -55, -40, -100, -56, 10, 88, 104, -56, -113, -42, -31, -105, -127, 37, -125, 47, -21, 127, -99, 68, -44, 109, -24, -71, 4, -119, -68, -65, -36, 109, 61, -13, 41, -88, 76, 105, 54, 21, -117, 33, 8, -64, -81, 1, -67, 27, 39, -99, 52, -102, 122, 44, -122, 65, 29, 7, -73, 82, 34, -96, -79, 6, -39, 24, 116, -19, -112, -54, -61, 19, 27, 73, -39, -64, -63, 51, 83, 7, 1, 71, -19, -103, -45, -106, 27, -3, -63, -18, 71, -110, 56, -85, -47, -12, -31, -77, -34, 96, -115, 75, -40, -52, 23, 17, -114, 103, 38, -86, 58, 26, 35, -94, -47, -42, 108, 121, -22, -49, -89, -88, -27, -55, 4, -14, -67, -110, -78, 8, 3, -57, -126, 115, 24, 42, -97, 38, -19, -22, -99, 57, -111, -22, -114, -103, 28, -93, -11, 105, -40, 115, 37, 73, -30, -84, -38, -42, 39, -95, -106, 58, -103, 38, 90, 23, 33, 91, -95, -37, -49, -71, 3, 53, -56, 45, 6, -104, 120, -127, 53, 98, -101, 86, -112, 41, 80, 65, -121, 37, -93, 124, 113, 31, -7, -128, 62, -27, 49, 23, -102, 42, -15, 89, 29, 73, -1, 107, -5, 107, -51, -5, 124, 69, -48, -7, 15, 101, -19, -118, 42, 12, 42, -123, 92, 107, 11, 13, 76, 50, -102, -16, -119, 123, 105, 32, 18, 44, 42, -24, -21, 122, 2, -91, 103, -105, 16, -109, 74, 118, 91, 58, 65, -108, -88, 19, 83, -46, 11, -119, -43, -71, 98, -50, 69, -14, 29, -25, 72, 36, -103, -35, 9, 20, 22, -16, 20, -70, -53, -71, -80, -105, 34, 16, 43, -104, -49, -15, -54, -91, 81, -50, -30, 29, 47, -121, -2, -1, -66, -122, 50, 66, 32, 9, 68, 61, -38, -6, 87, 43, -27, 58, 112, -46, 34, 8, 81, 45, 36, 122, -31, -54, -112, 76, 58, 67, -8, -80, -105, -48, 10, -22, -69, 122, 109, -116, 58, -16, 127, 105, 59, 43, -15, -36, -90, -44, 122, 69, -9, 91, 42, 36, 110, -47, -41, -7, -6, 48, 91, -22, -64, -56, 13, 116, -80, -98, -20, 121, -46, 79, 14, -7, -24, -28, -3, 122, -118, -81, -40, -83, 38, 77, 1, -62, 106, 83, -51, -126, -83, 44, -20, 82, 23, 20, 20, 78, 96, -101, 15, -30, -125, 17, 27, -89, -117, 35, -117, -45, 111, 101, 120, 84, 18, 78, 2, -61, 97, 90, 60, 118, 56, 79, 76, -97, 60, -102, 116, -40, 121, 65, -8, -55, 45, -103, -7, 1, -47, 35, 108, -34, 27, 66, -107, -26, 38, -33, 25, -75, 22, -9, 46, 33, 23, 58, -112, 106, -11, 72, 8, 82, 11, 29, -2, -33, -107, -6, -84, -84, -78, 77, 78, 70, 114, -69, 116, -40, -106, -18, 38, -119, -82, 61, 118, -76, -109, 1, -37, -97, 52, 46, 31, 82, 118, 40, 124, 126, -29, 62, -119, 74, -56, 93, 15, -63, 15, -45, 123, -37, 73, -100, -46, 20, -91, 125, -5, 75, 103, 30, 121, -43, 58, 68, -101, 53, -106, 94, -116, 99, 100, 78, 23, -25, -73, 62, -92, -47, 30, -98, -108, 16, -93, 100, -91, -110, -74, -110, -4, -67, -79, -81, 52, -39, 108, -36, -29, 116, 38, 127, -21, -1, 81, 120, 122, 40, -121, 67, 51, -77, 80, 65, 41, 100, 122, -41, -124, -90, -61, 101, -127, -114, -114, -61, 85, -91, 4, 61, -84, -106, -60, 70, -28, 68, 117, 88, 14, 62, 117, -30, -78, 67, 79, 112, 99, -105, -106, -39, 127, 19, 84, 2, -128, 20, 26, 34, -91, -112, -38, 74, -98, 81, 72, 73, -48, 49, 83, -40, -96, -13, 5, 37, -88, -59, 58, 15, 78, -109, 111, -49, 9, 103, -55, 1, -86, 80, 91, 100, 95, -51, 24, -45, -85, 48, 124, -82, -2, 42, -37, -17, 13, 67, -111, 58, 44, 42, -20, 41, -69, -103, 49, 112, 109, -44, 25, -123, -76, 123, -7, 81, -68, -5, 95, -11, 65, 96, 102, -96, 37, 74, -86, 90, -39, 125, -76, 62, 53, 64, -93, 19, 41, -15, 15, -122, 44, 86, -100, -59, 32, -82, 16, 20, -57, -97, 1, -9, 23, 109, 30, 108, 109, 20, -10, -70, -29, -93, -94, 119, 3, -94, 65, 108, -94, 82, -86, -111, 90, 88, 13, -2, 34, 41, 60, 53, -50, -105, 97, 122, -40, -45, -49, -94, -123, 74, 3, 98, 71, -32, -71, 70, 47, -39, -60, -24, 90, 23, -111, -91, 89, 92, -12, 35, -59, -15, 86, 116, -25, 27, -79, 23, 10, -115, 88, 58, 96, -49, 23, -113, 53, 50, 24, -2, 9, -72, 36, -57, 123, 75, -122, 118, 98, 80, 121, 126, 20, 96, -15, 83, -96, -58, 114, 50, -50, 35, 54, -50, -82, 95, -54, -55, 5, 63, 54, 104, 127, -11, -70, 32, 1, -118, -16, 15, -25, 28, -81, 19, -84, 58, -37, -42, 105, 78, 109, -110, -41, -14, 124, -24, 61, 66, -72, 28, 41, -49, -25, 26, -76, 50, 33, 23, -7, -92, -69, -128, 51, -60, 44, -101, -87, 124, 69, 88, -78, 52, -71, -29, 64, -5, -94, -75, -86, 8, 31, -41, 68, -32, 82, 117, -30, 121, -83, -2, -59, 52, -111, 28, 55, -30, 19, 7, 20, -34, 115, -35, -102, 109, -35, -126, 47, -99, 79, -12, -3, 108, 27, 114, 52, -43, -112, 73, 63, -22, -118, 92, 30, -110, 92, 123, -126, 46, 39, 86, 114, -83, 64, 68, -67, -74, -115, -24, -51, -94, -114, -40, -40, -51, -39, -75, -24, -74, 51, 78, 114, -1, -58, -121, -70, 122, -123, 89, 104, -75, -76, 101, -102, 4, -63, 70, 111, -93, 72, 116, 66, -84, -83, 4, 91, 96, 24, -33, -113, -88, -57, -76, 7, -79, -83, 55, -35, 2, 89, -47, 95, 62, -14, -97, -95, -101, 103, 38, 109, 59, 99, 0, 14, 34, -114, 13, 54, -118, 12, 101, -67, -48, -22, 122, -43, 106, -125, -22, -93, 112, 3, 80, 28, -121, 23, 36, 65, -77, -100, -104, 103, -17, -71, -102, -10, -16, 23, 21, -120, 57, 37, 65, -121, -22, -59, -111, -77, -17, -124, -114, -37, 43, 25, 52, -70, 104, -107, 89, 83, 26, 23, -126, 42, 13, -105, -112, -12, -107, 112, 59, 57, -84, 123, -106, -27, 31, 13, -109, 55, 97, 88, 72, -36, -38, 112, 119, -107, 5, 104, 107, -66, -3, -73, 9, -120, 26, 90, 41, -24, 40, 63, -111, 22, 43, 1, -35, 45, -72, -54, 74, 44, 93, 14, 13, -126, -124, 110, -8, 13, -112, -83, 127, 57, 5, -68, -111, -78, -38, -94, 119, -69, -108, -10, 64, -7, -84, 81, 15, -103, 125, 58, 69, -88, 1, -90, -48, -7, 108, 63, -6, -59, 68, -12, 100, -3, -30, 100, -94, 112, -69, 22, -81, 2, -41, 62, -78, -45, 106, -107, 46, 104, 112, -105, -5, 17, 80, -35, 46, 25, -82, -115, -122, -2, -113, 80, 49, 66, -59, -93, 47, -119, -54, 114, -114, -85, -59, 54, 13, 11, 58, -90, 59, -8, 60, -117, 37, 89, -9, 96, 109, 4, -73, 112, 56, 53, -105, -73, 4, -13, 37, 122, 84, -79, 14, -11, -112, 91, 23, -78, 39, 95, 99, -69, -69, -3, 53, -24, -61, -78, -118, -31, -71, -14, 119, -11, 91, 103, 68, -86, 86, -113, -96, 67, 49, 31, 93, -41, 28, 112, 7, 120, 32, -18, 35, -27, 6, 93, -120, 51, 125, -98, 81, -31, 18, -6, 84, -88, 111, 72, 4, 18, 106, -111, -5, -89, -121, -38, -59, 72, -102, 85, 94, 107, -24, 102, -117, 104, 88, 52, 44, -108, 100, -114, -37, -26, -110, -23, -94, 104, 47, 126, 34, 78, 61, -115, -108, -5, 49, -79, -114, -30, 86, -124, -52, 10, 1, -121, 59, 17, -112, 27, -99, -42, -73, -77, -82, 17, 52, -10, -36, 45, 83, -47, -11, -33, 32, 7, 50, -55, 74, -66, -73, 98, -29, 126, -122, -38, 60, 115, 119, 36, 54, 66, -10, -99, -100, -110, -48, 33, 45, 69, -87, 9, -63, -3, 32, 28, 45, 91, -80, 113, 79, 123, -106, 24, 16, 95, 98, -66, -127, 55, 99, 6, -71, 67, 124, -30, 116, -99, 106, 112, -89, -109, 61, -38, 89, 67, 25, -31, 81, -36, -78, -57, -30, -46, -9, -27, 48, 63, 109, -22, -102, -126, -49, -7, 106, -103, -127, -42, -50, 10, -57, 68, 124, 0, -62, -76, 112, 91, 62, 36, 32, 21, -121, -59, 88, 114, -5, 56, -12, 40, 104, -102, -6, 38, 127, -103, 50, -125, -36, 36, -41, 43, -86, 105, 3, -14, 46, -35, -87, 9, 59, 31, -91, -66, -64, -65, 2, -95, 118, 41, 68, 40, -36, 34, 21, 30, -99, 40, -67, -4, 21, 34, 19, -105, 84, -54, 38, -61, 124, -21, 2, 30, -65, 99, 122, -106, 16, 119, -11, 35, 58, -101, 58, -92, -80, -18, -33, 65, 115, -49, 72, -116, -107, 105, 29, 26, 123, 11, -107, 82, 14, 52, -41, 64, -14, -31, -107, -117, 95, -36, 14, 96, -75, -52, -56, 78, 87, 24, -47, 105, 84, 0, 100, 79, 95, 42, -54, -30, 115, -17, -21, -79, -46, -16, 82, -25, -90, -100, 71, -89, 67, -2, 111, 52, 68, -63, -72, -112, 73, -5, 73, -101, -56, -2, 121, 30, -35, -12, -42, 96, 25, -64, -57, 110, 90, -2, -126, 5, -7, 17, 58, -3, 119, -85, -121, 91, -33, 11, -40, 15, 85, 115, -82, 1, 0, 71, 10, 62, -117, -15, -6, 83, 112, -76, 10, 99, 69, 48, -15, 77, 43, -69, 29, -54, -121, 121, -114, -77, 30, -105, 20, -117, -44, 3, -69, -4, 0, 32, 75, 18, -49, -36, 106, -75, -16, -9, 96, 36, 102, 59, 126, -36, -18, 108, 47, 4, -6, -35, -55, -75, -38, -32, -82, -86, -3, 57, 125, 49, -13, -19, -83, -67, 73, 34, 41, 47, -103, -4, 71, -106, 53, 73, -104, 81, 85, 72, -92, 4, 103, -17, 70, 117, 47, -94, 39, 38, -116, 57, -74, 10, 105, -84, -26, -60, -55, 52, -46, -111, 117, 14, -91, 120, -11, 35, -67, -17, -71, -38, 120, 103, 106, 87, -95, 37, 42, -75, 13, -45, 18, -51, -46, -106, 29, 123, 112, -19, 5, 108, -47, -9, -35, 86, 29, 60, 73, -128, -86, -11, -120, 113, -38, 83, 120, -91, -5, -26, 88, -4, 107, -126, -38, -18, -127, 85, -82, 15, 93, -80, -45, 118, -63, -57, -18, -80, -24, 59, -128, -22, -73, -38, -61, -81, -116, 64, -19, -66, -62, -1, -1, 37, -46, 60, 3, 31, 16, 84, 45, 5, -10, 6, -39, -56, 24, -33, -29, -96, -68, 7, 117, -20, -119, 22, -119, -12, 45, 109, -25, -12, 65, -18, 78, 113, 84, -59, 17, -12, 85, -39, 61, -75, 48, -109, 24, -90, 46, 115, -126, -68, -30, 63, -15, 41, -94, -14, -16, -92, -90, 112, 44, -79, -122, -72, -112, -26, 57, 81, -101, -12, -98, 4, 118, 117, 49, -29, -37, -28, -103, 97, -51, 113, -52, 68, -56, 74, 5, 16, -16, 28, -103, -120, 41, -74, -92, 50, 70, 92, -125, -68, -37, -8, -37, -97, 121, 82, -1, -59, 84, -49, -6, -30, 112, -50, 84, -84, 56, 105, -55, 62, -115, 76, -55, -86, -19, -60, 43, 81, 80, 82, 94, -34, -127, -39, 88, 81, -16, 19, -77, -78, -57, 39, 19, 98, -100, 116, 102, -114, 56, 109, 79, 100, -122, -26, 7, 25, 63, -73, -36, -108, 52, -74, 104, -31, -48, -88, -53, -50, -99, -63, -83, 62, -29, -28, -98, -21, 112, -115, -35, 91, -62, -68, 109, 25, -40, -30, 25, -41, 1, -2, -102, -2, -124, -100, 42, 1, -57, 84, -78, -12, -95, 13, -117, 9, 112, -70, -3, 75, 30, 8, 98, -26, 4, 5, 106, 125, 115, 116, 6, -118, -39, -94, 20, 111, -114, 115, -46, -61, -18, 23, -47, 77, -16, -11, -32, -94, 31, -117, -51, 114, 40, -120, 127, -78, 50, 20, -5, -86, -83, 73, 3, 81, 67, -26, -4, 102, 89, 55, 21, -91, 10, 99, 87, -98, -2, -18, -7, -32, 33, 125, -37, -62, 20, 108, -54, -57, -29, -93, -122, -81, -95, 50, 73, 45, 5, 36, -23, -83, 15, -15, 36, 110, -66, 88, -21, 11, 54, -75, -20, 68, 14, -83, 69, 116, 45, -103, 95, -53, -64, 11, 43, 120, 43, 77, 111, -34, 12, -15, -8, -26, 65, -12, -51, 2, 7, -80, -106, 61, 124, -73, 13, 108, -19, -43, -66, -46, 103, -112, -73, -11, -48, -27, -30, -19, 78, -71, 54, 61, 61, 5, 121, -20, 126, 118, -22, -23, 38, -42, -117, 12, -101, -29, -114, 39, -3, -82, 123, -53, 68, 4, -59, 45, 58, -55, -10, 1, -61, -79, -20, -73, 78, 51, -122, 90, 34, -10, -87, 26, 105, 111, 43, -57, -4, 36, -121, 67, 83, 79, 33, 106, 76, 66, 43, -7, -89, 88, 40, -40, 51, -48, 71, -35, -14, -103, -109, 111, -58, 59, -52, -38, -49, 60, 91, -114, 4, 1, 5, -62, -27, 24, -46, -30, -118, -3, -76, 117, 88, 72, 127, -86, 100, -19, -40, 21, -91, 15, 125, 49, 124, 119, 117, -7, 30, -69, -52, -68, 106, 44, -27, 112, -123, 98, -79, 55, -77, 127, 113, -21, 5, 4, 48, 91, 109, 96, 53, 86, 114, -65, -44, 125, -100, -16, 0, 77, -21, -88, -37, -49, 66, -15, -94, 100, -63, -109, 30, -15, -123, -37, 110, -73, -53, 95, -74, 101, -17, 54, 65, 5, -30, 5, 105, -112, -121, -80, 58, -3, -85, -55, -101, -81, 63, -119, -26, -63, -47, 79, 74, 11, 66, -68, -68, -112, 52, -103, 64, 84, 100, -65, 59, 13, -15, -122, 122, 27, 89, 66, 119, 33, 28, -93, 124, 100, 43, -50, 68, 45, 90, 109, 47, 74, -19, 34, -41, 97, -37, 44, -9, 102, 59, -71, 15, -95, 68, 66, 42, 88, 89, -49, 36, 64, 81, 43, -64, 51, 107, 60, 49, -116, 87, -13, 7, -64, -29, 125, 123, 100, -111, 30, 118, -109, 113, 17, -118, 1, 28, -47, -36, 119, 56, -109, -73, 67, -72, 35, -111, 123, -5, 101, 18, -68, 120, 91, 65, 78, -88, 81, -109, -127, 48, 98, 88, 3, -25, 109, 102, 33, 85, -21, 2, -6, 124, 100, 29, -41, 102, -80, -68, -119, -47, 80, -99, 125, 113, 107, 34, 125, -101, -17, -48, 10, -33, -112, 108, 79, 48, 124, -68, -78, -83, -53, 20, 118, -105, 50, -37, -65, -75, -80, -104, -74, -104, -68, 57, -88, 47, 55, 99, -96, 55, -105, -54, -3, 6, 119, -36, 89, 96, 62, 19, 11, -90, 16, -29, 98, 113, 59, 115, -92, 104, -97, -60, 92, -98, 24, 119, 70, -22, 74, 11, -115, -127, 105, 112, 51, 112, 113, -79, 69, 112, 18, 37, -121, -31, 17, 56, -20, -69, -25, 20, -114, -93, -93, -16, 69, 104, -29, 24, -67, 115, -13, 115, 54, 15, -13, -123, -108, -6, -26, 33, 29, -23, 107, -99, 43, 117, -11, 24, -94, -8, 9, 41, -37, 40, -117, -54, 112, 52, -4, -56, -55, 1, 101, -14, 54, -78, -40, 90, -83, -92, -13, -107, 1, -51, 28, -64, -12, 117, 113, 40, 86, 60, 79, 41, 46, -18, -19, -56, -58, 63, -65, -76, 36, 110, -4, 96, 41, 73, 98, -58, 78, 56, -44, -88, -113, 91, 61, -81, -26, 64, 114, 2, 11, -30, 96, 36, -71, -16, 83, -109, 63, 76, 101, -19, 65, -54, -103, -40, 103, -24, 51, 82, 4, 56, 41, 66, 32, -43, -38, 12, 105, 47, 49, -42, 39, 13, -65, 9, -59, 29, 79, -105, 25, -33, 81, -62, -85, 22, 23, 57, 18, 115, 86, -94, 44, 6, -40, 118, -51, -28, -109, 15, -22, -25, -63, -60, 77, 123, -50, 119, -119, 81, -105, -40, -37, 84, -75, -77, -75, -50, 60, 102, 86, -62, -112, -32, -8, 0, 38, 115, 62, -112, 40, 33, 85, -43, 120, -7, 26, 122, -74, -89, -95, 78, -96, -54, 90, -106, 64, 11, 13, 41, 12, -88, -48, -67, 69, 107, -79, -39, -28, -46, -35, -22, -104, 57, -78, 77, -41, 108, 88, -106, 125, 58, -117, 15, 109, -74, -53, 126, -91, 85, 95, 94, -40, 98, -18, 59, 80, -121, 49, -36, 16, -64, -12, -35, -87, 98, -63, 79, -81, 71, 5, -92, -22, 19, -52, -19, 2, 89, -12, -102, 99, 83, 22, -33, 87, -99, -49, 126, 72, -88, -118, 37, 123, -106, -103, 8, -115, -92, 72, 119, -54, 21, 96, -72, -85, -90, -117, -50, 76, 39, 4, -26, 58, 16, -82, -54, 53, 36, -36, -25, -48, 126, 4, 47, 89, -115, 107, 79, 20, 26, 104, 59, -82, 27, 37, -105, 86, 51, 6, 42, 125, 27, -111, 104, 45, 121, -96, 44, -59, -23, -125, -21, 37, -24, 73, 57, -52, -2, 14, 37, -13, -111, -119, 5, -100, 27, 43, -86, 53, -84, -85, -63, -47, 74, -127, -128, 94, -34, -19, 93, 103, -66, 78, 81, 106, -10, -95, -47, 66, 77, 113, -73, 58, -71, -114, 3, -3, 42, -82, -29, 58, 51, -39, -103, 14, -81, -56, 25, 3, -83, 70, 88, 39, -98, 118, 124, -14, -15, -65, -92, 15, 33, 88, -16, -24, -118, 13, -104, -65, -86, 82, 115, 40, -42, -102, -114, -128, 39, -90, -94, -108, 105, 53, 3, 115, 68, 48, -69, -97, -91, -117, -64, 69, -22, 7, 66, 123, 17, -88, -99, -96, -100, 59, 6, 121, 75, 6, 2, 89, 10, 60, 4, -107, -73, -22, 96, -64, -118, 41, -42, -114, 8, -81, -76, 89, 51, -38, -104, 33, 85, 54, -103, 120, 86, 57, -22, -123, -52, -80, -90, 41, -127, 55, -95, 71, -77, -75, 54, -97, 43, 43, -51, -89, -70, -118, 104, -55, -25, 70, -96, -61, 96, -105, -75, 5, 39, 34, -100, -116, 61, 75, -99, 127, -46, 81, 20, -73, -34, -18, 126, 41, -74, 47, -76, -94, -125, 10, 18, 47, 32, -8, 103, 47, -70, 53, -109, 25, 20, 127, -78, 10, -88, -84, 18, 32, 103, 75, -83, -39, 68, 1, -52, 76, 80, 3, 35, -8, 77, 70, 15, -4, 4, 4, -22, 110, -64, 107, 99, -30, -114, -111, -125, -69, -86, -55, -15, -58, 17, 112, 115, 109, 38, 32, 72, 81, -50, -16, -89, 1, 88, 26, -87, -37, 4, -32, -22, 0, 63, 20, -43, -21, -106, -65, -33, 77, -113, -118, 100, 73, -24, -76, -42, -24, -20, 54, 0, -48, 110, 63, 118, 22, 76, 96, -3, -104, 108, -45, 41, -28, -120, 90, -10, -110, -31, -40, -36, 97, 57, 70, -69, -114, -35, 121, -6, -108, 92, -128, 91, 96, -102, 126, 47, -24, -86, 81, -125, 16, 86, 93, 79, 13, -124, -12, -17, 121, 123, 115, -27, 97, -60, -118, -30, 57, 21, -39, -119, 65, -111, -93, 6, -33, -52, -109, 23, 15, -121, 100, -55, 6, 76, -82, 68, 117, 108, -117, 119, 127, -32, 39, 119, -12, -89, -118, -19, 112, -121, 91, -26, 103, -128, -104, 57, -20, 74, 93, -62, -126, 70, 55, 52, 91, 70, 85, -49, -115, -96, 58, -17, 73, 106, -85, -9, -33, -10, -61, 127, -62, 19, -127, -92, -69, -34, 103, 55, 97, 123, -92, 69, 7, -46, -92, -53, 97, -94, -55, 59, -100, 9, 99, 22, 62, 42, 54, 2, -22, 12, -90, 20, 81, 102, -88, 93, -46, 45, -101, -23, 31, 25, 116, 60, -18, -84, -110, -36, 86, -125, 59, -23, -91, 109, -29, 84, 118, -72, 127, -109, 42, -106, -61, -119, 64, 2, -70, 63, 119, 120, 31, -7, 55, -14, -106, -31, 121, 45, -93, 91, -74, -3, 104, 4, -28, -96, 89, 82, 104, -124, -86, -61, -40, 40, -94, 56, 66, -81, -105, 60, 78, 65, -42, 79, 23, -86, -10, 80, -12, 124, 67, 61, 45, 100, -111, -57, 80, -38, -122, -75, 103, 58, 66, 31, 118, -27, 84, 3, -7, -7, -63, 126, -78, -4, -29, -30, 60, -116, 99, 38, -40, -21, -41, 26, 12, 9, 20, -113, -11, 33, -55, 98, 14, 98, -69, -52, 119, -43, -53, 104, 101, -68, -67, -83, 107, -19, -44, -20, -77, -127, -89, -115, -1, -110, -123, -105, -97, 39, -8, 58, -37, 72, 77, -1, 1, 63, 84, -104, 37, 100, 46, 125, 17, -128, -60, 55, -63, -69, -102, 96, -91, -65, 103, -127, -74, -5, -100, 41, -59, -100, 125, 100, -73, -99, 37, 56, -26, -33, 127, -25, 81, -32, 91, -37, 14, 45, -81, 5, -114, -27, -89, -87, -43, 64, 111, 12, -18, -116, -107, -13, -55, 95, 34, -23, -34, 44, -9, -8, 100, 2, -27, -106, -48, 85, 66, 36, -71, 113, -55, 120, 95, 85, -10, -17, -19, -74, 14, 65, -22, -77, -36, -81, -28, -71, 58, 122, 79, -35, 114, 35, 4, 34, -85, 99, 10, 114, -91, 44, -82, 71, 34, -28, -69, 4, -85, 116, 11, 71, -114, 106, 21, 10, -51, 73, -9, -105, -19, -106, -96, -87, -77, 82, -68, 80, 125, -49, -76, 28, 67, -76, -71, 120, 96, 50, 54, -44, 54, -67, 115, -19, -93, -66, -24, 66, -92, 13, 37, -23, 110, 109, 84, 53, -54, -7, 101, -15, -113, 123, 103, 62, 66, 97, 17, -101, 29, -113, 109, 71, -16, 13, -49, 86, 65, -29, 76, 28, -112, 6, -53, 124, 0, -34, -118, 9, -123, -5, -120, -112, 37, 37, -78, -98, -127, -48, 37, -102, -52, -119, -100, 42, 80, 62, -120, -115, -117, -47, -97, -94, -15, -65, -104, 80, 2, -122, -88, 64, -15, 89, 16, 74, 80, 1, -36, 98, 58, -91, 63, -91, 59, -77, -8, -83, -107, -73, 28, 0, 66, 47, 92, 65, 4, 50, 93, 97, -82, -113, -74, -127, -111, 122, -111, 53, -108, 118, -84, 69, -3, -8, -64, 39, -123, -51, -127, -127, -67, 56, -103, 44, -5, 96, -19, 45, 76, -50, -98, 62, -80, 48, -83, -87, 56, 19, -89, -95, 21, 13, 89, 11, 127, 61, 71, 81, 102, -112, 73, -83, 113, -30, 32, -38, -53, -108, -49, 62, -58, -107, 113, 97, -21, -125, 126, 25, -54, 12, -115, 105, 37, 22, -79, 108, 45, -106, 21, 1, 94, -19, -103, 2, -45, -62, 102, 76, 73, -13, -74, 82, 118, -46, 29, 35, -111, 39, -58, 77, 93, 41, 72, -13, -9, 117, 107, 121, -14, -40, 23, -126, 45, 67, -39, -23, 66, -108, 97, -121, -25, 0, 45, 56, 67, -109, -124, 63, -77, 73, -44, 67, -59, -68, 101, -48, 102, -14, 123, 65, -75, -120, -104, 18, 114, 31, -10, 80, 6, 115, 75, -31, 40, -38, -87, -15, 59, -77, -13, -126, -94, 49, -113, 56, 74, 127, 34, 78, -90, 27, 74, 12, 81, -34, 123, -21, 24, -121, -11, 26, 51, -38, 59, 110, 52, 91, 7, 55, -34, 126, 126, 96, -115, 68, 24, 68, 127, 57, -84, 103, -44, -97, -30, 34, -10, 105, 107, -66, 75, 123, -99, 38, -78, -102, 105, -96, -12, 46, -35, 35, 45, -126, -83, 0, -82, 101, -68, -41, -79, -52, 102, -61, -59, -74, 29, 14, -61, 86, 61, 118, -57, 118, 2, 111, 0, 117, -97, 83, -43, 117, 70, 88, 14, 33, 70, -8, -16, 91, -25, -27, 65, 111, 45, 124, -64, 113, -112, -44, -67, 117, -55, -98, 25, -83, 24, 26, 17, -48, -40, 97, 82, 36, 127, -5, 91, 41, -128, 20, 88, -74, -90, -108, -32, 88, 113, 106, 98, 3, 78, -118, 108, -13, 31, -24, 77, 78, 30, -25, -120, 0, 113, 27, -77, -15, 5, 97, 53, -17, -50, -67, 61, 79, -39, -1, -66, -2, 42, 79, -57, 18, -76, -1, -56, 113, -82, -115, 33, -51, 109, -88, 36, 22, 85, -35, 96, 25, 82, 13, -17, 80, -42, 103, -47, 46, 85, 18, -32, -33, 17, 14, 61, 25, 69, 36, -95, -46, -92, -122, 33, -43, 110, 40, -22, 126, -19, -76, 33, 42, -113, 8, 68, -53, -1, -74, 36, -92, -72, 4, -26, 124, 50, 56, -85, 103, 95, 115, 12, -92, 91, -101, 17, -111, 122, -71, -18, -88, 5, -107, 12, -57, 69, 49, 97, 53, 44, 0, 87, -85, -70, -58, -123, -25, 59, 90, 8, -1, -45, -17, -78, -119, -5, 57, -34, -69, 116, 36, -103, -20, 111, -49, -123, -102, -65, -16, 83, 4, -114, -112, 98, -65, -95, 100, 1, -69, 83, -37, -74, -117, 72, -93, -41, -95, 74, 33, 60, -81, -69, 3, 69, -115, 8, 114, 6, 30, 122, 91, 32, 64, 9, 125, -55, -18, 8, -29, -69, -100, 112, -51, 110, -65, -22, -127, 75, -61, 120, -84, -102, 45, 3, -28, -48, 57, 80, -29, -114, 80, 17, 114, 14, -10, 32, 82, 63, -95, 5, -60, -86, -14, 85, -39, -91, -17, 10, -69, 73, -62, 15, -127, -71, 20, 17, 89, -63, 2, -99, 113, -96, -113, -24, -24, -117, 127, 86, 31, 2, -6, -32, -76, 41, -94, 57, -30, -18, 21, 44, -1, 87, -18, -117, 69, -106, 118, 115, 100, -71, -42, -118, 10, -63, -19, -3, 4, 113, -83, -42, 45, -68, -70, -70, -7, -27, 120, -103, -39, -55, 27, -18, -122, -118, 31, 100, -91, 82, -93, -36, 68, 15, -47, -99, -104, 74, 55, -55, -68, -60, 115, 46, -21, 24, 5, 45, 33, 8, 96, -40, 29, -64, 66, 29, -83, 109, 23, -112, 80, 64, -29, 12, -66, 25, 125, 75, 44, 108, 108, -42, -69, -8, 58, 34, 35, 83, 63, -17, 51, -37, -13, 41, 22, -71, -119, 48, 13, -104, 114, 84, -10, -7, 90, -94, -36, -36, -53, -3, -42, -71, -110, -83, -128, -118, -98, 91, -16, -13, 68, -95, 16, -63, 13, 21, -67, 85, -33, -22, -90, -84, 79, -27, -18, -28, -15, 44, -112, 29, 13, -30, -13, -59, 52, -80, 92, -106, 116, -119, 86, -14, 109, -113, 119, 38, 49, -92, 9, -113, 72, 39, 19, 36, -25, -18, -48, 75, -76, -83, -15, -30, -70, -126, 104, 124, -11, 107, 84, 108, 63, 36, 7, -50, 95, -102, 3, 20, -8, 101, -90, 47, 40, 57, -38, -109, -112, 52, -17, 60, -55, -7, 70, -27, -57, 101, -59, -104, 34, 32, 59, -49, 63, 16, -110, 118, 35, 108, 90, 115, 86, -79, -51, 65, 77, 101, -84, -13, -94, 37, -26, -79, -62, -46, -60, 29, -122, -107, 122, -118, -47, -43, 120, -37, -27, 8, -79, 34, 57, -59, -112, 123, 113, -125, -57, -24, 124, -39, -121, -75, 125, 112, 3, 50, -7, -52, 2, -100, -77, 72, -50, -86, 95, 61, -50, -55, 89, 106, 71, 53, -106, 89, 67, -56, -64, -101, 41, -58, 39, -13, -105, -108, 62, -13, 65, 7, 64, -18, -84, -69, -84, 24, -67, 51, 122, -11, -121, 63, 7, 50, -24, 19, -41, 106, 34, -122, 84, 29, 104, -50, -52, 37, 63, 40, 3, -56, -70, 44, -5, -119, -41, -38, 107, 27, -109, -41, -20, 84, -106, -122, -114, 17, 25, -48, -88, 75, -127, -60, -20, 102, -60, 84, 116, 114, -25, -71, -18, -98, 122, 84, -69, 125, -107, 40, -10, -88, 32, -88, -80, -80, -20, 13, -36, 85, -97, 97, -75, -31, -28, 42, -83, 21, -120, -59, 98, -5, 36, -23, -89, -21, 38, -14, 44, 58, -32, 119, -46, -56, 87, 79, -6, -18, -70, -64, -106, 112, 13, 64, 95, 51, 114, 7, -54 );
    signal scenario_output : scenario_type :=( -128, 127, -8, -128, -24, -128, 42, -5, 127, -128, 107, 16, -128, 127, -128, 24, 127, -128, 127, 12, -128, -124, -128, -128, 127, 13, 127, 127, -128, 121, -128, -128, 127, 32, 127, 39, -128, -128, -128, -128, 1, -3, 127, 127, 0, -128, -128, -128, -128, 127, -28, -128, 127, -128, -128, 117, -128, -128, -128, -16, -128, 127, 127, -121, -29, -128, -57, 127, 95, 1, 127, -128, 127, 74, 122, 18, -128, -128, -128, -42, -128, 127, 42, -128, 127, -128, 127, -53, 76, 127, -97, 127, -128, -128, 127, -128, 66, 116, 127, 60, 127, 10, -128, -128, -128, -42, 54, 127, -64, 0, -6, -76, -74, -81, -44, -128, -2, -18, -24, 127, 127, 127, 127, 127, -128, -128, 127, -90, 90, 127, -128, -32, 127, 112, 47, -128, -128, -59, 109, 127, 116, 127, 90, 127, -117, -128, 80, 127, 127, 127, 127, 127, 127, -128, -85, -92, -85, 127, -60, -16, -128, -43, -128, -128, -92, -24, -100, 74, -128, -128, 70, -15, 127, 127, -1, 127, -52, 127, 31, -128, 127, -128, 127, 32, -128, 74, -128, 88, 127, 127, 127, 64, -73, 127, 127, -16, -100, 116, -128, -128, 127, 16, -128, 127, -6, -128, -15, -128, -128, -50, 24, 127, 127, 127, -55, 10, -128, -128, -128, -55, 127, 127, 65, 127, -87, 0, 26, 33, 96, 127, 102, 111, 21, 47, 127, 127, 127, 127, -64, -128, -107, 127, 118, 47, -128, -128, -128, -128, 127, 7, -124, 48, 100, -128, 119, 127, -58, 26, -95, -128, -128, -11, -128, 26, 73, 127, 127, 109, 127, 107, -128, -37, -33, -128, 111, 76, -128, 127, 23, -98, 127, -17, -78, -128, -128, -31, -128, -128, -17, 11, 42, 127, 127, 127, -74, 127, -128, -128, 18, 0, -128, -28, -128, -53, -12, 127, 78, 127, 127, 127, 127, -128, -128, -128, -128, -128, -128, -27, -128, -13, 97, 7, 127, 127, 10, 22, -36, 78, -71, -11, 112, 127, 127, 16, 127, -128, -27, 127, -128, -69, -32, 11, 68, 81, 127, 17, 127, 127, -128, 127, -128, 3, 127, -17, -128, 33, 127, 114, 55, -63, -128, -128, -124, -128, 127, 96, 93, 127, 11, 127, -119, -100, -128, -128, 39, 101, -81, 127, -71, 127, 127, -128, -128, -102, -128, 3, -73, 127, -29, -108, -38, -107, -6, -128, -128, 75, -128, -79, 127, -128, 55, 127, -128, 127, 87, -108, 127, 101, -42, 127, -128, 65, 127, -128, 127, -128, -127, -43, -128, 127, 78, -128, 50, -32, -128, -24, -85, -6, 59, 127, 127, 127, -108, 32, -128, 37, 127, 127, 109, 87, -11, -128, -128, -37, -128, -128, -18, 76, 127, 127, 127, -121, -128, -128, -128, -13, -108, -128, -100, -128, -128, 114, -128, 127, 53, -128, -128, -128, -128, -128, -128, -128, -12, -128, 127, -34, -18, 108, -128, -7, -128, -128, 91, -106, -128, -128, 54, -50, 53, -73, -87, -128, -128, -70, 39, 127, 127, 127, 127, 31, -128, 48, -128, -128, 60, 127, 127, 127, 127, -16, 127, -128, 127, -74, -119, 127, 127, 118, 114, 127, -32, -128, 50, -128, -55, 127, 63, 113, -128, -128, 123, -128, 50, 75, 123, 127, 127, -66, -106, -128, -128, -123, -128, 59, -128, -128, 31, 60, 127, 127, 127, -34, 127, -128, -128, -76, 107, 118, 108, 127, 22, 96, 127, -3, 43, 127, 31, -23, 127, -128, -128, 127, -54, -39, 127, -54, 49, 127, -6, 98, -128, -128, -128, 3, 127, 127, 127, 127, -102, 85, -128, -128, -128, -8, -118, -128, 96, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -128, 3, -95, -71, 127, 127, 127, -49, 127, -39, -33, 101, -128, 50, -128, -128, 66, -29, 127, 127, 127, 127, -48, 127, -128, -128, 52, 7, 127, 52, 127, -18, -128, -128, -128, -128, -128, -128, -95, -128, -128, -10, 127, 87, 127, -128, -128, 127, -118, 127, 127, -124, -65, -128, 71, 86, -52, -124, 127, -101, -128, 106, 119, -65, -39, 127, -128, -128, 127, -87, -128, -22, -114, 127, 127, -26, 36, -2, 127, 127, 127, -74, 79, -128, -13, 127, 127, -128, 95, -128, -93, 127, -17, -128, 127, -128, -128, 48, -128, 8, 127, -128, 45, -128, -69, 127, 37, 127, 127, 127, 49, 127, 5, 13, 58, -117, 127, 70, 108, -15, -128, -58, -128, -128, -128, -95, -128, -128, 127, -128, 127, 127, -128, -128, 66, -97, 127, 85, 108, -34, 92, 70, -7, 127, 48, -128, -128, -27, -128, 127, 127, -21, 127, -26, -113, 55, 0, 111, 127, 127, 122, 127, 49, -128, -128, -128, -128, 38, -54, 48, 127, -128, -32, 101, -7, -108, 29, -128, -128, -32, -128, -128, -128, 86, -101, 73, -124, -128, 121, -1, -52, -128, -109, 127, 39, 39, -128, -128, -128, -128, -48, 127, 127, -128, -34, -60, -128, 18, -128, 29, 2, -128, 116, -128, -128, -114, 16, -6, -15, 53, -128, -128, 127, -123, 127, 64, -128, -10, -128, -128, 127, 127, -88, 127, 117, 100, -16, 75, 127, 23, 127, 127, -13, 127, -26, 32, 127, 49, -128, -128, -128, 60, 71, 127, 98, -128, -128, -128, -95, 127, 24, -118, -128, -128, -128, -128, 127, -114, -128, -106, -128, -128, 31, -128, 24, 102, -128, 127, 123, -128, 127, -93, -128, 127, -128, 63, 87, 127, -42, 88, -121, -43, -128, -6, -128, -37, -31, 108, 127, 127, 127, 127, 127, 127, 127, 117, -22, -128, 57, -128, 74, 44, -128, -33, 8, -47, 101, -128, -45, -128, -43, 127, 107, 88, -109, -128, -128, -128, 123, -128, 118, 63, 39, 127, -128, 92, 127, 122, 127, 52, 127, -75, -128, -128, -116, -128, 127, -31, 127, 127, -128, 127, -60, -128, -85, 21, -128, 44, 127, -128, 127, 127, 127, 127, 127, -28, 127, -128, -60, -92, -128, 15, -128, 127, -88, -128, 66, -12, -5, 127, 127, 5, 127, 127, -128, 127, 98, -128, 127, -128, 127, 24, 127, 127, -128, -85, -128, 48, 127, 127, 127, 127, 53, 127, 127, -64, 38, -128, -128, 117, -128, -33, 18, -42, -128, -5, 37, -128, -128, 15, -128, -8, 113, 80, 44, 127, -128, 75, -91, -80, 127, 127, 127, 127, 127, 33, 96, -128, -128, -127, -128, -128, 127, 127, 53, 81, -128, -128, -128, -68, -128, -66, -128, -128, 127, -12, 127, 127, 127, -71, 127, -128, 38, 127, 108, 127, -128, -128, -128, -123, -50, 127, 39, 127, -69, 73, -128, -122, -31, 75, 127, 101, 42, 127, -80, -13, -18, -128, -128, -128, 68, -36, 127, -31, 127, 33, -33, 59, 80, 127, -74, 43, -128, 127, -128, 24, 127, 73, 127, 10, -128, 38, 28, -22, 127, -128, -116, 7, -69, 127, -31, -128, -128, -100, 85, -128, 127, -65, -128, 68, 64, -113, 74, 71, 127, 75, 127, -24, -50, -98, 23, 21, -74, 60, -128, 127, -68, 55, -48, 111, -128, 112, 29, -128, -128, -128, -50, -128, 127, 0, -73, -38, 58, 17, 127, 1, -22, -128, -52, 36, -75, 127, -128, -128, 127, 55, 127, -128, -108, 10, 127, 127, -128, -96, -128, -121, 127, 78, -68, -128, -128, -127, 118, 127, 127, 127, -128, -128, -128, -128, -128, 127, -128, 127, 127, -66, 127, -127, -54, 7, 127, 28, -128, -32, 0, -66, 127, 127, -114, -31, -121, 112, 127, 127, -118, -119, -128, -128, 116, -86, -128, -11, -128, -128, -123, -88, -128, -26, -73, -49, -34, 127, 49, 127, 127, 127, 127, -128, -128, -28, 127, 127, 127, 87, 54, -52, -128, 28, -128, 85, 127, 127, 127, 112, -113, 95, -128, 119, 34, -128, 68, -5, 88, 127, 127, -64, 6, -128, -117, 127, 24, 127, 127, 127, 127, 127, 127, 127, -128, 71, 127, 81, 127, 106, -81, 60, -128, 15, -128, -109, 31, 127, 76, 127, 127, 101, 117, 127, -92, 43, -128, -128, -128, -16, -124, -128, -114, -128, -32, 127, 127, 127, 64, -75, 65, -128, -7, 96, -128, -31, 127, 102, -7, -96, -52, 27, -116, 127, -32, -128, -34, -128, -128, -28, 127, 127, -58, 100, 127, 44, 119, -128, -128, -128, -49, -128, -98, 42, -128, 127, -128, -128, 39, 18, -1, 127, 63, -13, 127, 127, -13, 127, -87, -128, 127, -31, 127, 127, -128, 127, -128, -12, 127, 127, 127, 127, -128, -128, 127, -128, 127, 96, 0, 127, 127, 127, 127, 127, -128, 127, 127, -102, -124, -128, -128, 90, 2, -91, -109, -128, -128, 22, -128, 127, -116, -128, -26, 48, -42, -69, 24, -54, 60, 127, 127, 8, -128, -128, 111, 127, 50, 127, -128, 5, 113, 127, 127, 127, -7, -128, -128, -128, 109, -128, -88, 127, -128, 55, 127, 45, -70, -118, -18, 114, 29, 127, 127, 127, 127, -26, -128, -128, -128, -48, 122, 127, -10, 114, -128, -2, -128, -128, -53, -128, 127, -57, 127, -128, 47, 127, 3, 127, -38, -128, -128, -128, -128, -122, 60, 127, 127, 127, 73, 127, 127, 127, 127, 127, 18, 71, -128, -128, -128, -128, 108, -128, 54, 127, 127, 127, -74, -34, -128, 127, -95, 114, -28, -75, 127, 127, 127, 118, -36, 127, 71, -81, -113, -128, 66, -128, 48, 127, -128, 127, 127, -102, -26, 81, 18, 15, -92, -128, -128, -3, 127, 127, 37, -128, -128, -128, -128, -128, -128, -112, 100, -32, -128, -128, 39, -128, 127, 85, -128, 93, -128, 127, 127, 73, 63, -15, -128, -128, 59, 123, 81, -116, -128, -128, -39, 127, -97, -128, -3, -128, 127, -128, -48, 127, 52, -63, -97, 1, -128, 127, 111, -87, 127, -79, 70, 127, 58, 36, 127, -128, -128, 2, 127, 127, -128, 127, 57, -128, 93, 91, 127, 127, 34, -2, -128, 57, 18, 127, 127, 127, 127, 6, -24, -128, -128, -128, -128, 68, -128, 127, 127, -128, 127, 123, -128, 127, -128, -128, 127, -58, 127, -113, 112, -128, 38, 78, -79, 127, -128, -58, 53, -18, 11, 127, -55, 31, 117, 116, 127, -128, 108, 47, -128, 5, 127, 18, 6, 127, -128, 127, 127, 127, 127, 118, -128, -128, -58, -73, 127, -128, 17, -22, 127, -7, -15, -95, -128, 127, -33, 27, 127, 78, 127, -6, 127, -128, -97, -128, -128, -128, 127, 127, -128, 127, -128, 103, -128, 43, -10, -65, 127, 127, 127, 127, -128, -128, -128, -98, 103, 127, -85, 127, -29, -128, 127, 127, 127, 90, -128, -128, -128, 1, 127, 127, 64, 127, -111, 127, 127, -118, -53, -128, -128, -128, -27, 127, -128, -18, -128, 127, -53, 27, 85, -128, 127, 29, 127, 127, -128, -128, -128, -128, -93, 127, 127, 90, 127, -68, 127, 121, -68, 37, -128, -128, -128, -128, -128, 97, -128, 127, 91, -128, 50, -26, 127, 127, 127, 7, -119, -128, 64, 121, -128, -95, -128, -1, 127, 127, 127, -128, -2, 49, 44, -128, 127, -128, -128, -128, -107, -58, -128, -28, -75, 44, 48, -128, 54, -128, -88, 96, 127, 127, 1, 96, -121, 28, 127, -128, 49, 70, 127, 127, 37, 117, 74, 127, 127, 107, -128, -97, -128, -128, -128, -43, -2, -49, 24, 127, -80, 127, 102, 91, -128, -21, 47, 34, 127, 127, 121, 87, 127, 75, 127, 127, -65, 127, -128, -66, 74, 63, 127, 127, 122, -122, -102, -85, 127, 127, 127, -33, 127, -128, 112, 127, -128, 111, 92, -128, 58, 127, -47, 108, -128, -65, 123, -50, -73, -3, -59, -80, -98, -128, -128, 91, 127, 127, -128, -128, -93, 127, 127, 127, 69, 127, 127, -128, -128, -60, -128, 127, 127, 8, 127, 76, 70, 127, 59, 37, 127, -128, 108, 127, -128, 69, -128, 6, 127, 108, 127, 97, -114, 75, -3, -50, 127, -128, 127, -70, 127, -85, -128, 127, -74, 127, -128, -128, -106, 8, 127, 68, 127, 127, 68, 127, 127, 69, 127, 127, 127, 34, 127, -128, 111, 127, -112, -11, 73, -65, 121, -119, 16, -75, -128, 10, -128, -128, 21, -70, -128, -128, -128, -128, -44, 127, -45, 127, 113, -58, 127, 53, -116, -6, 102, -29, 127, 127, -42, 78, -128, -128, -128, -34, -102, 127, 91, -128, -128, 32, 73, -59, 127, 36, -128, 75, -128, -76, 127, 37, 17, 31, 127, 127, 127, -8, 76, 71, 127, 71, 119, -79, -128, -121, -128, -49, -128, -31, 71, -37, -92, 0, -128, -128, -92, -128, -128, -128, -107, -128, 127, 127, 69, -128, 0, -128, 80, 127, 18, 52, -128, 64, -63, 13, 127, 127, 121, 127, 127, 127, 127, -12, 127, -128, 127, -128, -29, 127, 127, 122, 127, 127, -128, 80, 47, 127, 36, 127, 48, -64, 76, 127, 127, -28, 124, 127, -118, 57, 123, 127, 127, 96, -21, -128, -73, -128, -128, -34, -8, -38, -43, -128, -128, 8, 68, 45, 127, 127, 49, 127, -6, 75, 127, 127, 98, 127, 33, -128, 108, -128, -128, -22, -128, 42, -128, 122, 127, -124, -18, -128, -128, -128, -3, -12, 127, -128, 57, 60, 13, 127, 127, 127, 127, -13, 127, 92, -128, 127, -128, -128, 127, 127, 127, 119, -53, 127, 127, 127, 127, 8, 127, 32, -118, 21, 23, 127, 0, 116, 34, 127, 127, -50, -78, -128, -18, -75, 50, 127, -5, 127, 127, 127, 123, -128, -33, 81, 127, 127, 127, 127, 127, 24, 29, 127, 70, 127, -128, -128, -128, -53, 127, 28, -128, 127, -48, 127, -44, 8, -128, -60, -128, -128, 50, 127, 108, -128, -65, -128, 127, 127, -128, 127, -12, -128, -121, -15, -128, -1, -128, -98, 127, 112, 127, 93, -34, -128, 101, -87, -128, 127, -21, -78, -128, -106, 31, -128, 127, -66, 0, 87, -128, -128, 64, 127, 127, 54, -109, -6, 127, 47, 127, 91, -128, 127, 66, -128, 127, -128, -128, 127, 65, -128, -31, -90, -123, 127, 127, 127, 127, 85, -128, 127, -128, -49, 127, -128, 127, 127, -71, 127, 127, -12, -70, -128, 87, 36, 127, 1, 87, 80, -128, 95, -128, 12, -128, -121, -128, -128, -47, 5, 127, 127, 127, -128, 21, 10, -31, 127, -128, -128, -23, -128, -128, -128, -128, -128, -128, 17, -128, 59, 13, -98, -12, 16, -50, 127, 127, 79, 127, -128, -45, -128, 114, 55, -128, -128, 90, -128, 127, 127, -128, -74, 127, -79, -7, -128, 2, -128, -38, -2, -128, -42, -128, -128, -128, -128, 39, -87, 127, 118, -88, 127, -86, -128, 78, 127, 127, 127, 127, -128, -128, -128, 49, -128, -29, 70, -128, 74, -128, -79, -128, 2, -128, -128, -128, -128, 127, -6, 112, -128, -127, -31, 127, 127, 127, 90, -128, -128, -65, -128, 127, 127, 16, -128, -36, -128, -128, 23, -128, 74, 52, 66, 127, -29, 127, 127, -118, 33, 98, 103, 79, 127, 127, 90, 17, -128, -128, -29, 127, 127, -128, 70, 12, -128, 127, 26, 127, 127, 37, 33, 127, -1, -128, -107, 88, -128, 78, 5, 127, -2, 0, 127, 2, 127, 54, 48, -128, 127, 127, -128, 1, -73, 123, 127, 127, 127, 80, -102, -128, -128, -79, 113, 127, -15, -128, -64, -128, 127, -6, 78, -79, -128, 123, -103, 101, 127, 127, 127, 127, 31, 127, 127, -103, 114, -128, -128, -128, -128, 127, 108, 127, 127, 122, -81, 107, 43, -128, 127, -44, 127, -59, 23, 127, -50, 127, 97, -128, -91, 88, -74, 127, 127, 127, 127, 127, 127, 127, 22, 127, -128, 127, -128, -15, 0, -53, 127, 118, 15, -128, -128, -128, -128, -117, -128, 43, -1, -128, 127, -128, 106, -121, 66, 44, 127, 127, 127, 127, 127, 127, -38, 127, 7, 107, 127, 127, -49, 48, 127, -79, 127, -60, 52, -45, -128, 127, 127, 100, 127, -128, -65, -128, 1, 127, 31, 1, -128, -128, -121, -128, -128, 127, -128, -128, -128, -128, 127, 127, -86, 127, -2, -121, -128, 108, -79, -128, 127, -128, -128, 127, -128, 16, -128, -128, -128, -128, 107, 92, 49, 50, 127, -128, 127, -50, -128, 127, -10, 127, 127, -128, -2, -128, -128, 127, -128, 111, 127, -65, 49, -55, 114, 127, -74, -26, 118, -71, 122, 127, 127, -128, -128, 43, -37, 127, 127, 32, -128, -128, -100, 114, 127, 127, 127, 127, 127, -52, 37, -124, -128, -95, 80, 127, 111, -81, -108, -128, -128, 12, -128, -73, -7, -128, 127, -23, -128, -128, -128, -128, -57, 127, 127, -60, -113, -128, 32, 38, 95, 127, 101, 31, 127, 127, -78, -38, 57, -128, 127, 127, 127, 127, -38, -50, 0, -97, 13, -47, 11, 127, 127, -63, 27, -128, -49, 127, -128, 71, -128, -128, 42, 78, 127, 127, -3, -43, -128, -48, 0, -128, 97, -128, -128, -128, -128, -128, 27, 101, 12, -26, -128, -91, -128, 45, 114, 60, 106, -23, -78, 127, 80, 34, -76, -128, -127, -128, -117, -128, -128, -111, 127, 63, -23, 127, -3, -5, 127, 93, -16, -128, -128, -128, 11, -10, -113, -128, -123, -128, 29, 127, 127, -42, 64, -33, 127, 127, -128, 127, -70, -128, -74, -128, -128, -128, -128, -68, 24, 95, 127, -38, 70, 127, 127, 127, -28, -37, -69, 123, -32, 127, -108, -128, -128, -128, -128, -66, -128, -29, 38, 86, 127, 127, -93, 127, -128, 127, 53, 127, -128, -128, 127, 127, 127, 18, -57, -128, -128, -128, -128, -98, -21, -128, 27, -128, -128, -128, -128, 47, 127, 127, 91, 92, -128, -128, 36, -86, 22, -128, 2, -128, -128, 127, -88, 127, -26, -128, -118, 85, -31, 127, 127, -22, -128, -16, -128, -128, 6, 17, -128, -111, -119, -128, -68, 127, 109, -22, 87, 68, -128, -128, -74, 112, -52, 106, 127, -122, -128, -92, -128, -128, 127, -128, 127, -128, -58, 127, -112, 127, -128, -53, 111, 127, 127, 2, -128, -128, -55, -116, -128, 102, -128, -101, 127, -74, 127, 127, -128, -87, 28, -116, 28, 127, 90, 127, 90, -112, 17, -128, 2, -128, -128, 103, 127, 127, -43, 58, -128, -128, 127, -128, 127, -128, 54, -45, -128, -80, -128, -128, -128, -59, 127, 127, 127, -128, 57, -107, -128, 127, 127, 127, 127, 100, -68, -24, -128, 127, 127, -128, 127, -128, -128, 127, -128, 127, -128, -21, -5, 17, 127, 127, 124, 127, 71, -106, 26, -128, 0, -128, -128, -92, -128, -2, -128, -128, -85, -117, 127, 127, 10, -128, -68, -128, -128, 127, -128, 127, -21, 127, 127, 127, 6, -128, -128, -55, -24, 79, 127, 127, -128, 79, -71, 127, 127, 127, -128, -81, -71, -128, 95, -128, 127, 111, -79, -128, -128, -128, 88, 127, 127, 127, -128, -128, -47, 27, 127, 0, -36, -43, -128, 127, 28, -31, -128, -128, -23, 68, -15, -112, 38, 127, -36, 90, 127, -128, -15, 117, -3, 127, -107, 127, 13, -128, -43, -128, 2, -33, -128, 73, 52, -128, -42, -79, -128, 34, 127, 127, 127, 127, -81, 127, -128, 57, 48, 74, 127, -74, 87, 88, 127, 127, 57, 127, 127, -23, 127, -78, 127, 21, 54, 127, -48, 127, 102, 42, -13, -36, 127, 127, 86, 52, 127, -86, 127, 38, 76, -57, -49, 116, -73, 127, 127, -128, 86, -128, -26, -128, -128, 127, 57, -128, 127, 7, 127, 127, 127, -59, -128, -128, -128, 127, 127, 119, -122, -128, -128, -24, 127, 0, 127, 127, -79, 127, -32, 127, 93, -128, 127, 71, -121, 113, -128, -128, 127, -128, 127, 127, -128, 127, 11, 127, 86, 80, 96, -22, -128, -3, 127, -7, -74, -54, 127, -18, 127, -27, -128, -128, -128, -5, -128, -45, 127, 11, 127, 127, 58, 127, 127, 127, 111, 127, -27, -128, -128, 127, 98, 127, 127, -128, -65, -128, -128, -79, -8, 5, 0, -59, -128, -69, -87, 127, -98, 127, 127, -128, 68, -76, -128, 127, -64, 127, 100, -128, -78, -128, 58, -128, -128, 127, -63, -36, 127, 15, 127, 102, 95, -128, 60, -128, -31, 127, 50, 73, 127, -128, -128, 49, -112, 127, 127, -23, 34, -128, -128, 127, -128, 113, 109, 127, 127, 127, -13, -128, 118, 127, 127, 127, -128, 127, 102, -97, 54, 127, 44, 95, 111, -128, 127, 3, -74, 123, 127, -49, 127, 121, 127, 57, 127, 127, 127, 107, -64, -95, -36, 127, 127, 127, 127, -65, -117, -128, -21, 70, -54, 127, 2, 122, 127, 45, 127, -8, -128, -50, -124, -16, 127, -54, 112, 127, -113, 127, -128, -16, -128, 52, 127, -21, 127, -60, -128, -128, -128, -128, -128, 127, 118, -118, -80, 103, -85, 127, 85, 26, -22, -55, -128, -93, -69, 3, -128, -38, 127, -80, 127, 127, -128, 50, -128, -128, 127, 127, 127, 127, -52, 127, -128, -128, 106, -128, 122, -85, 93, 127, -128, -128, -111, 93, -128, 87, -128, -128, 68, 12, -10, 127, -128, -128, 127, -37, -98, -65, -128, -93, 0, -128, 127, 127, -91, -128, 52, -128, -128, -128, -128, 101, 127, 34, 127, -128, 33, 78, -124, 86, -128, -60, -128, 127, 127, 127, -58, 127, -28, -128, -128, -128, 127, -128, 127, 91, -128, -122, -64, 24, 127, 127, 127, -65, -128, 76, 33, -113, -128, 7, -128, 34, -8, -128, -68, -98, -128, 24, 127, 127, 127, 100, -128, -116, -128, 28, 101, 8, 127, -74, 127, 116, -128, 23, 116, -91, 127, 111, -13, 12, 116, 127, 127, 39, 127, 17, -128, -128, -74, -128, -128, -128, -128, 95, 127, 127, 90, 127, 127, -128, 127, -128, -128, 127, 127, 127, 85, -28, 10, 98, -55, -17, -128, -128, -128, 80, 127, -74, 60, -128, 127, 54, 11, 127, -90, -128, 33, -68, 127, 127, -128, -64, -5, -128, 127, 127, -128, -128, -117, -47, 127, 127, 127, 127, -116, -128, -6, 38, -68, 73, 92, -128, -38, -128, -44, -128, 47, 47, 127, 127, -78, -128, -128, -128, -128, 127, 127, 127, 127, -73, 127, -78, -128, 127, -128, 60, -128, -128, 127, -119, 127, -54, -128, -128, -128, 47, -128, -128, 127, -128, -38, 127, 10, 127, 127, 127, 127, -21, 127, 127, -128, 127, -128, -70, 113, 127, 127, 127, 127, 127, 127, 127, 127, -128, -93, 127, 127, -73, 127, 124, -128, -29, 107, -90, 5, -49, -128, -114, -13, -57, -128, -23, -128, -128, -123, -3, -43, 117, 127, -128, 127, -93, 65, -128, 118, -54, -128, 71, -128, -101, 50, -128, 127, 75, 27, 127, -128, 127, 74, -128, -32, -128, -128, -74, -128, -128, 118, 127, 93, 91, 127, 1, -128, 127, -128, -128, 127, -128, 11, -16, -59, 0, -128, -11, -128, 21, 127, 127, 127, 127, -98, 73, -21, 11, 127, 98, -58, -28, -76, 127, -47, -124, 96, -103, 127, 127, -75, 127, -128, -128, 127, -128, 63, 127, 81, -2, 127, 127, -128, -92, 127, -128, -60, 127, -33, -112, 127, 127, 127, 57, -128, -128, -58, -128, 127, 124, 38, 127, 6, 66, 127, 74, -96, -23, -128, -100, 117, 127, 127, -128, -128, 127, -11, 100, -17, -128, -103, -128, -79, 127, -113, 127, 127, 127, 127, 127, 127, -13, -128, -128, -128, -128, -128, -93, -128, -128, 127, -128, 65, 127, 16, 48, 127, 127, 38, 127, -8, 50, -128, -43, 71, -128, -128, -10, 63, 127, 48, 127, -128, -38, 1, 31, -24, 92, 114, 1, 127, 117, 127, 97, -128, -128, -70, -128, -128, 29, -128, -128, -128, -128, 127, 127, -128, 127, -128, 17, 127, -21, 0, -33, -128, -57, -114, -128, 127, 114, 127, -59, -128, -15, -106, -12, 10, -128, -124, 127, -128, 127, 127, -128, -116, -55, -128, -95, -128, -128, -128, 55, -128, -96, 127, -128, 96, 127, 127, 127, 27, -128, -103, -128, 12, -21, 70, 33, 127, 127, 127, 127, -26, 127, -85, -128, 38, 127, 127, 127, 127, -128, 127, -128, 121, 21, -128, 127, -80, 71, -128, -90, 81, -128, -128, 3, -128, -54, 127, 38, 33, 127, -128, -50, -128, -128, 92, 79, 127, 127, -5, 127, 11, -128, -78, -128, -128, -128, 78, 127, -28, 49, -128, -128, -128, -128, 127, -38, -24, 127, -101, -128, 127, -128, 127, 127, -128, -128, -123, -116, -128, 127, -128, -116, 127, 127, -11, 93, -39, 127, -21, -45, 127, 101, 127, 127, -16, -88, 75, -128, 33, 24, 127, 116, -106, 127, 127, 91, 107, 127, -128, -128, 127, -128, -38, 127, -117, 127, 127, 10, 13, -111, -128, -128, -128, -128, -16, -26, -128, 74, -93, -102, -128, -128, -128, -128, -128, -128, -128, -45, -68, 81, 127, 93, -128, 57, -128, -128, 127, -59, 127, -2, -17, 127, -128, -38, -108, -128, 127, 127, 127, 127, -128, -128, 45, 74, 127, 91, -116, -128, -128, -128, -58, 127, 127, 127, 127, -1, -95, -128, -128, -128, -128, -50, -128, 10, 71, 127, 127, 117, -74, -109, 127, 127, 127, -113, -97, -128, 127, -85, -44, 127, -128, 127, -109, -98, -91, -91, -128, -128, -128, -81, -64, -128, -57, 18, -95, 127, 127, 127, 52, 127, 127, -102, 127, 37, -128, -128, -128, -128, -23, -128, 57, 69, -48, -48, -90, 109, 127, -128, 57, 102, -112, 127, 5, -128, 95, -128, -128, -128, 127, 57, -85, -128, 50, -18, -113, -50, -128, -128, -49, -128, -17, 34, 8, 127, 127, -22, -5, -128, -128, -128, -12, -97, -128, -128, -128, 127, 45, 65, 95, -128, 114, -128, 124, -75, 86, 127, -128, 87, -128, -128, -128, -128, -128, -128, 127, 127, 127, -22, 24, -128, -128, 127, -31, -96, -26, -128, -128, -13, -71, -18, 121, 127, 127, 127, 1, 34, -17, -74, 127, 111, 127, 127, 103, 127, 127, -59, 127, -128, 0, -128, -128, 0, -11, 127, 127, 127, 127, 58, -128, -128, -128, -128, -90, -100, -31, 127, -121, 127, 85, -128, 127, -128, -92, -128, -116, 79, 49, 127, 127, 127, -36, 127, 127, -128, 127, 127, -53, 24, -128, -128, -22, -128, -128, 81, 127, -98, 69, 101, 95, 127, 127, 127, 127, -7, 127, -121, 127, 102, -128, -128, -128, -128, 114, -60, 49, 127, -128, 43, -128, 57, -121, 127, 63, -128, -128, -106, -128, -68, 127, 127, -16, 127, 111, 121, 127, 0, -128, -64, -128, -128, 23, 58, -128, -63, -80, -128, 78, 86, 127, 127, 127, 96, 127, 74, 127, -128, 49, -79, -128, -128, 11, -128, -64, 127, -128, -43, -47, -128, -100, 127, -128, 127, 12, 12, 127, 127, -26, -45, 127, -128, -7, 43, 37, 69, -70, -87, -57, -111, -128, -128, -109, 127, 127, 127, 127, -1, -128, -128, -29, -128, 127, -128, -128, 127, -128, -6, -22, -66, 127, 96, 127, 127, -128, 127, -85, 49, 127, 31, 127, 127, -128, 127, -128, 127, -1, 10, 81, -128, -95, -128, -128, -81, 50, 127, 127, 127, -2, 124, 5, -128, -128, -128, -17, 45, 127, 127, 79, 127, 26, -128, -59, -49, -71, 111, 127, 114, -128, 88, -128, -128, -63, -128, -128, -128, 3, 10, -128, 38, -128, -128, -128, -128, -128, -128, -124, -117, 39, -34, -8, -128, -128, -128, -128, 93, -128, 127, -106, -7, -37, -128, 127, -90, 127, 31, -128, -128, 38, -85, 127, 127, 127, 127, 79, 124, 127, 127, -128, 127, -123, -79, -128, 58, -128, -81, 127, 127, 78, -31, -27, -128, -128, -128, -128, -128, -128, 127, -128, 127, 127, -85, 38, -128, 26, -116, -128, 75, -128, -128, -69, -128, -128, -128, -128, -39, -54, -42, 127, -128, -44, 127, -128, 127, 127, 127, 127, -73, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 47, -128, -128, 127, -128, -50, 33, 127, 127, -117, 127, 127, -128, 127, 6, -128, -57, -128, -128, -121, 127, 127, 127, 127, 127, 127, 127, -128, -93, 23, -22, -36, 24, 57, -128, 127, -10, 127, -68, -70, -128, -128, 127, 44, 121, 127, -128, -128, 86, 127, 127, 127, 109, -128, 91, -128, 0, 127, 33, 15, 23, 100, -128, 127, -128, -128, 116, -128, 106, 127, -98, 124, 85, -128, 127, 127, -128, 127, -128, -128, -128, -128, 127, -21, 73, -128, 53, -63, -128, -128, -128, 85, 127, 127, 127, 117, 127, -128, -36, -49, -34, 127, 127, -39, 127, 127, 123, 127, 93, 45, 127, 127, 127, 127, 127, 98, 127, -37, -128, -128, 119, -128, 127, -66, -128, 90, 127, 65, -80, 127, -122, 122, 127, -128, -48, 60, -128, 36, -128, -1, -123, -128, -112, -53, -47, 127, 102, -121, 32, -128, -74, 5, -47, -128, -128, -128, -128, -63, 127, 127, -128, 127, -123, -128, 127, -128, -128, 127, -128, 127, 127, -128, 22, 26, 127, -15, -101, -23, 85, 93, -44, -128, 26, -128, -128, -128, 1, -128, 57, -21, -128, 127, -88, -68, 127, 28, -13, 127, 117, -106, 43, -128, -59, -128, 87, 127, -128, -96, -128, -128, 37, 127, 59, 52, -6, -128, -128, -128, 127, 74, 127, -128, -128, -128, 73, -50, 127, -11, -128, 127, -128, 43, -109, -128, -22, -128, 127, 127, 10, -128, -13, -128, -128, -128, -6, -128, 111, -71, -128, 127, 111, 127, 127, 127, 127, 127, 127, 127, -128, -5, -63, -128, -53, -128, -128, 127, 127, 127, 127, 127, 16, 127, -128, 100, -128, -128, -39, -1, 127, -128, 95, 127, 121, 127, 58, -128, -128, -128, 48, 127, -47, 127, -54, -128, 127, -1, -128, 16, -128, 48, -128, 127, -58, -7, -3, -98, 127, 24, 33, 1, 127, -85, -119, -38, 127, -18, -78, 127, -8, -128, 103, -106, -21, -128, 119, -128, 127, 127, 31, 27, -128, -37, -127, -128, 127, -33, 23, -128, -128, -128, 22, -128, 127, -45, -78, 127, 127, 55, 127, -54, -128, -128, -128, -128, -128, -128, -128, -128, -128, 54, -100, 68, -27, -24, -128, 127, -2, 33, 66, 107, 127, -42, 127, -53, -128, -128, 107, -128, 127, 86, -124, -128, -128, -58, -128, 85, -27, 16, 127, 127, 127, -128, -113, 65, -100, 127, 127, -128, 124, 127, -91, 127, -69, 3, 127, 127, 108, -17, 21, -93, 127, 127, 114, 86, -113, -128, 127, -81, 127, 24, 65, -75, 63, -96, 92, 43, -52, 127, 127, 127, 127, -128, -128, 124, -106, 5, 127, -128, 100, 127, -3, -128, -55, -109, 64, 127, 127, 85, 127, -63, -128, 127, -117, 34, -42, -128, 127, 76, 58, -28, -128, -128, -128, -128, -128, -91, -128, -128, -45, -128, 127, -2, -5, -36, -128, -59, -86, -117, -128, -128, -128, -128, -59, 98, -73, 127, -124, 127, 15, -98, -97, -128, 127, -128, 127, 127, -18, 113, -128, -128, 127, -112, 95, -12, -128, 127, 127, 127, 16, -79, -3, -97, 127, -128, 64, -128, -54, 127, -128, 127, -58, -128, -23, 127, 127, 75, -128, -116, -39, -128, 27, 100, 12, 58, 5, -128, -119, 127, 127, 127, 127, 16, 127, 127, 127, 127, 127, 127, 101, 127, 100, -128, -70, 127, 127, 119, -63, -128, -128, -111, 127, 127, -15, 5, -128, -93, 106, 78, -92, -128, 57, -11, -111, -128, -128, -96, 37, -5, -128, -128, -24, -128, 127, 127, -93, 107, -128, -96, -128, 127, 127, 127, 127, -128, -27, -54, 43, -128, 121, 11, 0, 6, 127, -75, -74, 119, -128, -128, 2, -128, -128, 127, 11, -128, -34, 93, -128, 1, 100, 127, 127, -85, -12, -128, -128, 127, -59, 127, -128, -128, 127, -128, -128, -128, -128, -121, 69, 127, 127, 117, -92, 78, -128, -59, 127, 54, 127, -128, -124, 55, -13, 57, -128, -76, -91, 127, 127, 10, 127, -80, 127, 127, -128, -128, 18, -16, -127, 59, 0, -128, -78, -59, 127, 127, 127, -128, -128, -81, -128, -60, 127, 73, 127, 127, 18, 42, -128, -63, -1, -128, -128, -128, 1, -128, 127, -52, -128, 127, 33, -128, -85, 127, 24, -93, 111, -26, -69, 127, 21, -39, -128, -128, -128, -59, -128, -128, 55, -73, -128, 43, -52, 16, 127, -55, -128, 101, -128, 127, 127, 43, 127, -5, -128, 0, -128, -128, 108, 127, 68, 127, 127, -76, -128, -128, -128, 81, 75, 127, 127, -128, -128, -24, 127, 127, 127, 127, 78, -128, 127, -118, -128, -111, -69, -81, 127, -128, -109, -128, 0, 127, 52, -128, -128, -128, -12, 127, 10, 127, 127, 87, 127, 127, -8, -91, -128, 87, 127, 127, -57, 127, -16, -37, -31, -128, -128, -128, -128, 127, -128, 24, 127, -18, -128, 73, 44, -111, -128, 66, -128, -128, 70, -128, -113, -128, -128, -95, 0, -128, 33, -128, -128, 127, -128, -128, 74, -128, -107, -95, -124, -128, -128, -57, 29, -7, -114, 113, -128, -33, 127, -64, 127, -7, 36, 124, -128, -12, -128, -128, -128, -128, -114, -118, -73, 16, 127, -128, -38, -55, 127, 127, -128, 17, -11, 127, 127, 127, 127, 85, 127, 66, -45, 57, -128, -128, 81, -128, -48, 127, 15, 80, 127, -128, -92, -27, 127, 88, 127, -24, 97, -12, -11, 127, -107, 37, 127, -103, 29, 80, 127, 127, 127, 18, -128, 127, 0, -96, -128, 22, -128, 100, 127, -128, -58, -128, -128, 13, 127, 127, -98, 117, -128, 8, -124, -71, 127, -52, 127, 127, 127, 127, 123, 39, -128, -128, -128, -128, -117, 127, 114, 127, 127, 127, 29, 127, 32, -128, -128, -128, -59, 127, 127, -128, -28, -95, 127, 127, -63, 127, -128, -128, 17, -128, -124, 87, -128, 71, -78, -128, -128, -95, -93, 75, -29, -103, -101, -128, -128, -128, 55, 13, 127, 127, -13, 127, 60, -128, -5, -128, 78, 127, 87, 127, -68, 127, -128, 28, 28, -128, 127, -106, -128, 127, -128, 127, 42, 127, 49, -123, -28, -128, -64, 79, 33, -128, 76, -128, -128, 127, -65, 70, -98, -128, -128, -128, -69, 117, -37, 16, -15, 127, 127, -55, 48, 127, -128, 127, 47, 0, -31, 60, -100, -128, -128, -128, -52, -128, -69, -128, -128, -42, 127, 127, -21, -128, -37, -128, -128, 121, -3, 127, 91, -128, 11, 66, -128, 93, -114, 26, -13, -114, -21, -128, -63, -65, -128, 16, 1, -128, 127, -44, -28, -85, -111, -108, -128, -27, -128, -106, 57, 88, 58, -128, -128, -71, -128, -123, -128, -128, -128, 113, -1, -128, 127, -107, -75, 106, -128, -128, -128, -128, -128, -107, -128, -49, -29, 33, 127, -3, 127, 108, -128, 127, -64, -128, 80, 127, -128, 24, 59, -128, 127, 127, 127, 127, 49, 127, -102, 127, -78, -128, 127, -63, 76, 31, -90, 100, 127, -49, -60, -107, -54, 58, 127, 127, -128, -128, -128, -57, -128, 127, -128, 53, -64, 113, 127, -66, 0, -128, -128, -127, -10, 100, 127, -42, 75, 127, 127, 127, -6, 127, -128, 22, 127, 127, -69, 127, -128, -128, -128, -128, -128, 71, 127, 127, -68, -128, -95, 127, 127, -128, 127, -128, -43, 127, 66, 127, 127, 127, 127, 127, 1, -63, -3, -128, -128, -128, -128, 127, 107, 127, -128, 33, -128, 21, 127, -128, 127, -128, -128, -108, 10, 127, 127, 127, 112, -128, -128, 127, -128, 127, 127, -128, -128, -128, -128, -128, 127, 50, 113, 50, -128, 127, -128, 127, -113, -127, 55, -128, 127, 57, -128, 127, -13, -80, 127, -10, 11, 48, -128, -48, -128, -128, -128, -58, -111, 127, 127, -128, -48, 127, -128, 127, 127, -128, 127, 127, -57, -128, -128, -121, -54, -73, -128, -128, -128, 28, 127, 1, 24, -128, -128, 103, 76, 127, 127, 127, 108, -128, -128, -24, -10, 127, 0, 39, 127, -15, 6, 127, 23, -128, -3, 127, -21, 127, 127, -128, -57, -128, 80, 127, 127, 127, 127, 47, -128, 127, -128, -114, 11, 127, 127, 18, 32, 127, -128, 127, 127, -128, 127, -128, 127, 102, -128, 107, 127, 123, 122, -128, -128, -98, -128, 64, 36, -128, -128, -128, -128, -128, -128, -27, -128, -128, 95, -128, 127, 127, -128, 76, 127, 127, -73, 17, -128, -108, 117, -81, -38, 49, 7, 127, 127, -128, -128, 100, -128, 127, 57, -128, -87, -128, -128, -39, 36, 127, -16, 31, -69, -128, -6, -128, -34, -128, 43, -34, -128, 127, -107, -128, 127, 18, -128, -117, 0, -128, -18, 127, 127, 43, -128, -128, -106, -128, 98, 127, -128, -6, -128, -128, 5, 127, -128, 0, 127, -122, 127, -27, -128, 127, -78, 127, 127, -128, 127, -128, 114, -106, -128, 127, -128, -44, 122, 127, -16, 127, -74, -128, 127, -128, 127, 127, -128, -12, -106, 118, 127, 127, 112, -128, -128, 74, 68, 127, 127, 2, 127, 127, -128, -128, -128, 55, 127, 50, 127, -128, -15, 127, 90, 127, 127, -128, 127, -128, -36, -28, -128, 127, -128, -98, 73, 74, -128, 108, 127, -128, 127, -128, -88, 33, -70, -128, -128, -128, -128, -128, -18, 127, 75, 15, -128, -128, -128, -128, 127, -43, -87, 95, -128, -10, -75, -128, -128, 119, -16, 49, 127, -13, -128, -1, -36, 127, 95, -128, -33, -97, 108, 127, -87, 23, 127, 45, 124, -95, -128, -128, -128, -128, -128, -128, -128, -97, 127, -128, 50, 124, -17, -27, 127, -18, -128, 93, -107, -128, -128, -66, -37, 101, 127, 127, 127, -26, 127, 127, -128, 127, -128, 33, 18, -128, 109, -128, -128, 42, 127, 65, 127, 127, -3, 127, 127, 86, -92, -128, -55, -128, -49, -128, -74, -128, -112, -66, -128, 127, 0, -34, 55, -70, 55, -55, -117, 127, 127, 47, 127, -128, 16, -128, 13, 127, -93, 127, -8, -128, 127, -128, -128, 127, -128, 127, -128, 24, -52, -12, 127, -128, 127, 127, -128, 127, -128, -68, 58, 102, 127, 127, -128, 127, -128, 36, 127, -128, 37, -128, -21, 90, -47, -128, -128, 113, 66, 127, 127, -108, -70, -128, -128, 127, 42, 127, -128, -58, -128, -128, 127, -90, 127, 127, -128, 127, -128, 127, -5, 22, 69, -128, -128, -123, -49, -52, 66, -128, -1, 127, -114, 127, -102, 98, -23, 127, 127, 48, 78, -128, -128, -128, -128, 17, -96, 127, 121, -28, 79, -128, 5, -122, -128, -26, -128, -128, -128, 24, 21, 127, -69, 55, 127, 127, -70, -23, 127, -65, 127, -128, 8, -128, 127, 127, -128, 127, 12, -50, 127, 127, -128, 127, 127, -43, 29, -128, -75, -128, 127, 57, -98, 85, -128, 70, -1, -128, -128, -128, -53, 127, 127, 127, 37, 44, -37, -38, 127, 127, 55, 48, -128, 92, -128, 127, 127, -128, 127, -128, -128, 107, -128, 127, 116, -70, -128, 127, -128, -45, 127, -128, 127, 127, -128, 127, 127, -117, -90, 64, -128, 27, 127, -68, 33, -111, -128, -128, -128, 48, -76, 127, -128, 127, -128, -127, 127, -117, -128, -63, 28, -93, 127, 2, 11, 81, -128, -2, 66, 42, 64, -128, -80, -128, -59, 3, -34, 127, 78, -127, 81, -60, -128, 49, -128, 65, 10, -12, 127, 22, 111, 29, -128, -128, 127, -87, 127, -15, -22, -128, -128, 108, -50, -128, 127, -59, -128, -128, -128, 0, 59, 127, 93, -3, 127, -128, 127, -21, 127, 127, 26, 76, -34, -128, 58, -57, -128, 44, -15, -128, -117, 53, 127, 127, 127, 127, 127, -76, 127, -128, 127, -100, 127, 44, 10, -128, -75, 127, 103, 11, -128, -87, -128, 127, 127, -106, 127, 127, 22, -36, -75, -128, -128, -128, -76, -1, 127, -128, 127, -128, -128, 127, -128, 45, 127, 43, 127, 127, -102, -128, -128, -55, -128, -42, -22, -128, 55, -128, -128, 127, -128, 63, -128, -128, -128, -128, 74, -8, 127, 127, -128, 12, -75, 127, 127, 47, 63, 127, 127, 127, 109, -103, -128, -128, -128, -128, -128, 92, -128, -128, 36, 127, 127, -128, -78, -29, 127, 127, 127, -128, -116, -49, -128, 60, -128, 127, 127, -128, 127, -128, -111, 127, -68, -63, 127, 32, 81, 48, -128, -128, -128, -128, -128, -128, -128, -128, -128, -27, 127, -8, 127, 95, 22, -29, 127, 111, 3, 127, -128, 127, 127, -103, -128, 49, -128, 127, 127, -128, -7, -12, -53, -68, -128, -128, -128, -128, 127, 127, 127, 127, 85, -128, -64, -128, -69, 127, -128, 7, -128, -55, 107, 127, 127, 127, -128, 127, -128, -128, -10, 58, -128, 127, -79, -42, 127, 98, 58, 127, 127, 127, 127, -66, -128, 109, -128, -121, 127, 32, -27, -128, 26, -128, 101, 127, -128, -128, -71, -128, -128, 127, -128, -49, -33, -128, 127, 127, 127, 127, 114, -128, 127, 76, -124, -128, 24, 93, -128, 127, -23, -58, 127, 127, 127, 127, 127, -128, 127, 13, -73, 127, 85, -32, 127, -128, -128, 127, 48, 111, 127, -128, 101, -11, -128, 127, -128, -17, -128, -128, 127, 127, -85, 127, 127, -128, 127, -128, -124, 127, 127, 127, 127, -128, -28, 12, -128, 127, -128, -58, 127, -128, 127, 127, -87, 127, 5, -112, 103, -34, -128, 37, 127, 54, -37, -97, -128, -111, -95, 127, 86, 127, -128, -128, -26, 127, 127, 127, 127, -128, -128, -128, -128, -128, -107, 119, -70, 127, 21, 127, -74, 127, -128, 0, 113, -128, -128, 64, -128, 90, 127, -112, -128, -78, -128, 127, 127, -3, 127, -53, 65, 127, 127, -29, 48, -96, 127, -42, 127, 127, -128, 127, -122, -128, 63, -49, 127, 127, -128, 15, 127, -88, 127, 108, 13, -18, 114, -86, -128, 114, -128, 2, 127, 127, 127, 55, -55, 27, -128, -128, -103, -76, -128, -128, -36, -73, -128, -128, -128, -53, 127, 127, 32, 127, -128, -107, -128, -48, -64, -128, -128, -128, -128, -128, 32, -128, -128, -32, 70, 26, -68, 127, -128, -68, -10, 127, 127, -24, -93, 97, -128, 60, -57, -80, 127, -128, 127, 127, -128, 127, -96, 1, 127, -128, -1, 127, 10, -128, -28, -128, -93, -127, 127, -128, 127, 109, 127, 127, -100, 127, -63, 127, 127, -128, -49, -128, -128, -128, 15, -47, -128, 127, -128, 122, 52, -128, 59, -38, -128, -16, -128, -128, 31, -128, -128, 5, -128, -128, 1, 127, 127, 127, -74, 52, -107, -128, 97, 123, -113, 127, -128, 113, -21, 122, 127, 26, 127, 127, 127, -34, 27, 7, -44, 127, -8, -128, 21, 71, -1, -38, -128, -128, -128, -124, 127, -103, 127, 127, 31, 127, 127, 117, -128, -128, 127, 59, 127, 24, -128, -128, -128, -21, -48, -128, 127, -42, 127, 127, -42, 55, 127, 127, -37, 122, -128, -128, -7, 75, 114, 127, 127, 91, 127, -3, -113, -128, -121, 96, 48, -47, -78, 114, 127, 71, 127, -128, 127, 127, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, 127, 38, 107, -128, -128, -128, -128, 127, 127, 127, -128, 16, -128, -128, 100, 127, 127, -42, 127, 127, 87, 85, 127, 117, 127, -128, -39, -128, -10, -36, -128, -128, -59, 50, -128, -128, 127, -29, -128, 127, -128, 76, 127, -101, -128, -128, 45, -75, -44, -128, -128, 10, -128, -128, -128, 0, -128, -87, 127, -23, 127, 58, 127, 127, 127, 101, -128, -38, -128, -31, 31, 116, 127, 2, 24, -85, -128, -128, -107, -128, 33, -28, -11, -128, -64, 3, 47, -128, 117, 127, -128, 123, 127, -128, 127, -128, -128, 127, 127, 127, -86, 2, 34, -128, 127, 127, -128, 127, 127, -128, 127, 80, -122, -128, -128, 27, -128, 107, 127, -128, 127, -114, -128, 127, -128, 127, 127, 127, 97, -33, -24, -128, -128, 127, 0, -128, -2, -128, -128, 127, 127, 127, 127, 127, -128, -5, -128, -54, 112, -128, -55, 101, 44, 127, 36, -8, 102, -79, 127, 92, -13, 127, 127, 121, 127, -128, -128, 127, -128, 23, 127, 91, 127, 76, -128, -128, 10, 127, 13, 127, -18, 127, 127, -128, -128, 26, -37, 127, 127, 42, 100, 113, 123, 127, 114, 127, 47, -128, -128, 29, -128, -34, -81, -128, -128, -7, -96, 127, 73, -128, -128, -21, -128, -128, 127, -128, 127, 80, 127, 127, -88, 127, -128, -128, 29, 45, 127, 127, -3, 127, -128, -128, 127, 34, -128, 127, -7, 95, 127, -24, 127, 127, 127, 86, 127, -75, 29, 81, -111, 127, 8, 127, -55, -86, -128, -128, -128, -23, -50, -31, -69, -128, 127, -113, 127, 127, 127, 22, 127, 28, 97, -128, -111, 127, 5, 44, 42, 127, 127, 127, 0, -91, 127, -128, -53, 127, -128, 127, 127, -128, 127, 113, -128, -36, -95, -128, -106, 58, 127, 101, 127, 127, 127, 68, -87, -100, 33, -39, -18, -128, -91, -55, 127, 127, 127, 127, 68, -39, -128, -128, -57, 97, 127, -128, 127, -128, -96, 44, 68, 127, -128, 109, -128, -128, -128, -37, -128, 116, 92, 127, -12, -8, 27, -128, 34, -128, -128, -71, -128, 42, -128, 127, -128, 124, 127, -128, 71, -128, -128, -128, 106, -128, 127, 18, -128, -128, -128, 18, -128, 127, 127, 117, 127, 111, -128, 127, -128, -54, 127, 33, 127, 127, 127, -13, 88, -128, -81, -16, -128, 39, 127, 106, -78, 127, -112, -97, 91, 127, 127, 101, 127, 23, -128, -58, -65, 127, 127, 127, -6, -121, 127, -128, -107, -128, -128, 127, 63, 127, 102, -128, -128, -16, -128, -96, 127, -128, 98, -33, 7, 116, -112, 127, -47, 107, -42, -128, -21, -128, -75, -24, -118, 127, -86, -128, 117, 113, -117, -50, -128, -128, -16, -27, 49, 13, 127, 1, 127, 34, -128, 98, -128, -60, 80, 127, 127, -90, -128, -92, -128, 122, -5, -128, 127, -49, 127, 127, 96, 127, 127, -128, 12, 42, -128, -128, 64, -128, -128, 127, 108, 106, -128, -117, -128, -128, -69, -2, -128, -70, -97, -65, -114, -128, -128, -128, 109, -107, -124, -128, -95, -128, 127, 106, 127, 93, 96, -128, -128, 24, -47, 127, -127, -128, 34, -128, 111, -44, -26, 127, 127, -70, 127, -128, -118, 127, 22, 127, 127, -1, -55, -76, -128, -10, -128, -128, 127, -113, -128, -128, -128, -128, 127, 71, 96, -78, -128, -128, 102, -71, -128, -92, -128, -128, 0, -128, -78, -8, 102, 127, 127, 127, 123, 127, 127, 8, -128, -106, -128, 127, 127, -128, -79, 96, -21, -128, -16, -34, -128, 127, -97, 5, 127, 127, 127, -23, -128, -90, -128, -128, 127, -128, 97, 81, 12, 127, 127, 119, -128, -29, -128, -116, -128, -128, 28, 10, -128, -23, 74, -10, 127, -128, -16, -128, 58, 127, 78, 127, 127, 127, 127, -63, 64, -128, -32, 127, 127, 127, 18, 36, -45, 127, 127, 127, 121, -128, 127, -118, 127, 127, 64, 127, -114, -92, -128, -128, -128, -128, -116, -128, 71, -128, 127, -60, -128, -128, -73, 127, 127, 127, 127, 17, -85, 127, 93, -66, -128, -128, 12, -128, 39, 127, -113, 26, -128, -28, -128, 121, 127, -43, -75, -55, -128, -128, -128, 127, 95, 68, 97, -128, -113, -128, -128, -128, -128, -128, 122, -52, 127, 112, 26, 127, 127, -23, 127, -128, 86, -128, -6, 127, -128, 127, -48, 57, 127, 0, 127, -80, -123, 58, -81, 127, -128, -85, 127, 24, 127, 127, -90, -27, -128, -55, -128, -44, 127, 96, -128, -121, -13, -73, 23, 127, -98, 6, -60, -32, 48, 127, 48, -128, -128, 127, -15, 88, -122, -128, 58, -2, -128, 90, -128, -128, 127, -118, -128, 127, 74, -71, 127, -128, 127, 37, -128, -38, -128, -95, -128, -128, -128, -48, -128, -128, -128, 33, 52, -128, -128, -128, -116, -103, 73, -128, 127, -128, 127, 33, -128, -111, -128, 127, 121, 70, -73, -128, -128, -128, 106, -128, 13, -114, -128, 127, -128, 32, -78, 87, -128, 127, -10, -128, -128, -122, -18, 127, -17, 127, 32, 127, 127, -128, 85, -128, 127, 2, 127, 57, -44, 127, -128, 101, 127, -101, -53, 98, -93, -128, -31, 2, -10, 60, -128, -128, -26, 127, 113, 127, -116, 12, -128, 45, 127, 108, -116, -128, 127, -128, 127, 66, 127, 92, -100, -128, -128, -128, -128, -128, -128, -57, -128, -16, 127, -128, 127, 78, -128, 127, -109, -128, 69, -128, 87, 127, 59, 127, 127, 102, -128, 13, -50, -11, 127, 127, 127, 127, -53, 87, -128, 31, -128, -128, 127, -88, 127, 127, 112, 127, 114, -128, -1, -128, -128, 34, -128, -128, -128, 7, -128, -128, -128, -128, 75, 127, -15, -128, -128, -128, -128, 127, 127, 127, 127, 127, 127, 127, 127, -8, 127, 127, 55, -128, 87, -128, 127, -112, 44, -128, -128, 85, 127, 127, -42, -60, -128, 63, 127, 127, -122, 127, -92, -16, 127, 127, 101, -109, -47, 127, -128, 127, -44, -1, 127, 118, 57, -128, -128, -128, 50, -128, 109, -33, -90, 112, -128, -128, 127, -49, -128, -128, -28, -124, 127, 127, 127, 127, 127, 127, 39, 127, 44, 127, -73, -128, -26, -128, -31, -92, -128, 11, 127, -128, 10, -22, 127, 127, 127, 16, 75, 81, 127, 127, -128, -16, -128, -48, 64, 69, 127, -29, 117, 127, 127, 127, 127, 127, 127, 127, 127, -11, 127, 127, -58, 127, -128, -128, -52, -128, 48, -128, -48, 127, 85, 65, -128, 28, -70, -128, -69, -128, -128, -128, -128, 127, 127, 2, 127, -128, -128, 127, -111, 101, 39, 76, 96, 127, -128, -2, 127, 127, 127, 6, -128, 21, -128, -81, 32, -128, -57, -128, -128, -39, -69, -128, 127, -86, -128, -12, -49, -128, 127, -128, -121, 127, -68, -6, 127, -128, 103, 127, -38, -91, -128, -93, -128, 85, -128, -5, -64, 127, 34, 127, -128, -128, 17, -128, 127, 127, 107, -128, 55, -114, -128, -93, 16, -128, 127, 127, -119, -128, 22, -128, -38, -128, -42, -118, 98, 127, 93, 127, 127, 55, 12, -70, -128, -128, 103, -128, 63, 86, 127, 127, 127, 8, -128, -128, -103, 127, 127, 127, 127, 127, 127, 127, 127, -128, -128, -74, -49, -70, -116, -128, -68, -128, 78, 33, 39, 127, 95, -71, -37, -128, -128, 36, -128, 107, 127, -32, 122, 127, -128, -50, 81, -92, -18, 127, -85, 39, -100, 102, 75, 2, 78, -128, -128, -8, 49, 93, -48, 54, 127, 127, 15, 127, 73, -128, -70, 90, -65, 116, -29, 127, -12, -69, 127, -128, -31, 127, 6, 127, -128, -76, 47, -106, 127, -69, 127, 127, -13, 127, -55, 127, 127, 127, 127, 127, 1, -63, 127, 127, 49, 1, -128, -13, -87, -128, 127, -128, -128, 127, 127, -8, 127, 127, -128, -13, 74, -128, 29, 127, -128, 70, 127, -128, 127, 47, -57, 12, -128, 47, -128, 69, 95, 80, 127, 127, 127, 127, 127, 100, -128, -87, -128, -128, 36, 127, 24, 93, -128, 113, -128, 127, -128, -128, 127, -128, 127, 127, -42, 127, 16, 107, -52, 127, 127, 12, 31, -119, -128, -112, -128, -128, -128, 28, 49, -128, 127, -128, 127, -116, 26, -128, -128, 16, 127, 127, 106, 85, -128, -48, -128, 54, -128, -28, -85, -112, -128, 123, -128, -78, 127, 85, 127, 127, 127, -86, -128, -73, 71, 18, -128, 64, -128, -59, -128, -49, -128, 12, 127, -8, 108, 45, -124, 52, -128, -68, 117, -128, 127, 123, -37, 31, -128, -128, -90, 58, 38, 127, -111, 127, 45, 127, 127, 127, -38, 31, -128, -128, 127, -59, 127, 127, 122, 127, 127, 127, 127, 91, 127, 127, 86, 127, 127, -123, 93, 127, 127, -26, 127, -128, -49, 127, -92, 127, 113, 127, -127, -78, -128, -128, -128, -128, -17, 112, -93, 127, 127, -97, 127, 127, -128, 127, 127, -60, 127, 114, -128, -128, -128, 127, 127, 127, 127, 66, -128, -121, 117, -128, 127, 53, -128, -128, -128, -128, 22, 8, 31, -102, -128, -128, -128, 48, 26, 127, 127, 27, 127, -13, 45, 127, 127, 74, 28, -23, 127, 73, 45, 103, 127, 11, 127, -128, -128, -21, -58, 127, 71, 127, 18, 127, 127, 119, 127, 0, 127, -114, 127, -43, 127, 10, -11, 31, -43, 3, 0, 127, 127, 127, 127, 127, -128, 31, -128, 0, 127, 127, -128, 127, -128, 127, 18, -128, 127, -128, 37, 1, -128, -128, -128, -128, -128, -128, -128, 11, -128, 127, 16, 66, 127, 124, 127, 88, 127, 127, 127, -48, 49, -128, -128, -58, 127, 127, 71, -22, -128, 3, -128, 74, 114, 7, -109, -50, -128, -128, -128, 47, 124, -128, 127, 60, 85, 127, 127, 127, -103, 127, 119, -128, -128, -128, 2, 2, 127, -27, 127, 11, 98, 63, -98, -52, 12, 60, 127, 127, 127, -128, 57, -128, -74, 44, -128, 107, -52, -128, -28, 8, -128, 0, -128, -128, -73, 127, 127, -49, 127, 75, -128, 127, -128, -128, 127, 127, -128, 127, -69, 23, -119, 127, 48, -128, -128, -128, -128, 127, 127, 127, 5, 52, -128, 100, 28, 127, 127, 127, -11, 5, 66, -128, 60, 127, -128, 127, -48, 55, 21, 123, 95, 111, 87, -95, 127, 36, 127, 107, 39, 2, -128, -1, 127, 127, 127, 127, -29, 127, 78, -128, 127, 1, -13, 54, 31, 127, 127, 127, -128, -95, 32, -39, 127, 23, 50, 127, -128, -88, -118, -128, 98, -128, -128, 127, -50, 127, -43, 127, -50, -128, 43, 127, 13, 58, 127, -88, 127, 117, -128, 17, -116, -78, -128, -54, -128, 103, 127, -11, -69, -128, -128, 73, -6, -128, 33, -128, -128, -128, -128, -128, -47, -15, -128, 63, -128, -128, -18, -128, -128, -128, -128, 63, -98, -128, 107, -128, -90, -128, 60, -69, 127, -88, -101, 127, -128, -1, 127, 54, -34, -122, 18, -128, -128, -122, -53, -128, 127, -128, -128, 127, 76, 127, -128, -48, -128, -128, 127, 127, 127, -60, 119, 127, -128, 127, 86, -128, 127, 39, -128, -128, -128, 112, 127, 11, 127, -128, 33, 13, -11, -128, -12, 102, 127, 127, 127, 127, 6, -128, -100, 127, -128, 127, 127, -36, 103, -128, -128, -116, -128, 58, -93, -128, -96, 38, 127, -86, -36, -54, -128, -27, -128, -128, -45, 47, -121, 127, -128, -128, 127, -54, 127, 28, -128, -122, -50, -128, 127, -101, 127, 127, -39, -128, -128, -45, -128, 127, 8, -36, 74, 55, -47, 101, -24, 127, 57, 127, 127, -15, 127, -128, 36, -92, -79, 97, -69, 127, 127, 127, -29, -44, -128, -128, -3, -68, 127, 113, 119, 26, 1, 127, -128, 50, 127, 68, 47, -128, -48, -44, 47, 102, 127, 74, 1, -128, -128, 16, -113, 127, 127, 127, 127, -128, -128, -111, 33, 127, 24, 79, 127, -16, -49, -100, -128, -112, 127, 16, -8, 127, -128, 127, -70, 127, 32, -128, 32, 127, 119, 100, 127, 108, 33, 127, 127, 127, 127, -128, -103, 17, -128, 127, 127, 36, 127, -128, -128, 127, -28, 127, 127, -39, 31, 127, 127, -111, 66, -128, 127, -7, 118, -128, -15, -128, -128, 127, -87, 127, 90, -53, 127, -117, 116, -128, -128, 57, -128, -106, 73, -128, 127, 53, -128, 127, -128, -128, 127, 127, 73, 127, 52, -79, 127, 127, 96, 80, -73, -128, 52, -128, -128, 127, 16, 42, 113, -119, -54, -45, -128, 26, -49, 127, 127, 127, 81, 26, 49, -32, -128, -128, 98, -127, 117, 127, -128, 127, -108, -128, 127, -128, 0, 57, 113, -93, -92, 127, -36, 127, 127, 27, -18, -47, -52, 127, 127, 127, 127, 36, -128, -79, -63, 116, 127, 127, 66, 127, 95, -128, -128, -128, -42, -88, 68, 127, 127, 127, 127, 90, 127, 108, 127, 127, 11, -10, -128, -128, -128, 127, 52, 106, 127, 127, 127, 127, 95, -128, -78, -26, -10, 127, 127, -128, 127, 127, 63, -128, 66, -128, -128, 127, -65, -128, 68, 127, -86, -53, -118, 42, -128, 48, 127, 49, 127, -23, 95, 113, -128, -47, 50, -50, 95, -60, 127, 109, 74, 127, -122, -128, 43, -128, 127, -90, 75, -16, -128, 127, 127, 127, 0, 92, -128, -128, -128, -15, 97, 111, 127, -128, 18, -42, 7, 127, 88, 127, 124, 71, -18, -54, 127, 86, 127, 8, 93, -128, -85, -7, -128, 127, -128, -43, 122, 0, -118, 127, 15, -128, -75, 21, -70, -24, -128, -128, -128, -128, -128, -128, -101, 118, -5, 127, -128, 39, 127, -86, 127, -128, 127, 127, -128, -17, -128, 85, 55, 127, 127, 127, 127, 127, -47, -128, 78, -37, -128, 127, -128, 22, -18, 127, -128, 0, 127, -128, 90, 26, -22, 127, 127, -38, -31, -128, -128, -128, -128, -128, -128, 66, -38, -128, 127, 127, -128, 127, 127, -128, 118, 114, 127, 127, 90, 127, -128, 75, 127, -128, 106, 127, -85, 127, 127, 127, 127, 127, 121, 127, 127, -128, 10, -73, -128, -57, 127, -128, -128, -36, -75, -128, 127, -128, 112, 38, -128, 111, 11, -58, -21, 13, -128, 42, -86, -128, 127, 85, -13, 127, -128, -128, -42, -114, -128, 15, -128, -128, 48, -66, 127, 92, -45, 127, -128, 127, 127, 78, -116, -128, -27, 127, 127, 127, 97, 7, -15, 10, -128, 127, -85, -128, -122, -75, -128, -85, 127, 127, 65, 121, -58, -124, -81, 118, 127, 127, 127, -74, -128, -128, -128, 127, -128, -44, 122, -128, -24, -128, -128, -128, -96, -128, -128, 127, 42, -28, 127, -128, 21, 81, -128, 127, -128, -50, -128, -81, 93, 127, 32, 127, 76, 68, 38, 127, 57, -128, -127, -128, 6, -128, 21, 127, 127, 127, 127, 127, 127, 127, 127, 127, 48, -27, -128, -128, -128, -5, -54, 24, 88, -37, 127, -33, 47, -97, 112, -128, -13, 127, -128, 127, 79, -118, 127, 107, 127, 127, -26, -128, -128, -128, 55, -111, 5, 58, -128, -90, 73, 5, -128, -128, 24, -128, 3, 127, -128, -54, 6, -128, 93, -59, -128, -128, -128, -128, -128, -128, -128, 50, -128, -64, -31, -121, 76, 114, 66, -128, 81, 10, -124, -128, -128, -119, 127, 127, 127, 127, 75, 127, 103, 127, -109, -128, -128, -128, -128, 91, 127, 68, 127, 8, 127, 127, 127, 127, 106, -128, -128, -128, -128, 26, 44, 127, 112, 127, 127, -58, -128, -55, -128, 2, -128, 78, 71, -128, 76, -128, -128, 28, 36, -128, -45, 127, 11, 127, 127, -128, 85, 127, 85, 127, -128, -128, 31, 45, 127, -75, 107, -128, -55, -34, 37, -28, 127, -16, 13, 127, 49, 127, 0, -128, -128, -96, 69, -100, 127, 38, 127, 127, -128, 127, -128, -128, 127, 127, 127, 113, 85, 127, 108, 64, -128, 127, 42, -24, 127, -128, 127, 50, -117, -128, -128, -128, -37, 127, 49, 127, 127, -128, 88, -128, -128, -123, 47, 127, 127, 127, 109, -128, 127, -128, 127, 127, -128, 127, -128, -106, 127, -128, 127, 127, 116, -32, 48, 127, 127, 127, 88, -100, -68, 95, -28, 127, 127, -102, 127, -88, -128, 88, -15, -17, 127, -114, 68, 127, -98, 127, 127, -1, 127, -128, -70, 127, 60, 127, -102, -128, -128, 127, 17, 79, -128, -128, -22, -76, 127, 85, 68, -52, -128, 127, -128, 127, 127, -128, 127, 100, 127, 127, 0, 74, -128, 119, 127, 54, 127, 127, 95, -87, -128, -128, -128, 53, 73, 36, -15, -8, -128, 57, 127, -128, 80, 127, -26, 50, 127, -128, 127, -128, 101, -91, 16, -86, -22, -128, -128, 102, -91, -128, -32, -123, 27, -97, 109, 8, 50, 6, 39, 127, -21, 127, 10, 33, -128, 127, -128, 66, 33, -128, 0, 127, 127, 127, 102, -18, -38, -128, -128, -128, 86, 28, 7, -16, 36, -128, 127, -128, -114, 70, 18, 127, 127, 127, 127, -13, 27, -49, -53, 103, 127, 127, 127, -6, 127, 0, 103, 127, 127, -43, 127, -128, 10, 54, -128, -59, 57, -127, 58, -128, -128, 127, -88, -128, -38, -128, 68, 127, 127, 66, -34, 127, -128, 118, -128, -128, 127, -128, 127, -79, -118, -128, 1, -101, -128, 111, 10, -17, -128, 42, -128, 50, -116, 70, 127, -128, 127, -15, -121, 58, -128, 0, -114, -128, 42, -128, 127, 127, 127, 73, -106, -128, -128, -128, 127, -128, 127, 127, -128, 127, -128, -128, 127, -32, -128, 127, -128, -128, -128, 27, -128, 73, 75, 127, 127, -15, -128, 75, -128, -128, -27, -128, 127, -66, 127, 55, -128, 127, -128, 45, 127, -128, 127, -127, 0, -78, 16, 127, -44, 122, -128, -116, 127, 127, 127, 127, -128, -111, -128, -128, 127, -80, 17, 127, -128, 127, 127, -48, 102, -128, -128, 69, -17, 78, 8, -128, 127, 97, 127, 127, -128, 57, 16, -44, -24, 13, -128, -128, -43, -18, 127, -34, 127, 76, 127, 127, -128, -128, -78, -59, 127, 127, -52, 127, 127, -128, 127, -128, -117, 127, -128, 127, -116, 79, -85, -73, 11, 111, 91, 127, 127, -128, 127, -128, -128, 127, -8, 10, -128, -128, -2, 28, 127, 127, 127, 127, 106, -128, 127, -128, -128, -63, 44, 42, 127, -29, 127, 127, -128, 48, -128, -28, 127, 127, -23, 127, -71, -128, 80, -128, -86, 127, 29, 127, 127, 127, 127, 127, 111, 54, 11, -127, -128, -128, -128, 127, -128, 127, 127, -128, -128, 48, -128, 48, 127, 127, 127, 127, -128, 127, -107, -128, -128, -128, -124, -128, -128, -128, 127, 54, 127, 127, 31, -128, 26, -128, 2, -70, -58, 127, -5, 127, -128, 96, -108, -128, 127, -128, -128, 127, -128, -128, -128, -128, -128, 59, -128, -18, 127, -87, 80, -33, -128, -128, -128, -22, -98, -128, -68, -128, 50, 127, -112, 3, 28, 127, 127, 127, 55, 28, 127, 57, 100, -128, -128, -86, -128, 88, 127, 127, 50, 127, 127, -10, -90, 127, -26, -128, -123, -121, -128, -128, -13, -68, -128, 50, 52, 87, 127, 127, 8, 127, 127, 127, 127, -45, -128, -128, -128, -128, 127, 127, 33, 127, 85, 127, 127, -95, 36, -18, 107, -60, 42, -98, 29, -109, 127, -128, 1, 127, -128, 127, -11, -128, 127, -128, 127, 26, -128, -128, -75, 127, -48, 127, 111, -128, 127, -128, 127, -128, 29, -44, -119, 127, -128, 106, 98, -128, -128, -128, 2, 10, 127, 127, 2, -128, -36, -128, 121, -128, 50, 127, -128, 127, -101, 127, 127, 127, 49, 124, 68, -128, 127, 127, 29, -53, 76, -128, -128, 127, 127, 0, 127, 3, -128, -21, 0, 112, 127, 127, 127, 127, -121, -128, -52, 81, 64, 127, 127, 57, 127, -23, -128, -128, -128, 76, 112, 127, 127, 127, -27, -128, -128, 38, -128, 127, -60, -5, 66, -93, 127, -128, 127, -128, 80, 127, -23, 50, -128, -28, 127, 127, -93, -128, -128, 123, 127, -3, 127, 76, 127, 127, 127, 127, -50, 127, 127, 127, -119, 87, -128, 88, 127, -128, -58, 119, -11, -70, -128, -128, 127, 127, 0, 127, -75, -107, -128, -128, -128, -128, 15, 43, -128, 127, 86, -128, 65, -128, -10, -27, -69, 127, -33, 127, -128, 127, 95, -128, 127, -128, -11, 127, -128, -128, 127, -128, 127, 127, -128, -13, 127, -128, 127, 127, -128, 69, 31, 127, -124, 127, 64, -128, 21, -60, 58, -128, -16, 127, -128, 6, 127, -128, 64, 127, 127, 127, 127, 127, -128, 127, -128, 43, -55, -96, -18, 17, -2, 31, 127, 116, 127, 49, 70, 127, 123, 127, -109, 8, -128, -128, 127, -128, 116, -17, -128, -124, -128, 79, 127, -86, 127, -128, -128, -128, -128, 127, 127, 127, 127, 127, -128, -128, -95, 88, 127, 127, 7, 65, 0, -112, 21, -128, -80, 0, 127, 127, 127, 96, -128, -47, -122, -81, 66, -63, 127, 38, -128, -128, -128, -58, -128, 127, -128, -128, 22, -90, 44, 101, 127, 127, -39, 117, -128, -128, -23, -128, 70, 38, -128, -128, -16, -74, 90, 127, 127, 108, -128, -42, -128, -128, 127, -71, 127, -73, -128, -70, 127, 118, 127, 95, -128, 38, -128, -128, -60, -128, -128, 88, -37, -128, 127, -128, 127, 127, -85, 88, -8, 127, 127, 127, 127, -108, -107, -8, 127, 127, 127, -128, -128, 8, 127, 127, 18, -128, -128, 47, 127, 127, -128, -26, -128, 127, 127, 127, -36, 127, -10, -128, 91, -10, -128, 127, -128, 119, 127, -128, 127, -86, -128, -37, -128, -128, -128, -112, -128, 58, 127, -58, -128, -1, -45, -70, -2, 15, 5, -10, 127, 64, 127, 127, 47, -128, -128, 58, -128, 23, 127, -24, 124, 127, 103, 101, 127, 127, -98, -79, -128, -128, -87, -128, -95, 127, 1, 87, 127, -48, -33, 23, 127, 11, 127, 127, 64, 127, -122, -128, -128, 48, -128, -27, 1, -128, 127, 127, -128, 127, -128, -128, -128, -128, -128, 127, 55, 127, 127, -70, 42, -128, -128, 127, -128, 127, 127, -128, 127, 127, 17, -43, 112, -128, 73, 127, 2, 127, 66, 127, -48, 49, 127, 127, 117, -128, -59, -128, -128, 127, -128, 127, 127, 6, -45, -60, -128, 27, -12, 127, 127, -75, 3, 108, -128, 38, 127, 127, 127, 86, 1, -36, 63, -128, 12, 127, 75, 103, -128, -128, -128, 127, -22, 70, 127, -12, 127, -128, 127, -38, -128, 127, -128, -117, -98, -128, -128, 127, -44, 127, 127, 127, -102, 117, -106, -128, -64, -128, -128, -128, 44, 107, 107, 66, 127, 127, 127, 127, 127, 60, -128, 47, -128, 38, -108, 127, -97, -128, 36, -128, -48, -128, -128, 63, 113, -128, 59, 27, 45, 127, -128, -128, 127, -17, 127, -95, 16, -18, 27, 127, 97, -128, 127, -128, -37, 127, -128, 127, 123, 127, 127, 127, 17, 127, -128, 52, -39, -7, 52, 69, 127, 127, 127, 107, -76, -128, -128, -81, -65, -114, -128, -128, -128, -108, -85, -57, -63, 127, -100, 111, 127, 48, -91, -124, -128, -128, -128, 33, -76, 127, 27, -128, -128, -128, -128, 127, -85, 118, -24, -90, -128, -128, -128, -108, 17, 60, -29, -121, -128, -128, 53, 113, -128, 121, -128, -79, -128, -107, 127, -69, 127, 127, 127, 78, 15, 90, 127, 127, 127, 127, -119, -100, -128, -128, 50, -128, 127, 12, -128, -45, -128, 127, -71, 127, -38, -128, -23, -128, 127, -114, -128, 16, -128, 127, -101, 98, 127, 71, 127, -22, -128, -53, 76, 127, 127, -102, -86, 127, -29, 127, 127, -128, -128, 59, -128, -128, -128, -24, -128, -88, 71, -114, -128, -68, 127, 47, -53, 127, -128, 127, 90, 15, 0, -128, -128, -128, 13, 127, 127, -128, 33, 127, -108, 127, 127, -66, 50, 127, -75, 97, 127, 127, -128, 24, 127, -28, 127, -128, -12, -128, -128, 53, -92, -122, 127, 111, -106, 127, -128, -113, 127, 100, -58, 127, 127, -48, 127, 127, 127, 37, -102, -128, -128, -88, 127, 127, 127, 92, -128, -128, -128, -128, 127, 117, 95, 127, -95, 45, 127, 117, -42, 127, -128, -87, -128, 48, -75, -8, 127, 127, 127, -128, 127, -128, -108, 23, -57, 127, 112, -60, 127, -128, -79, 95, 87, 127, 127, 127, 127, 127, -128, 127, -128, 22, 127, -128, -86, -128, -128, -128, -128, -128, -128, 117, 81, 127, 127, 109, 127, 127, -65, 127, -128, 10, 13, 1, 127, -3, -128, -128, -128, 96, -113, -39, -24, 45, 127, 127, -49, -128, -128, -128, -128, 22, 127, 127, 23, -128, -128, 21, -128, -44, 98, -128, -119, -85, -128, -128, -50, -79, -87, -128, -128, -101, -28, -63, -69, 10, 127, 127, -24, -11, -128, -128, 127, 32, 127, 127, 127, 52, -128, -128, -123, 52, -38, 127, 37, 57, 127, -128, 127, 38, 127, 127, 49, -27, -128, -128, -128, -128, -63, -73, 127, 127, 127, -128, -128, 127, -128, -128, 127, -128, -128, 103, -49, -128, -128, -2, 117, 88, 44, -128, -128, -128, -76, -128, 127, -18, -128, -55, -113, -75, -123, 1, -103, -22, 27, 114, 127, 6, 127, 127, -118, 127, 91, 127, 127, 127, -128, -128, 24, 76, 127, 68, -128, -128, -128, -128, -128, -116, -49, -11, -128, -128, 26, -128, 127, -27, 127, 127, -128, -63, -128, -128, -128, -73, 127, 86, 127, -128, -123, 127, -128, 127, 127, -128, -128, -55, 80, -128, 127, 47, -128, -95, -128, 107, 127, -76, 127, -29, 22, 127, 127, 127, 127, 113, 127, -71, 127, 127, -128, 44, -81, -26, 127, 127, 88, -128, 76, -128, -128, -64, -86, -128, -27, 127, -128, 127, 10, -42, 127, 71, 58, -128, -128, 127, -128, 127, 127, -128, 0, -128, -27, -69, 55, 127, 87, 127, 127, 127, 33, 127, -128, 127, -22, 127, 58, -128, -3, -1, 74, -8, 127, 127, -64, 127, -12, -128, -128, -128, -128, 127, -128, 127, 37, 23, 127, -68, 127, 127, -69, -128, 112, -128, 71, 78, 127, -11, 127, 29, -128, -81, -128, 127, -100, 127, 127, -87, -111, -128, 23, 127, 27, 127, -90, 127, 100, 127, -78, 52, 15, -128, 127, -128, -59, -57, -128, 74, -80, 117, 127, -128, 127, -111, -128, 85, 127, -88, 127, 127, 123, -33, -26, -128, -128, 79, 127, 127, 81, 127, -21, -128, -128, -98, 23, -128, 127, -128, -88, 12, 7, 127, 127, 127, -34, 127, -78, 63, 18, -128, 98, 93, -55, 15, -11, 37, -119, -6, -128, -128, -128, 0, -128, 127, 36, -128, -128, -128, -128, 127, -22, 118, 127, 127, 127, 127, 2, -128, -39, -128, -108, -128, -37, -128, 111, 119, 97, 127, 73, -64, 7, -128, -54, -23, 31, 127, 23, -76, -128, -128, 85, -128, 127, -98, -128, 117, 127, -128, 100, 127, 17, 1, 92, -31, 127, -97, 34, 114, 101, 127, 127, 80, 60, -128, -128, -114, 103, -128, 127, 127, -38, 127, 127, -128, 113, 127, -15, 127, -28, -128, 127, -128, 107, 127, -3, 7, -79, -1, 127, 127, -128, -27, -128, 8, -128, 127, 12, 127, 86, -79, 127, 63, -128, 50, 22, -34, 127, -128, -64, 127, -128, 127, 27, -128, 127, -2, 127, 43, 127, 113, -128, 54, -80, 123, 127, 127, 127, 127, -128, -128, 114, -128, 118, 127, -128, 53, 2, -33, 127, 127, 36, 127, -8, -128, 127, -108, -34, -128, 109, -128, 127, 127, -128, 127, -128, 96, 28, -128, 127, -128, -128, -128, 54, -38, 127, -17, -128, -128, -128, 47, -128, -128, 127, -128, 127, 127, 55, 43, -128, -128, -128, -128, 80, -78, 127, -128, 91, -128, -128, 127, 127, -2, 96, -64, -70, 102, 65, 55, 127, -128, 127, -128, -102, 55, -128, 60, 127, 127, 127, -70, 127, -49, -128, 108, 71, 127, 93, 5, -79, -128, 127, 39, -87, -86, -128, 70, 127, 127, 127, 93, 127, 90, -128, -108, 54, 127, 127, -26, 85, 23, -128, -128, 69, -128, 70, -111, -128, 127, 127, 27, 127, -71, 58, 127, -128, 39, 127, -128, 21, 127, 127, 127, 3, -128, -128, -128, 37, 127, 127, 75, 37, -81, -128, 98, 127, -118, 127, -71, -113, 63, 71, 127, 127, 127, -114, 66, 8, 6, 127, 127, 109, 53, -128, -128, -79, -128, -87, -128, 127, -128, 127, 100, -10, -32, -128, -128, -5, -111, -128, -128, 113, -50, 42, -128, -128, 48, 127, 127, 127, -128, -128, 127, 43, 108, 127, -128, 127, 127, -128, 127, -128, -36, 127, 63, 127, 127, 107, 87, 127, -116, 127, 127, 127, 127, 47, 127, 6, 127, -128, -128, -29, 88, 127, 7, -128, -128, -128, 28, 127, -70, -128, -128, -128, 10, 27, 127, 127, -128, -128, -2, -85, -124, -47, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 127, -117, -128, 60, -128, -64, 127, -31, 15, 23, -128, 127, 127, -22, -128, -128, -128, -66, 11, 96, -128, -128, 111, 86, 127, 127, 11, 127, -80, 1, 127, -29, 71, 118, 88, 127, -93, 127, -128, -85, -128, -128, 127, -128, -3, 127, 127, 127, -128, -79, -128, 127, -64, -52, 127, -47, 127, -128, -80, -73, -128, 90, -128, -128, 64, -128, -13, 106, 7, 127, 73, -106, 127, 33, 0, 127, -128, -29, 127, 101, -91, 127, -128, -128, 44, 33, 127, -53, -128, -53, -128, 127, 15, 127, 127, 109, 127, 127, 127, 127, 127, -128, -128, 22, -52, 127, 127, -57, -10, -102, -128, -128, 127, -128, 22, 68, -128, 127, -68, 127, 127, -36, 127, 127, -128, 127, -109, -16, -128, 127, 93, -128, 12, -128, -128, 127, 127, 127, 28, 55, -44, -128, -128, -128, -128, -114, 59, 127, 127, -47, 127, -128, -128, 127, -10, -58, -95, -128, 127, -47, -13, 127, 49, -12, 127, 92, -11, 127, 127, 127, -80, 13, -58, -55, 127, -128, -128, -49, 18, 127, -119, 127, 127, -128, 127, -87, -11, -128, -128, -75, 64, 75, 127, 127, 127, 29, 127, -128, 127, -47, -6, 17, -107, -128, 127, -68, 17, -45, -75, 127, -128, 69, 127, 127, 127, 85, 50, -86, 127, 127, 68, -74, 15, -100, 102, 47, -97, -128, -128, -128, -128, 103, 49, 127, 127, 127, 127, 127, -27, 108, -49, -34, 127, 86, 127, 127, -6, -128, 127, -128, -44, 60, -128, -29, -44, 49, 127, 86, -128, -128, -70, 127, -44, 127, 66, 127, -113, 63, 127, -128, 127, 23, -128, 127, -128, 127, -128, 47, 127, 50, -6, -128, -128, -128, 91, 13, -76, 28, -1, -55, -107, -128, -128, -128, 59, -122, -65, 127, 23, 127, 127, -5, 127, -68, -39, -128, -128, 78, -128, -106, 127, -128, 66, 127, -73, 127, 79, -33, 127, 106, 127, 127, 50, -128, -128, 112, -128, -1, 26, -128, -128, -64, -128, -63, 117, -26, 127, 50, 127, -128, -16, -128, 127, 127, -128, -128, 27, -101, -128, 1, -128, -75, 85, -128, -70, -128, -128, -112, 42, 127, 127, 127, -23, 87, 127, -102, 127, 127, 127, 127, 127, 45, 127, -58, 127, 26, -121, 98, -75, 127, -59, -116, -128, -128, -128, -37, -11, -90, -128, 127, -128, 127, 23, -128, -128, -128, -128, -21, -128, 55, -22, 127, 127, 59, -128, -128, -106, 127, 127, 127, 123, -81, -128, -128, 5, 74, 101, 127, 91, 39, 127, -1, -128, -128, -128, -128, -128, -128, -128, -15, -128, -64, -128, 92, 8, -128, -42, -128, 78, 127, 36, -107, -128, -128, -128, -128, -128, -128, -128, -128, 92, 127, 50, 127, -108, 42, 127, -50, 127, -15, -128, 3, -91, -90, 127, -128, -128, 127, -128, -107, 127, -128, -128, 52, -128, -128, -128, -123, 127, 127, 127, -128, 10, -128, -103, 127, 127, 127, 127, 127, 127, -44, 127, 7, -128, 107, -128, 127, 127, 127, 127, -63, -128, -128, -128, -128, 0, -108, -114, -128, -128, -128, -128, 127, 7, 34, 127, -128, 127, 71, 127, 127, 127, 108, 127, 127, 127, 127, 127, 63, 127, -80, -128, 95, -128, -18, 127, 127, 7, 127, 127, 65, 29, -128, 63, -91, 64, 33, -128, -128, -109, 64, 127, 114, 127, -3, 127, 127, 43, 65, -128, -128, -128, 117, -80, -118, 127, -128, -128, -128, -128, -128, -128, -128, -128, 37, 127, 33, -121, -21, -106, 127, 127, 127, 127, -128, 55, -128, 88, -100, -109, 127, -44, 127, -66, 85, 127, 127, 54, -128, -128, 127, 91, 127, -128, -71, 127, -68, 127, 127, -13, 16, -128, -128, -128, -39, -128, -28, 127, -128, 97, 127, -128, -128, 78, -128, -119, 85, 127, 90, -128, -39, -128, -128, -128, 86, -128, 127, 127, -128, 127, 27, -128, 102, 127, 2, 127, 32, 127, -6, 127, 91, -60, 127, -128, 98, -128, -79, -48, -128, 127, -124, -98, -128, 116, -128, 39, -123, -128, 127, 95, 127, 8, -128, -128, -122, 121, 127, 127, 127, 22, 42, 127, -128, -121, -118, -128, -21, 127, 24, 34, 127, 24, 34, 54, -128, -128, -128, 32, 26, 7, 96, -128, -128, -117, -128, 109, 64, 127, 127, 127, 127, 127, 2, 81, -113, -128, -122, -101, -127, 127, -101, 127, 127, -24, 11, -128, -128, -128, -128, 92, 127, 43, -87, -102, 21, 28, 36, 127, -128, -93, 127, -5, 10, -123, -128, 127, 127, -7, -33, -128, -128, -128, 1, 96, -123, -128, -128, -55, -52, -16, 39, -98, -128, -128, -128, -128, -7, -124, -128, 127, -128, 13, 127, 75, 5, -36, -128, -128, -52, -128, 127, 127, -128, 127, -114, 127, 96, -66, -128, -128, -128, 127, 16, 127, -128, -71, -121, -128, -7, -128, 127, -87, 88, 127, -21, 12, 71, -49, -90, 22, 18, 58, 127, 127, 127, 117, -128, -59, -128, -92, -128, -128, 15, -97, -128, -128, -128, -1, -128, -43, 127, 127, 127, 127, -79, -128, -128, -128, -128, -128, -128, 121, -128, 127, 127, -128, -128, -69, 36, 117, 127, 127, 93, 64, 3, -128, -128, 127, -128, 88, -108, -128, 90, -11, 127, 119, 127, 127, 127, 127, 127, 127, 127, 45, -111, -80, 22, 26, -122, -86, 24, 7, -88, -128, -128, -23, 59, 127, -108, -114, 75, 124, 59, 127, 127, 31, 127, -54, -128, 127, -48, 69, -33, -128, 96, -128, 121, 127, -10, -128, -113, -128, 0, -43, -128, 53, 47, 127, -10, 127, -128, -23, 127, -32, -79, 5, -128, -128, -128, -128, -128, 92, 127, 127, 7, 127, 24, -122, 47, -37, -15, 127, 50, 127, 127, 127, -32, 69, -128, -128, 127, -13, 53, -128, -6, -122, 5, -128, -128, -128, 127, 43, 127, 127, -128, 127, -90, -128, -70, -128, -117, -128, -55, -128, -11, 127, 127, 127, 127, 66, -128, -128, -128, -128, 26, 127, 127, -128, 127, -128, -128, 127, -37, 127, 27, -12, -128, -128, -128, 127, 39, -128, 73, -91, -55, -87, -128, 58, 91, -54, 127, -6, -128, -128, -68, -33, 127, 127, 79, 127, 127, -128, -118, -54, 127, 109, -97, 80, -128, -128, 47, -128, -81, -128, -3, -118, -128, -128, -128, 80, 127, 127, 127, 90, -64, -128, 127, -128, 113, -10, -128, 127, -128, 18, 127, -128, -33, 127, 127, 127, 127, -128, 70, -128, -39, 33, -21, -128, -128, -6, -128, -128, 127, -13, 127, -128, 45, -128, -128, 127, 33, -128, 114, 127, -128, 127, 16, -128, -106, -128, 122, -128, -128, -49, -6, 127, 127, 127, 23, -6, -128, -128, -128, -128, 127, 75, -43, -128, -128, -31, -7, 127, 127, 127, 127, -54, 53, 127, 124, -124, 127, -91, -128, 127, -128, -128, -103, -128, 13, 27, 127, 127, 57, 123, -128, 57, -128, 26, 127, -128, 18, -32, 127, 127, 127, 127, -107, 127, 123, -128, 127, -128, 127, 76, 127, 127, -81, -128, -128, 13, -128, 103, 127, -111, 127, 127, 127, 127, 127, 127, -128, -128, -34, -128, -128, -128, -54, -15, -57, -128, -128, -128, -29, 127, -86, 127, -79, 127, -95, 88, 127, -128, -128, 57, -128, -38, 127, -128, 121, -122, -128, -128, -128, 116, -128, 127, -101, -34, 79, 3, 79, 127, 127, 0, 95, 111, -5, -13, 109, 127, -8, -128, -128, -128, 12, 87, 127, 127, -71, 127, -111, -128, 24, -128, -23, -128, -48, 8, 33, 127, -128, -128, -124, 96, 127, 39, 127, -128, -128, 52, -81, -128, 75, -121, 63, 113, -118, -34, -109, -22, 127, 57, -128, 109, -128, 127, -8, 92, -92, -108, -123, -128, -128, 127, -7, 124, 31, -128, -128, 0, 127, 127, 58, 127, -23, 69, -2, -17, -128, 101, 11, -128, 5, -128, -96, -128, -128, 127, -128, 12, 127, -6, -23, 127, -3, 127, 10, 16, -68, 78, 127, -103, 38, 92, 127, 127, 127, -54, -60, -69, -128, -49, -128, -1, -31, 15, 127, 37, 29, 127, 127, -52, 127, 73, 114, 93, -75, -128, -128, -16, 127, 127, -64, 127, -128, -39, 48, 117, 127, 127, 127, 127, -65, 111, 127, -81, 127, 65, -128, 127, -128, 93, 13, -23, 127, 127, 53, 127, -8, -53, -128, -114, -128, -128, -128, -128, -73, 127, 54, 127, -22, -91, -128, -58, -128, -1, 127, -10, -128, -7, -128, 100, -128, 102, 127, -128, 78, -128, -128, -128, -128, 127, -128, 59, 127, -128, -128, -128, -90, -13, 127, 86, -47, -128, -95, 127, 127, -128, -48, -113, 112, 127, 127, 127, 91, 127, 109, 127, 127, 127, -118, -128, -81, -128, 127, 0, 127, 55, -108, -128, -128, -128, -128, -12, -128, 107, 127, -112, -128, -128, -128, 127, 127, 127, 127, 127, -53, -128, 50, -128, -60, 15, 127, -95, -124, 95, 127, -76, 75, 127, -128, 127, 127, 27, 127, -24, 127, -22, -128, -68, 108, -52, 68, 127, -6, 127, -38, -128, -43, 127, 47, 127, -128, -128, 50, 127, 127, 8, 95, -128, -128, 127, -78, 127, 127, -54, 91, -50, -127, -5, -128, 127, -128, 127, -128, -119, 37, 71, 127, 127, 38, 127, 57, -128, -128, -128, 80, 45, 107, 64, -128, -117, -128, 127, -102, 127, 100, -122, -128, -128, -128, -102, -13, 127, 127, 127, 11, 127, -65, -75, 127, -128, 127, 127, -128, -119, -128, -37, -80, -76, 127, 127, -128, 127, 13, -128, 127, -128, -128, -68, -128, 127, -22, 116, 127, 2, 127, 127, -128, 102, -68, -128, 127, -128, 21, -128, -103, 127, 127, 127, 127, 127, -128, -128, -73, -37, -6, 127, -54, 127, 127, 127, 97, 39, -50, -128, -122, -23, 127, 127, 127, 127, -116, 127, 113, 45, 88, -80, 13, 127, 127, 127, 78, 127, -128, 0, 127, 106, 127, 127, -128, -38, -44, -128, -128, 127, 34, -116, 127, -128, 76, 97, -128, -128, -128, -128, -76, 37, 127, 127, 119, 116, -128, -128, 16, -128, 96, -128, 47, -27, -96, -59, -87, -128, -97, 127, 91, 127, 16, -128, 68, 43, 127, 81, -128, 88, 127, 0, 42, -71, -128, -128, 31, -127, 119, 86, -112, 127, -3, -42, 127, -128, 106, -128, -128, 127, -55, 102, 42, -27, -128, 8, -128, 53, 127, 64, 127, 127, 60, 86, 122, -31, -128, -128, 55, -128, 127, 23, 2, -101, -128, -36, -128, -27, -26, -103, 27, 127, -128, 73, 127, 114, 127, 127, 127, 127, 127, 127, 127, 58, 127, 127, 127, -39, -128, -128, 127, -128, 127, 127, -118, -128, -128, -128, -128, -128, -128, -128, -128, -79, 11, -101, -76, -102, -128, -128, -16, 127, -128, 127, 127, -57, 127, -48, -2, 127, -128, -29, -128, -128, 55, 127, 127, 90, -1, -45, -128, -23, 60, -128, 81, -128, -50, 127, 68, 127, 127, -74, 127, -81, 66, 127, 127, 69, 127, -128, -128, 101, -121, -18, 127, -128, 122, -98, -38, 127, 127, 127, 127, -37, 127, -128, -39, 127, 127, 127, 127, 127, 127, -21, 33, 28, 127, 127, -91, 10, 50, -58, -128, -101, -106, 85, 127, 96, 127, 76, 127, 32, -69, -128, -128, -128, -128, -128, -54, -128, -57, -128, -128, 57, -128, 2, -128, 34, 44, 15, 10, -128, -128, -85, -128, 87, 127, -73, 127, 28, -33, 127, 42, -90, 63, -96, -128, -33, -128, -79, -128, 71, 127, 127, 49, -128, -128, -128, -128, -128, 70, 37, 127, 85, -90, -128, -128, 37, -102, -128, 88, 2, -12, 127, -53, -16, 127, -107, 127, 127, -73, 65, -128, -128, -13, 10, 127, 127, 12, -128, -128, -128, -128, 127, -128, 127, -128, -107, 127, -90, 127, 70, 127, 127, -128, 127, -128, -8, 127, 127, 127, 127, 127, -128, -128, -128, 74, 127, 127, 127, 17, 127, -128, -128, 65, 127, 127, 32, -128, -52, -128, 34, 127, -128, 29, -8, 23, -128, 127, -103, -43, -11, -128, -128, -128, -128, -34, 68, 127, 127, 127, -15, -93, 127, 108, 127, -68, 15, -128, -128, -52, 90, 127, 127, 127, 127, -128, 127, -64, -48, 127, -128, -128, -128, -128, -68, -128, 65, 127, -23, 127, 49, -106, -128, -128, -128, 93, 127, 127, -10, -128, -128, -33, 127, 127, 127, 127, 75, 127, -92, -128, -47, 117, 127, 38, -85, -128, 58, 87, 68, 59, 127, -86, -128, -17, -24, -128, 127, -101, -15, 127, 1, 127, -24, 2, 38, -109, 36, -128, -128, 7, -128, -47, -17, 3, 127, -128, -128, -23, 45, 127, 127, 127, 127, 127, 127, 127, 127, 50, -128, -128, 53, -128, 127, 117, 69, -76, -107, -128, -128, -128, -128, 116, 127, 96, 127, -111, 97, 114, 127, 127, 88, 127, -128, 98, -128, -47, 127, -128, -45, 71, -128, 6, -26, -128, -128, -128, -128, 60, -81, -128, -24, -128, -128, 59, 24, 42, 127, 16, 127, 127, 127, 127, 98, 127, -128, 86, 15, -128, -128, -39, -128, 107, 127, -122, 81, -128, 80, -106, 28, 8, -70, 127, -102, 127, -49, -55, -128, -73, -128, -128, -128, -128, 74, -81, -128, 122, -128, 127, 95, -6, 0, 98, 127, 2, 127, -128, -36, 127, -45, -101, -128, 65, -128, 127, 107, 114, -107, 10, -128, -90, 6, 127, 116, -128, -96, -68, -116, 127, 29, -128, 127, -128, -116, 127, 117, 127, -33, 98, -128, 5, 127, -103, 28, -128, -128, -49, -17, -107, 92, -11, 127, -75, 127, -95, -128, 127, -128, 127, 95, -128, -86, -128, 127, 127, 17, 127, 127, -18, 1, -128, -128, -128, -127, 127, -78, -128, -128, -128, 101, -128, 74, 127, -10, 127, 127, -74, 42, -128, -128, -7, 85, 127, 127, 118, 127, 127, -93, 54, 69, -119, -128, 79, -128, -128, 3, -128, -128, 85, -128, -128, -128, -128, 10, -122, -128, 127, -128, -85, -128, -128, -24, -128, 29, -122, -128, -93, -128, -128, -29, -48, -123, 127, 65, 127, -39, 127, -21, -128, 127, -128, 127, -96, 127, -45, -74, 33, -16, 127, -112, -32, -48, 58, 127, -79, -76, -128, -128, -66, 112, -128, 127, -49, -128, -106, -128, -8, -128, 127, 63, 18, -87, -128, -128, 127, -86, 127, 127, -44, 127, -128, -128, 127, -6, -50, 6, 43, 127, 127, 127, -128, 114, -128, -43, 92, -128, 97, 0, 127, 127, 127, 12, 127, -43, -128, -108, -128, -63, 111, 79, -114, 127, -66, -78, 71, -42, -128, 92, 127, 81, 127, 127, -100, 127, 127, -16, 22, -112, -128, 16, 1, -128, 45, -128, -16, -128, -106, 81, 127, 127, 127, 127, -128, 127, -128, -66, 0, -128, -128, -128, -36, 17, -122, 127, -128, -69, -121, -128, 127, 93, 127, 113, 11, 127, -128, 127, -128, -128, 127, -128, 127, 127, 59, -26, -128, -44, -26, -32, -128, -128, -70, -128, 81, 127, 24, -75, 95, 127, 98, 127, -24, -128, -128, -8, 60, 28, 127, 127, 127, 127, -128, -15, -128, 44, 28, -128, -128, -128, 24, -128, 16, -128, -128, -128, 97, 127, 127, 127, 127, 2, -128, -128, -128, -128, 127, 80, 127, 85, -128, -49, -128, -128, -128, -128, -11, -74, -23, -128, -128, -95, -128, -42, 107, -128, -45, 73, -128, 111, 127, -128, 127, -31, -128, 80, -107, 127, 127, 127, 127, 127, 127, 57, -102, -48, 127, -96, 127, -128, 127, -32, 107, 127, -128, -3, -128, 13, 127, 127, 127, 127, -5, 76, 53, 91, 127, 127, 127, 60, -128, 127, 53, 127, 127, -128, -128, 58, 33, 127, -123, -128, -128, -128, -85, 45, 45, 127, 127, -76, -128, -128, 79, -16, 127, 97, 43, -128, 109, -21, 45, -128, 85, -128, -128, 127, -6, -103, -128, -107, 127, 49, 127, 102, 24, -93, -128, -37, -38, 127, 3, 127, 127, -128, 103, 1, 3, 15, -128, -74, -128, -128, -128, -112, -128, 91, 95, 127, 31, 45, 127, 127, 127, 95, -128, -12, 127, -101, 127, 127, -114, 0, 127, 127, 95, 127, -33, -128, 90, 5, -17, 127, 127, 127, 127, 127, -128, 127, -112, -92, 50, -128, -128, -128, -128, 63, 127, 21, -71, 63, 76, 118, 127, 108, -75, -128, 26, -28, -128, 127, -128, -74, 127, 45, 31, 127, -128, 58, 127, -106, 117, -128, 12, -128, 127, 127, 127, 127, 68, -128, 47, -60, -93, -128, 2, -128, -128, 127, 0, -6, 127, -17, -103, -128, -128, -26, -12, 127, -60, -13, 127, 127, 127, -50, 127, -128, -48, -49, 108, 26, 36, 127, 1, 71, 127, -31, 81, 127, 28, 58, -38, -128, -128, -128, -128, 127, 44, -128, 112, -32, -128, 127, 127, -128, 127, 3, -128, 33, -128, -128, -128, 59, 127, 6, 127, -128, -128, 123, -128, 0, -128, -128, 70, 127, -74, 17, -128, -36, 127, 101, 36, -86, -128, -128, 29, 49, -128, -113, 127, -128, -1, 52, 92, -70, -128, -57, -22, 127, 127, 27, 127, -128, -128, -128, -128, 121, 107, 127, -128, -76, -112, -21, 85, 127, -66, 127, 52, -23, 127, -55, 53, -100, -128, -128, -34, -15, 127, -128, -128, 127, 108, 34, 127, -128, 86, -128, -76, 127, -128, 127, -12, -70, 127, -128, 127, -59, 127, 86, -128, -128, -128, 63, -128, 127, 36, -128, 127, 38, 37, 127, -93, 127, 127, -128, 127, 112, -128, 127, -128, -69, -52, -128, -128, -128, -73, 33, -128, 127, -26, 101, -128, -122, 127, 76, 95, 127, -128, 17, -119, -128, -128, -128, 127, -128, 127, -74, -128, 127, -73, 34, 127, 103, 123, 127, 127, -17, 127, 0, -128, 79, 5, -128, 127, -111, -90, 127, 74, 127, 127, -128, 127, -47, -128, 127, -10, -38, -128, 50, -128, -128, 127, 34, 127, 127, -128, -128, 100, -128, -79, -24, 127, 5, 127, -119, 127, -128, 127, -128, -128, 127, 127, 127, 127, 127, -22, 127, -128, -45, 127, -106, -5, -73, -96, 127, 101, 8, -39, -128, -128, 127, 108, 127, -66, -128, -114, -71, 127, -48, -85, 57, 55, 1, -92, -128, -128, -33, -50, 127, 127, 127, 127, -128, -128, -128, 124, 127, 127, 127, -128, -128, -63, -29, 127, 127, -75, 44, -128, 37, 86, 127, 127, 127, 127, 127, -33, -70, 26, 127, -68, 114, -5, 127, -98, 127, -74, 118, 127, 18, -128, 123, -128, -21, 90, -95, -50, -128, -23, -22, -128, -111, 22, -16, -2, -74, -128, -128, -5, -128, -114, -114, 117, 116, 93, 127, -114, -128, -128, -128, 73, 96, -128, 111, 0, -128, -128, -116, 78, 127, 127, -88, 127, -98, -128, 127, -112, -64, 127, 113, 127, 64, -128, 93, -128, 127, -106, -28, 127, 127, 127, -45, -16, -27, 127, -34, 127, -78, -76, 127, -54, 91, -128, -128, -23, 127, -113, 127, 0, -128, -23, -128, 88, -128, 109, 127, -64, 127, 127, 127, 123, -23, -23, -128, -6, 121, 127, 127, -3, 13, 45, 127, 127, 127, 127, -128, -78, -128, -128, -128, 24, -128, -124, 127, -128, 117, -128, -44, -13, -10, 127, -128, -29, 87, -92, -7, -42, -128, -128, 5, 12, 43, 127, -128, -128, -128, 76, 80, 91, 49, -128, 127, -103, 127, -10, 127, -128, 86, 127, -128, 127, -128, -37, 59, -128, 127, -121, -128, -15, -128, -128, 16, -32, 127, 127, -31, 66, 127, -128, 127, 58, -128, 95, -101, -128, -128, -111, 127, -21, 127, 127, -128, -96, 127, -128, -65, 127, 31, 127, 127, -66, -128, -128, -47, 88, 47, 127, -11, -54, 127, 16, 127, 7, 127, 127, -102, 12, -128, -128, 103, -128, 127, -103, -128, 127, -128, 127, 127, 127, 127, 127, 127, -128, -86, 127, 59, 127, -128, -103, 0, -128, 92, 127, 127, 127, -88, 10, -128, -128, -128, -128, -10, -128, -128, -128, 23, 75, 127, 127, 127, -128, 32, -128, 44, 127, 127, 127, -127, -128, 121, 28, -69, 127, 127, 127, 127, 127, 127, -128, -112, 22, 127, 127, 127, -74, -128, 127, -79, -128, 18, -118, 127, 78, 127, 8, 58, 63, -128, 127, 7, 127, -80, 127, -81, -128, 127, -128, -128, 121, 70, -52, 78, -128, -86, -128, 75, 0, -128, -45, 32, 8, 127, -101, -128, -90, -128, 69, 127, 116, 127, 127, 127, 127, 28, 22, -88, 29, 127, 127, 127, 127, 127, 123, -128, -128, -90, 127, 70, -27, -128, -128, -128, 47, 127, 127, 127, 21, 117, 64, -76, 49, -128, -128, 18, 127, -43, 127, -128, -65, -33, -106, 127, -48, -48, -128, -128, -128, -97, 127, 88, 127, 13, 127, 127, 43, -98, -111, -128, -86, -21, -128, -128, -128, -54, 127, 127, -24, -128, -128, -128, -101, -87, 127, 23, 109, 127, 70, 58, 127, -39, -128, 28, -128, -128, -128, -128, 18, -128, -23, 127, -128, 33, -128, -128, 53, -128, 123, -24, -128, -128, -128, -55, 127, 2, -36, -23, -76, 76, -112, -128, -128, -128, -128, -128, 127, -128, 108, 127, -128, 127, -95, -128, -69, -128, 26, 127, -63, 127, 127, -128, 44, -128, -128, 127, -128, 127, -10, -98, 127, -11, 127, 127, 127, 127, 34, 127, 127, -128, 127, -97, -128, -128, -128, -128, 107, 92, -52, 127, -106, 127, -128, 127, -96, -118, 127, 127, 127, 127, -112, -49, -128, -128, -122, 127, -128, 127, 127, -128, -128, -128, 81, 6, 127, 71, 113, 127, 127, 16, -128, -128, 11, 127, 127, 13, -128, -128, -128, -128, 127, 13, 127, 127, 127, 127, 58, -128, -103, 93, 127, 127, 127, 28, 101, 127, -128, 127, -128, -86, -95, 7, -23, 57, -16, -127, 31, -128, 23, -128, -128, -26, -96, 119, -42, -128, -111, 127, -128, 127, 127, -8, -128, 24, -101, -93, -128, -128, -123, -22, 127, -87, 127, -128, -128, 53, 127, -13, 127, -34, -128, -87, -113, -128, -75, 63, 127, 127, 127, 127, 127, 127, -32, 127, -128, -128, -52, 86, 127, 8, 49, 98, 96, 16, 127, 17, -128, -52, 53, 97, 127, 127, -90, 127, 127, 127, 127, 127, 127, 127, -128, 6, -55, -21, -128, 18, -80, -128, 127, 121, 24, 127, 85, 65, -80, -128, 16, -27, 80, 59, -22, 12, -31, 127, -128, 127, -128, 127, -31, -98, 60, -11, -128, 78, -79, -128, -128, -128, -75, -128, 15, -18, 127, 127, 127, 127, -128, 127, -128, -128, 127, 98, 127, -45, 127, -128, 21, 127, 127, 127, 103, 127, 52, 127, -16, 63, 127, -128, 59, -128, -73, 36, -128, 85, -128, -1, -128, -128, 127, -58, -128, -5, -128, -128, -47, -27, 127, -11, 54, 127, -118, 127, 96, 70, 106, 127, 127, 127, 21, -128, -128, 47, 127, -22, 127, -128, 2, 1, -50, 127, 123, 127, -26, -128, -128, -128, -22, -128, 127, -128, -128, 114, 53, 127, 39, 127, 127, -128, -128, 44, -128, 87, 127, 12, 127, 127, 108, 127, 107, -17, -5, -128, -128, -123, -8, 127, 127, 127, 90, -128, 1, -108, -11, -128, -128, -128, -49, 127, 127, 127, 127, -128, -103, 63, -128, 127, 127, -28, -113, -128, -128, -106, -65, -128, 127, -57, 68, 24, 90, -128, 116, 103, -128, -48, -128, -128, -128, -55, 112, 43, 24, -128, -128, 127, 42, 38, -128, -128, -128, -10, -117, -128, 123, -36, -128, 127, -128, 36, 95, -128, -128, -128, 107, 127, 0, 127, -128, 34, 127, 127, 96, 60, 127, -87, 65, 116, 69, 127, 127, 127, 127, 47, 81, -128, 66, -128, -128, 127, -128, 127, 127, -85, 127, 92, 54, 101, 127, 127, 127, -65, 127, -128, -128, 127, -128, -128, -96, -128, -128, 127, -128, -128, 106, -128, 23, 127, 47, 127, 63, 2, -128, -76, -128, 43, -128, -27, 127, 31, 127, 127, 127, 57, 127, -88, -128, -49, -128, 123, 71, 127, 93, -76, 58, -128, -128, 34, -128, 127, 10, -128, -128, -128, -128, -128, -47, -128, -128, -128, 50, 15, 127, 78, -128, -37, 127, 22, -128, -113, -128, -128, -128, -128, 127, 127, 3, -128, -88, -128, 52, 127, -38, 45, 42, -107, 59, -8, 53, 127, 127, 28, 127, -128, -128, 106, -78, 127, 127, 127, 127, 127, 127, 39, 127, -64, -106, -128, -128, -71, -128, -128, 127, -86, 127, 3, -128, 121, -52, -13, 127, -54, -73, 85, 127, 127, -128, -81, 116, -128, 127, 127, 127, 80, 6, -128, -128, -128, -128, 127, 116, 121, -128, 52, -128, 127, 127, -58, 127, -112, -128, -63, -93, 117, 108, 127, -128, 127, 52, -128, -128, -128, -113, -128, -128, -128, -128, -28, 127, -58, 70, 127, -75, 98, 73, -128, -128, -128, 16, -128, 22, -44, -128, -128, -128, -128, -128, -109, 127, -128, -48, 26, -128, 127, 71, -65, -128, -128, 24, -128, 2, 127, -128, -21, 52, -128, 63, -32, -128, -111, -76, -128, 127, 127, 127, -102, -128, 66, 127, 127, 127, 64, -118, -50, -128, -128, -65, -128, 93, 27, -128, -13, -128, 55, 127, 127, -85, -128, -128, -128, 127, 39, 37, 10, -128, -128, -128, -128, 103, -128, 127, -128, 18, 74, -128, -66, -90, 98, -12, 127, -92, -128, -90, -128, -112, 127, 60, 45, -88, -128, -128, -128, 58, -128, -3, 7, 86, 127, 127, 127, 127, 127, -26, -128, -128, -128, -128, 109, 127, 79, 112, -5, -128, 127, -76, 127, -22, -128, 127, -128, -128, 127, 71, 127, 127, -128, 127, -128, 127, -59, 78, -18, -78, 127, 127, 6, 127, -128, -57, -17, -128, 0, 127, -29, 93, 0, 127, 26, -128, 127, 58, -102, -75, -113, -128, -27, -57, -128, -128, -113, -128, -128, 127, -111, -128, 6, -128, -33, -113, -128, 127, 50, 127, -50, 34, -128, -128, 0, -128, -128, -128, -80, -128, 127, -12, 15, 127, -128, 127, -128, 98, -87, 102, -73, 127, 127, -128, -59, -128, -128, -8, 127, 127, 127, 127, -128, -128, -128, 11, -128, -37, 10, 127, 127, 127, -53, 52, -128, -128, 127, -34, -1, -128, -128, -128, 127, 37, 127, 127, -27, 0, -90, -128, -128, 127, -76, 127, 127, -80, 127, 127, 8, 64, -128, -128, -22, 64, 100, -128, -34, -90, -128, -68, 92, -128, 58, 127, -42, 85, -128, -128, -128, 23, 127, 127, 127, -128, 98, -23, -128, 127, -128, -128, 127, -71, -128, -123, 17, -109, -24, 80, -128, 121, -128, -128, -48, -97, 127, -118, 122, 86, 109, 127, -52, -128, -128, -50, -6, -71, -18, -121, 55, 127, 127, 127, 127, 127, -128, -128, 91, -128, 38, 66, -128, -128, -128, -128, -36, 2, 127, 127, 54, 11, 38, -128, -64, -34, -65, 0, -128, 92, -128, 127, 127, -90, 127, 127, 127, -128, -113, 34, 127, -13, 127, 127, 39, 80, -128, -59, -128, -128, -128, -127, -128, -128, 116, -128, 111, 127, 90, 127, -128, -128, -128, -128, 91, -128, -128, 127, 111, -128, 127, 36, 127, 27, 127, -128, -17, -3, -128, -128, -102, -91, 117, 0, -106, -128, 27, -12, -128, 92, -128, -128, -5, -128, -128, 24, 127, 127, 127, 18, -128, 123, -57, -128, 127, 127, 127, 127, -24, 12, -113, 127, 127, 127, -128, 24, 127, -106, 38, -128, -128, 127, 127, 76, 127, -128, 96, -128, -128, 81, 101, -39, 127, -8, -58, 127, 127, 127, 47, -128, -58, 85, -128, 127, -50, -42, -128, 10, -103, 127, -37, 47, 127, -86, 127, 127, -128, 17, 90, 106, 91, -39, 127, -127, -128, 127, -128, 43, 127, 103, 127, -17, -128, -128, -128, -3, 127, -13, 127, -128, -128, 127, -128, 21, -80, 16, 127, 127, -71, 54, -128, -128, 6, -128, -90, -128, -128, -128, -128, -38, 24, -108, 106, -128, -128, -128, -128, -60, -98, -128, -114, 64, 36, -128, -59, -91, -24, 127, 95, 127, 127, -6, 127, 78, -23, 52, 127, 100, -128, 31, -10, -128, 127, -128, 45, -127, -128, 69, -128, -13, -23, -128, -107, -128, -128, -128, -128, -128, -128, -128, 100, 127, -24, 71, -102, -128, -69, -128, -128, -128, 118, -128, 127, -92, -128, -128, 71, -128, 127, 127, 127, 123, 127, 12, 12, 34, -128, 127, 66, -128, 127, 116, -128, 127, 127, -64, -128, -38, -128, -128, -29, 127, -49, 127, -69, -128, -128, 24, -128, 3, -93, -128, -128, -128, 59, 127, 127, 127, -52, -128, -49, -59, 37, -128, -128, -128, -128, 127, 127, 3, 127, -128, -128, 66, 127, 124, 121, -128, -128, 88, -128, 127, -128, 79, -7, -128, -7, -128, -121, 127, -23, 127, 127, -128, -128, 53, 127, 27, 127, -128, 37, -128, -128, 127, -128, -128, 127, -128, 6, 127, -128, 127, 127, -66, -34, -128, -128, 38, 127, -2, -128, -73, -128, 116, 127, -91, -128, -36, -128, -128, 127, -128, 127, 127, 127, 64, 127, 23, -128, -52, -128, -128, -128, -128, -128, -109, -91, 127, 127, 127, 127, 127, 127, 127, -97, 127, 127, 63, 127, -111, 127, 5, -128, -128, -12, -128, 119, -70, -128, -128, 85, 81, -57, 127, -128, -91, -128, -128, -44, 127, -27, 107, 127, -128, 68, 127, 127, 127, 55, 86, 127, 101, 127, -63, -116, 26, 34, 127, 127, 127, 127, 127, -128, 13, -128, -128, 127, -128, 127, 127, -80, -28, -74, -128, -128, -43, 106, 127, -128, -48, -118, 127, 18, -43, 127, -128, 127, 11, -128, 92, -128, -128, 75, -128, 70, 127, 5, 127, -128, 127, -29, 127, 127, -128, 22, -116, 127, -23, 127, 127, -128, 127, -128, 42, -113, -128, 127, -128, -108, 73, 127, 127, -76, 127, -128, -55, -107, -128, -43, 127, 33, 127, -42, -71, 123, 59, -11, -128, -114, -128, 86, -50, 21, 118, 127, 114, 127, -31, -128, 36, -128, -128, -128, -128, -128, -27, 127, -27, 127, 127, 127, 127, 113, 106, 127, 127, 127, 127, 127, -128, -128, 44, -65, 127, -11, -50, 127, -86, 12, -49, -128, -53, 79, 23, -93, -128, 86, -128, 65, 127, -114, -128, -128, -128, 43, 127, 127, 127, 127, 78, -3, 50, -128, 58, -128, -48, 127, -128, 127, 87, -128, -128, -128, -128, -128, -76, -128, 127, 127, -128, 1, 127, -3, 97, -128, -57, -128, 81, 127, -28, 127, 127, 127, 127, 127, -128, -128, 127, 127, -128, 127, 58, -128, 38, -128, -128, -128, -97, -128, -16, 127, 127, -109, 58, 103, 127, 127, -91, 127, -116, -128, 127, -128, 127, 127, -128, -128, -128, -5, -32, 127, -42, -128, -128, -128, -6, -128, -128, -31, -128, -16, 127, -119, -128, -15, -128, 127, 127, -128, -21, 116, 127, -10, 93, 100, 127, 127, -60, -128, -23, -108, 127, -17, 17, 127, -97, 127, 108, 32, -81, 16, -128, -70, -88, -128, -54, -65, 8, 47, 113, -128, -128, -128, 88, 22, -128, 60, 127, -80, 101, 127, -128, 127, 127, 31, 127, 127, -127, 50, 31, 127, 127, 127, 127, 127, 127, 127, 127, -128, 127, -96, -128, 127, 127, 127, 3, 127, 127, -86, 5, -71, -128, -128, 66, -128, 97, 0, -128, 127, -128, 127, 127, 127, 127, 59, -128, -43, 55, 127, 127, 127, 127, 37, 45, 57, 127, 127, -18, -128, -128, 127, 127, 85, -53, -128, -128, 127, -34, 70, -128, -108, -71, -128, 127, 43, -80, 127, -128, 127, -101, -86, 127, -23, 127, 127, 127, 127, -128, -33, -128, -128, -128, -128, 59, 127, 127, 64, -128, 17, -128, 48, 127, 127, -50, 96, -48, -112, 78, 43, -128, 127, -29, -128, 127, -128, -128, 81, -128, -128, 127, -128, -15, 127, 127, 127, 127, 127, -128, -128, 24, -128, -128, 34, -128, -1, 127, 127, 127, 127, 49, -93, 0, 127, -7, -128, 60, 73, 127, 127, -128, 127, 127, -18, 24, -128, -128, -128, 21, 127, 127, 127, -31, 127, -103, 31, 127, -42, 127, 44, 127, 127, -128, -128, -65, 127, 127, 127, -63, -128, -128, -128, -17, 127, 127, -87, -69, -21, 127, 95, 127, 127, -128, -123, -128, -128, -128, -108, -128, 127, 34, -128, -29, -128, -117, -96, -128, -128, -128, -128, -26, -96, 127, 44, 127, 22, -128, -118, -11, -75, 127, -66, 127, 13, -128, 127, -128, -128, -49, -128, 119, 127, 12, 127, 127, 127, 127, -16, 127, 127, -57, 24, -128, -128, -128, -128, -108, 90, 127, 24, 127, -128, -128, 127, -128, 107, 127, -71, 127, 33, 127, 127, 127, 55, 127, -128, -128, -128, -128, 127, 127, 69, 127, -128, -128, 127, -128, 52, -128, -128, 75, 111, 127, 127, -128, 65, -91, -128, -39, -96, -128, 127, -63, 52, -44, 97, 127, 127, 127, -128, -128, -92, 33, 127, -128, -18, -33, 127, 127, 127, 127, 119, 114, 127, 95, 127, -78, 122, 127, 26, -128, -26, 75, -128, 127, -39, -128, 106, -128, 117, 116, -92, -128, -128, -60, 17, 69, 75, -128, -128, 127, -22, -128, 127, -128, -31, 127, 108, 127, 127, 108, 64, -128, -128, -128, -128, 57, -100, -128, -128, -88, -33, 127, 5, 127, 127, -128, 24, -128, 113, 127, -23, 127, 44, 16, 127, 96, 127, 127, -128, 86, -128, -128, 16, 36, -128, -5, -128, -26, -128, 111, 127, -128, -112, -128, -123, 127, 127, -48, -73, -128, -10, -113, -128, 127, -128, -18, 127, -128, 127, -47, 73, 127, -123, 127, -128, -17, 127, -128, 127, -128, -128, 127, -100, -128, -63, -128, -128, -49, 11, 127, 127, 127, 100, 93, 34, 32, -106, 127, 127, -53, -128, -106, 114, 87, 127, 70, 108, 127, -2, 127, -128, -86, -128, 106, 50, -128, 127, -128, 22, 102, -128, -90, -128, 76, 127, 86, 127, 127, 127, 47, -128, -128, -124, 12, 127, 122, 88, -81, -128, -15, 127, 24, -93, 117, -87, 127, 21, -100, -128, -123, -34, -69, 127, 26, 127, 127, -122, 127, -128, -11, -42, 66, 70, 127, 127, -128, 127, -119, -128, -39, 24, 92, 91, -128, -32, -128, 127, -32, -103, 127, -128, 107, -44, -128, 127, 79, -128, 122, -116, -103, -36, -128, -39, -64, 15, -103, -128, -128, -128, -128, -90, 107, 127, 37, 127, -38, 127, -10, 127, 127, -128, 127, 116, 60, -128, 65, -128, 33, -36, -128, 127, 101, 24, -128, -96, -128, -49, -128, -128, 127, -121, 127, -57, -128, 70, -128, 127, 127, -128, -45, -128, -128, -7, 127, 127, 127, -128, -42, -112, -128, 127, -128, 78, 21, 49, 127, 127, 80, 127, 7, -96, 127, -80, -26, 127, -128, -128, 98, 86, 127, 127, 68, 127, -128, 127, 127, 127, 7, 127, -128, 70, 127, -128, 127, -128, -87, 127, 22, -15, 127, -92, -128, 10, 74, 127, 127, 127, -128, -128, -13, -128, 53, 17, 15, 127, 127, 127, 127, 127, 127, 116, 73, -128, -42, -128, -63, 127, -128, -38, -128, -128, -113, 101, 127, 127, 70, 127, 127, 127, 54, 127, -128, 127, -54, 81, 42, -27, 127, -103, -16, -92, 42, 18, -128, -128, -128, 12, -33, -16, -50, -118, -128, -114, 127, 127, -11, -75, 11, -128, 127, -102, 93, 74, -113, -38, 127, -128, 39, 76, -128, 28, -128, 127, -127, 127, 127, -22, -128, 85, -128, -58, 32, -128, -128, -128, -128, -15, 127, -109, 127, 127, -13, -16, -128, -5, -128, 0, 6, -128, -38, 127, 127, 127, -128, -128, 127, -128, 127, 23, 76, 127, 73, 127, 127, 127, 98, 127, -55, 127, 127, -128, 127, -128, -107, -128, -128, -50, -128, 0, 33, 127, 127, -43, -128, -54, -128, -38, 127, 127, -87, 114, -128, -128, -15, 127, 45, -5, 108, -128, 116, 22, -128, 127, 127, 127, 78, 0, -128, -128, -128, -8, 127, 37, 127, 127, -128, -128, -29, -128, 11, 10, -128, -108, -92, 127, -122, 31, 127, -128, 127, 127, 93, 127, -87, -128, -109, -5, -128, -76, 127, -128, 88, 127, 33, 127, -8, -128, 127, -47, 127, 124, -128, 43, -117, -10, -128, 43, -88, -128, 59, -128, 116, 127, -128, 85, 22, -128, 127, 101, -68, -92, -90, -124, -128, 79, -81, -128, -128, 17, -128, -34, 108, -128, -11, 127, 127, 127, 127, 16, -128, -128, 27, 17, 127, 127, 127, 127, 64, 127, 127, 60, 127, -128, -128, -128, -60, 29, -128, 127, 55, -65, -17, -128, -128, -128, -128, -128, -128, -128, 127, 127, -128, 127, -128, -128, 15, -128, -124, -128, -128, -128, -128, 127, 127, 48, -36, -128, -128, -128, -43, -128, -128, -128, 127, -63, 127, -52, 71, 127, -96, 127, -128, -128, -128, -128, -108, 91, 33, 127, -116, -93, 127, 101, 127, 0, 16, 50, -113, -128, -36, -128, -128, 127, -128, 127, -128, -68, 127, -128, 127, 48, 22, -91, 50, 127, -31, -73, -55, -128, -128, 127, 127, 24, 33, -128, -128, -128, 117, 127, 52, -128, -128, 16, 48, 59, 127, 127, -45, 52, -128, -128, -52, -128, -128, 127, -128, 124, -7, -128, -21, -117, -128, -128, 127, -128, 90, 113, -128, 28, 95, -128, 36, 127, -128, 127, 24, 127, 60, -37, -128, -128, 127, 127, 127, 85, -128, -128, -128, -128, -15, -39, -128, -128, -128, -128, -16, -128, -32, -98, 127, 29, 55, 8, -21, -128, 86, -128, -76, -74, -128, -70, -128, -128, 127, -128, 127, 127, 127, 127, 12, -7, -128, -8, -52, -128, 85, -128, -128, 127, -28, 86, 127, 58, 43, 24, -128, -128, 22, -128, 54, 127, -128, 127, -128, -128, 127, -128, 127, -88, -128, 92, 127, -32, 127, -128, -128, 127, 127, 127, -91, 36, -128, -107, 127, -128, 69, -128, -24, 78, 127, 79, 127, 57, 127, 127, -128, 127, 127, 111, 127, -64, 116, 127, -128, 53, -128, 108, -128, -70, 127, 15, 127, 127, 127, 5, 127, -128, -128, 103, 70, 127, 127, 127, 97, -114, 127, 127, -128, 127, -128, 28, -128, -128, 50, 88, 127, 127, 127, -121, -128, -27, -106, 127, -33, -128, -128, -63, -128, 59, 100, 53, -17, 39, 127, -38, -31, -90, -128, 31, 1, 127, 1, -57, -87, -128, -128, -128, -128, 100, 13, -93, -32, -128, -128, 24, -112, -128, 17, 127, -128, -36, 38, -108, -128, -128, -97, -23, 85, 127, 127, 86, -10, 117, 127, -2, 71, 127, 11, 127, 52, 33, 127, 21, 127, 127, 127, -128, -128, -103, 78, 127, 127, -85, -128, -128, -121, -128, -34, 127, -127, 127, -86, -74, 127, 127, 127, 127, 127, -63, -128, -85, 68, -15, 127, 127, 18, 127, 127, 50, 66, -128, -117, 127, 127, 107, -54, -128, 127, 57, -73, -128, 17, -128, 127, 127, 42, 117, -47, -128, 127, 8, -75, 32, -128, -128, 17, 75, -107, 95, 127, 127, 95, -128, -128, -128, -3, 127, 70, 80, 57, 127, 23, 127, 127, -128, -128, 17, -109, -128, 47, -128, -128, -69, -102, 127, 127, 127, 127, 127, -119, 74, 97, 23, 127, 127, 127, 127, 1, 127, -128, 42, -112, 15, 127, 127, 78, 127, -128, -128, 24, -128, -128, 127, -12, 65, 127, -80, -96, 68, -128, 100, -91, -52, -85, -68, 86, 17, 127, -128, 127, -26, 23, 113, 127, 127, 127, 127, 127, -128, -34, -128, -128, -128, -128, -88, -7, 127, 28, 127, 127, -128, -53, 42, -128, -128, -128, 93, 87, -44, 37, -128, -128, -111, -59, -103, 111, 127, 127, 127, 127, 127, 127, -60, 79, -128, -34, 127, -92, 127, -128, 112, -48, 127, 122, -128, 114, -128, 54, -36, -43, 127, 47, 127, 127, 106, 127, -128, 127, -128, 93, -128, -128, 127, 111, 127, 127, -85, 127, -113, -128, 127, -128, -128, -6, -128, 38, 45, -128, -15, -128, -128, -128, -128, -128, -116, -128, 101, 127, -128, 127, -71, 127, 127, 37, 118, 65, 127, 127, 49, 118, 127, -128, 96, 122, -39, 127, 127, 127, 127, -39, -128, 1, -118, -128, -128, -128, -75, -128, -128, 127, -47, -100, -128, -128, -128, -101, 127, 127, 127, 127, 127, 127, -38, 53, -75, 64, 127, 127, 36, -128, -117, -128, 127, 127, -111, -10, -98, 33, 97, -128, -128, -26, -128, -55, 106, 127, 114, 80, 127, 124, -18, -38, -128, 28, -28, -128, -18, -128, 127, -128, 127, 34, -128, 127, -39, 127, -128, -128, 5, 64, 127, 127, 127, 127, -128, -128, 127, -70, 38, 127, -107, -43, -58, 127, -128, -2, 58, 28, 76, 127, 114, -128, -128, -118, 127, 127, 127, 53, -128, 38, -128, 127, 127, -128, 127, -107, 36, 127, 127, 87, 88, 127, -128, 127, -107, 127, 18, 5, 127, 127, 33, 12, 103, -113, 127, -128, -128, 127, -116, -88, 127, -128, -128, 91, -36, -128, -106, -128, -128, 127, 16, 127, 127, 127, 127, 95, 28, -119, -128, -44, 29, -128, 29, 127, -128, 127, 127, -128, -53, -17, 33, 127, 127, 31, 87, 127, 127, -128, -91, 127, 59, 127, 127, -121, -128, -128, -128, -49, 127, 127, -26, 39, 79, 31, 43, -128, -28, 127, 24, -128, -128, 1, -17, 127, 85, -128, -43, 127, 98, 127, 17, -66, 127, -128, -16, -43, 127, 127, 127, -123, -128, 23, -22, 127, 127, -113, 60, -128, -39, 127, -128, 127, 127, -6, 127, 127, 127, 127, 127, 127, 127, -128, 73, 64, -47, 127, 127, 48, -128, 127, -55, -128, -44, -97, -65, 103, 127, 127, 102, 127, 109, -128, -113, -65, -128, 114, -118, 48, -128, -43, 7, -128, 57, -12, 127, 127, 55, -128, 8, -63, 71, 127, -55, 59, 127, -73, -42, 127, -128, -54, 34, 13, 127, 13, 1, -128, -128, -128, 5, 24, -128, -22, -111, 127, 127, 127, 36, -128, 79, 53, -27, -5, -128, -128, -73, -128, 127, -80, -58, 127, -57, 127, 127, 58, -63, 45, -128, -128, 119, -128, 76, 50, 54, -128, 127, 127, -128, 127, 79, -128, 127, -128, -97, 38, -128, 127, -22, 127, 127, 127, -97, -50, 31, 93, -128, 47, 127, -128, 21, 127, -128, 127, 47, -118, 127, 36, 127, 127, 6, 127, -128, -128, -128, -128, -128, -128, -128, -128, -101, -128, -118, -128, -128, -85, 127, 127, 127, 12, -128, 80, -128, -113, 127, 0, -100, 127, -128, -26, -128, -128, 127, -128, 58, 127, 127, 127, 10, -128, -128, 87, 127, 127, 70, -128, -128, -128, -128, -128, -128, -15, -128, -128, 127, -128, 95, 127, 127, 127, -28, -128, -128, -128, 71, 127, 127, 127, 127, 127, -128, -113, 127, -128, -128, 127, -90, 0, -128, 76, -128, 127, 78, 1, -128, -123, -103, 54, 127, -103, 3, -78, 85, 127, 21, -128, -124, -63, -38, -78, -128, -128, -128, 127, -128, -29, -52, 127, 26, 34, 17, -128, -128, -119, -128, -128, -128, -128, -128, 127, -106, 127, -128, -86, 127, 21, 127, -78, -21, 116, -128, -128, -63, -128, -128, 8, 127, -18, 127, 2, -128, 76, 18, -128, -97, 1, 27, 127, 127, -49, 38, 127, 0, 28, 87, 127, 112, 127, -32, 3, -128, -128, 7, 36, 69, 114, 127, -128, -18, 70, -44, -38, 127, -21, -128, -2, -128, 127, 127, 127, 127, -128, -44, -128, 85, 102, -128, -50, -27, 127, 127, -43, -128, -128, -128, 29, 17, -128, -101, -100, 2, -128, 100, 127, -128, 127, 45, 127, 127, 127, -50, -128, -128, -98, 127, 127, 24, 127, -128, 118, 127, -103, 127, -128, 127, 33, 39, -6, -98, -128, 42, -28, -128, 127, -128, -128, 102, 127, 119, 113, -22, 28, -23, 96, 127, 45, -2, -128, -128, -128, -128, -38, 127, 127, -128, 127, -128, -128, 127, -128, -128, -128, -128, -113, -79, 127, -124, 75, -31, 127, -87, -128, 127, -128, 121, 127, 127, -17, 127, 63, 127, 127, -90, -69, -128, -128, 100, 127, 109, 127, 127, -128, 2, 109, -128, 2, 8, 127, 127, 54, -65, -50, -1, 31, 31, -128, -128, -128, -128, 68, -128, 75, 127, 127, 45, 127, 59, -128, -39, -128, -101, 127, 91, -17, 127, -68, 127, 127, 75, 127, 13, -128, 127, -128, -114, 127, -128, 127, 96, -58, -15, 127, -128, 49, 127, 29, 111, 127, -29, 121, 69, -128, -128, -128, -18, -128, -116, 90, 127, 127, 127, -79, -17, 127, 34, 127, -76, 127, -55, -128, 106, -128, -93, -128, -128, -111, 127, 127, 127, 127, 127, -101, -128, -87, -73, -128, -128, 45, -128, -128, -28, -48, -128, -38, 122, -128, 127, -128, -128, -98, -128, -128, -128, -73, -13, -50, -12, 127, 16, 118, -27, -69, -68, 127, -76, 127, 91, -128, 127, -128, 127, 103, -128, -32, -128, 127, 127, 127, 127, 127, 109, -16, -128, -128, -128, -128, 127, 12, 127, -60, -128, -34, -75, 0, 127, -97, 127, 121, 127, 127, 127, -1, -98, 127, 127, -103, -96, -12, 70, -18, 8, 127, -113, 127, -24, -24, 127, 78, -78, 108, -128, -91, 127, 127, 55, 127, 127, -44, -39, -128, -128, -128, -128, -111, -38, 127, 127, 127, -90, -128, -128, 64, 43, -128, -65, -128, -128, -128, -128, 127, 127, 127, -128, -85, 7, 127, 127, 127, 127, -1, -128, -128, 38, 27, 127, 127, -44, 127, -18, -8, -63, 127, -65, 127, -2, -128, 27, -128, 118, -128, 47, 108, -102, 127, 98, -128, -117, -70, 109, 48, 6, -113, -128, -86, -128, -60, 3, 60, 127, 58, 118, 47, 127, -102, 106, -101, -128, -21, -49, 127, -128, 127, -114, 11, -128, 109, 86, -29, 127, -128, -47, 127, -57, 10, 127, -76, 93, 127, -128, 127, 15, -128, -63, -128, -128, 127, -39, 127, 127, -128, 6, -128, -128, 127, 127, -107, 127, -47, 68, 32, 127, 118, 80, 39, -128, -66, -128, -128, 127, 13, 28, -128, -128, 49, 127, 2, 127, 127, -17, 127, 127, 127, 127, 127, -76, 127, 12, 117, 66, -128, -128, -12, 81, 24, -128, 6, -128, -59, -63, 28, 127, 127, 127, 112, -128, -128, -128, 127, 93, -119, -128, -53, 127, 100, 127, -128, 7, 127, 32, -128, -33, 102, 127, 38, 15, -128, -128, 107, -97, 127, 127, -128, 127, -128, -49, 28, -128, -29, 127, 88, 127, -5, -21, 3, 127, 15, -58, -128, -128, 127, 50, 26, 127, 38, 127, 123, 127, 127, -48, 127, 106, -128, 127, -128, -128, 127, -128, 0, -128, -128, -24, -128, -128, -103, -128, 113, 127, 103, -119, 127, -86, -38, -74, -32, -15, 127, 127, 127, 127, -6, 127, 103, 127, 127, 81, -15, -128, -128, -121, -128, -128, -128, -128, 52, 127, 127, 127, 2, -128, -103, -108, 3, 127, -15, -100, 127, -128, -63, 127, -128, 44, 118, 127, 119, -34, 127, -128, 31, 127, 127, 58, 121, 127, -128, 127, -117, -128, 127, -79, 65, 27, -128, -6, -3, -128, 75, 91, -128, 127, -6, 109, 114, 17, -81, -128, -81, -1, 127, 127, 127, 127, 127, -128, 93, -86, -43, -17, -24, -128, -128, -96, 127, 127, 119, 127, 26, 91, -64, -17, 3, 49, 127, 90, -88, 42, -128, -29, -128, -128, 127, 11, 127, -73, -21, -90, 127, 88, -64, 127, -128, 37, -128, -128, 127, -68, -128, 127, -53, -78, 127, -128, -128, 127, -128, -42, -112, -128, -117, -128, -128, -128, -96, -128, -81, -128, -128, 26, -112, 70, 32, 16, 29, 113, 127, 127, 127, 117, 18, -128, -2, -92, -5, -75, -128, -128, 10, 127, -108, 127, -128, -128, -128, 59, 109, 32, 127, -111, -7, 127, 127, 127, 127, -48, 97, -39, 127, -29, 127, -128, -13, -128, -128, 127, -66, -16, -128, -128, -128, 127, -5, -74, 54, -128, -128, -86, 68, 60, 31, -90, -128, -128, -128, 127, -37, 127, -128, -128, -79, 91, 127, 127, 127, 98, -128, 31, -128, 127, 33, 127, -1, 34, 102, 37, 63, 127, 39, -128, -12, -128, -128, -118, -128, 127, 127, 5, -95, -128, -63, -128, -68, 102, 127, 43, 127, -34, -23, -123, 127, -109, 127, -2, -128, 127, -124, 127, -112, 49, 88, -128, 22, -128, -128, -23, 44, 127, 127, 127, 28, -128, -128, 13, 54, 127, 106, -121, -128, -128, -128, 127, -128, 53, 127, -128, 79, 127, -13, 127, 127, 31, -17, -128, 127, 32, 108, -128, -65, -128, 16, 124, 3, 8, -128, -128, -128, -128, -128, -128, -108, 0, -85, -128, 127, -128, -128, 127, -103, -128, 127, 48, 7, 57, 58, -119, -54, 127, -128, 57, -128, -128, -128, -128, -128, 127, -65, 26, -122, -38, -128, -128, 127, -128, -57, 127, 6, -23, 127, 101, 71, -13, -33, 127, 127, 127, 127, 127, 117, -128, -128, 127, -128, 127, 127, -128, 1, -39, -128, 85, 54, 12, 127, -128, 60, -128, -128, 2, 119, -128, 127, -108, -80, 127, 59, 64, -128, -60, -128, -13, 127, 109, 7, 100, 119, 127, 127, 45, -109, -10, 127, 45, 127, 12, -123, -116, -128, 127, 127, 3, -31, 127, 32, 24, 124, -128, -128, -128, -128, -128, -100, 43, 127, 127, 127, -124, -8, -128, -128, 127, -92, 127, 127, -87, 127, -49, -128, 69, 73, -128, -23, 124, 127, -31, 127, 68, -128, -17, -128, 81, 127, 127, 127, 127, 127, 123, -28, -128, 57, 76, -66, 22, 53, -39, -128, -128, 127, -95, 1, 127, 44, 119, 53, -128, 127, -101, -128, 16, -128, -128, -103, -128, 124, -128, -26, 108, 93, 37, 127, 12, 127, 127, 127, 127, 127, 76, -128, 49, -128, -128, -128, -128, -1, -128, 127, -123, 38, 127, -128, 29, 127, -52, 44, 102, -70, -128, -64, -128, -128, 127, -128, 122, 113, 43, -15, -128, -55, 113, 127, 127, 85, 127, -128, -101, 24, 45, 127, 127, 127, 127, 127, 127, -122, 43, 108, -128, 127, -93, 93, 64, 75, 44, -128, 18, -128, 45, 127, -69, -128, -128, 127, -97, 57, 22, -64, -44, -127, 18, -116, 48, -128, -112, -128, -128, 76, 24, 127, 53, 127, 127, -128, 127, -128, -128, 80, -79, 127, 127, 127, 127, 127, 127, -37, -128, -111, 70, -128, 127, -128, 127, -45, 21, -128, -96, 127, 79, 127, 86, -68, 48, 127, 127, 127, 127, 127, 127, -69, 127, -128, -69, -31, -11, 127, -31, 10, -128, -87, 69, -128, 127, 42, -128, 37, -16, -128, -128, 90, -128, -128, 127, -128, 111, 68, -33, 127, 127, 88, -64, 127, 58, -80, -128, -128, -75, -114, 44, -128, -128, 1, -128, -128, -75, -128, -119, 42, 7, 127, 127, 53, -128, -53, -128, -128, 33, 127, 90, 127, 127, 113, -128, 28, -87, 10, 127, 127, 127, 127, -75, 31, 127, 127, 127, 127, 28, 24, 127, 127, 127, 127, 127, -68, 127, -5, 69, -1, 50, 127, 11, 127, -128, -128, 43, -58, 127, 127, 106, 123, 102, 90, 127, 42, 23, 127, 86, 127, -32, 127, 18, -1, 58, -128, -52, 57, 127, 127, 39, 127, -128, 127, 127, -128, 21, 21, -128, -128, 63, 127, 45, -86, 101, -128, 85, -128, 8, -69, 75, 127, -128, 127, 127, 96, 127, 24, 127, 114, -128, -128, -128, 88, 127, 37, 127, 127, 101, 127, 127, 113, -69, 17, 127, 127, 97, 127, 74, 11, -111, -128, 0, -128, -53, 127, 127, 127, 127, 127, 98, -16, -128, 39, -128, -69, 11, -71, 127, 127, 106, -16, -128, -128, 127, -128, 127, 127, -128, -32, -128, -128, -128, -128, -128, -63, -128, -128, -1, 127, 0, 127, 21, -128, -81, -128, 127, -50, 86, 127, 127, 127, 127, -38, 8, -128, -128, 127, 95, 127, 50, 127, 114, -128, 127, -128, -128, 127, 127, 79, 127, 127, 43, -128, -128, -71, -43, 127, 127, 75, 127, 127, 38, 127, 70, -128, -128, -70, 88, -13, -70, 64, -128, -128, -128, -128, -128, 114, 66, 127, -107, 101, -81, 96, 127, 127, 127, 34, -128, -128, -128, -128, 73, -128, 127, -76, -122, 127, -31, 127, 48, -109, -98, -18, -69, 127, -37, -128, -5, -17, 127, 127, -68, -128, 39, -66, 127, 118, -128, 127, -57, -128, 79, -128, -128, -128, -71, -95, -128, -5, 127, 127, 127, 127, 127, 127, 127, 127, 127, 22, -128, 43, -64, -128, -128, 43, -96, 127, 127, 100, 127, 31, 127, 127, 95, 127, -128, -128, 59, -100, -18, -68, 92, 122, 127, 1, 76, 127, -2, -34, 127, -128, -59, 58, 127, 127, 127, 127, -119, -128, -23, -128, -17, 127, 24, 127, 127, 127, 127, 127, 6, -128, 10, 65, 127, 123, 109, 127, -118, 92, -128, -128, 127, -128, 88, -114, 44, 103, -128, -23, -128, -13, -15, 127, 127, 15, 127, 127, -128, 127, 49, 101, -90, -128, -122, -114, -36, -128, -128, 127, -122, 127, -37, 127, 34, -128, -128, 2, -15, -64, -70, -128, -128, -52, 127, 127, 34, -81, -128, -128, -128, 114, 127, 0, 121, -36, 93, -50, 127, 127, -79, 127, 127, 65, -128, -34, -128, -128, 127, -128, -16, 92, -113, 127, 127, 0, -1, -128, -128, 127, 7, 93, 57, -128, -128, -10, -128, 13, -128, -2, -117, -34, 127, -128, 127, 127, -128, -8, 127, -80, -128, 127, -128, -48, 127, 127, 109, 127, 87, -2, 127, -128, 127, -22, -50, -26, -69, 13, -128, 93, -128, 127, -54, 1, 127, -128, -43, -1, -128, -95, -128, 58, 127, -128, 49, 80, 103, 70, 127, 3, -128, 74, 127, 127, -68, -128, 127, -29, -103, 127, -128, -128, -128, 73, -52, 58, 127, 43, 36, 5, -128, -128, -128, -79, 75, 29, 96, 127, -16, -128, -73, -8, -11, 96, -128, 59, -8, 2, 127, -128, 87, 127, 8, 127, 127, 127, 31, 108, 127, -128, 27, 109, -64, 69, 127, 127, -102, 127, -50, 127, 106, 127, 68, -21, -128, -128, -78, -128, 12, 127, 12, 79, 2, 10, 127, 31, -128, -96, -128, -128, 119, -128, 127, 21, -128, -117, -128, 53, -75, -128, 45, -128, -128, 81, 127, -39, 127, 127, 127, 127, 119, -111, -128, -128, 127, 88, 127, 127, -128, -87, -128, 8, -38, -128, -24, 42, 127, -80, 59, -128, -128, -74, -24, -128, -54, 75, 127, -85, 71, 127, 91, 127, 127, -128, -128, -128, 68, 127, 127, -107, -3, -128, -128, -128, -128, 28, 127, 127, 127, -81, -128, -128, -128, -128, -128, -128, -49, -128, 127, 127, 127, 127, 45, -70, -128, -128, -128, -128, -124, 17, 127, 127, 127, 79, -128, -128, -128, -128, 0, 127, 127, 127, 127, 32, 127, 127, 8, -96, -128, -10, 32, -128, 74, -66, -128, 24, -128, -128, -71, 29, 103, -63, -128, -58, 127, -128, 127, 127, 127, 127, 34, -32, -128, -128, -5, -128, -6, -128, -13, 44, -128, 127, -128, -128, 127, -11, 7, -21, -128, -76, -128, -128, 127, -92, -128, 127, -128, -128, -76, -128, 119, 79, -128, -128, 55, -128, 127, -32, 23, 127, -33, 31, -128, -16, 127, -39, 127, 47, -111, -128, -128, -128, -119, 127, -47, 127, 127, -44, 127, -128, -128, -128, 127, 48, 127, 96, -128, -128, -128, -13, 127, 127, -16, 90, -12, -128, 50, 127, 32, 127, 34, 48, 127, 127, 127, 108, 54, -128, 127, -128, 32, 127, 127, 127, 0, -128, -128, -128, -128, -128, -128, -128, -42, 70, 127, 127, 127, 127, 127, 127, 127, -79, -128, -5, 116, 26, 0, -29, -128, -112, -128, 1, 117, 38, 127, -102, -128, -128, 22, -55, -128, -57, -26, 60, 123, -24, -128, -128, -18, 64, -128, 108, 2, 127, 127, 127, 127, 127, -106, 127, -112, 5, 127, -128, 58, 70, -128, 13, -128, -128, -45, 0, 127, 127, -47, -128, -45, 59, -128, 127, -128, -128, 127, -128, 127, 127, 95, -37, 127, -128, -128, 18, -39, 127, 127, 45, 3, -128, -128, 117, 127, 127, 127, 127, -128, -128, -128, -52, 127, -128, 118, -128, -128, -48, -128, -90, -128, -128, 31, -128, 127, -78, -128, 127, -128, -55, 127, 127, -21, 127, 127, -28, 127, 127, 127, 127, -80, -128, 74, -128, 123, -36, 127, 127, -128, 34, -128, -127, 127, 127, -128, -17, -118, -100, 127, 127, 127, 127, 80, -128, -128, -128, -128, 127, 32, 127, 26, -93, -128, 127, -59, 127, 71, -128, -128, -128, -128, -70, 80, 127, 57, 127, 127, -5, -7, -128, 66, -128, -128, 127, -128, -128, 118, -81, 127, 127, 127, 127, 59, 127, -128, -128, -57, 127, -49, 127, 26, 114, 12, -128, -36, -128, 113, 127, 127, 127, -128, -128, 37, -128, 21, 127, -128, 127, -128, -87, 127, -121, 127, 7, 108, 43, -128, -128, -128, -33, -128, -39, 18, 127, 127, 127, 127, 127, -90, -128, -24, 127, -128, 127, -36, -128, 127, 37, 127, -128, -90, -52, 127, 127, 37, -88, -128, -31, -128, -116, 127, 2, -128, -97, -118, 127, 50, 127, 127, -76, -71, 76, -128, 127, 127, 127, 127, 127, 127, -128, 127, -22, -127, -128, -128, -128, 101, 127, 127, 86, 127, 127, 38, 127, -128, 127, -50, -17, 97, -128, 127, -128, -5, 127, -65, 127, -97, -92, -33, -33, 127, -108, -128, 34, -128, 87, -13, 127, 127, -128, 127, -18, -128, 96, 127, 107, 127, -128, -53, -32, -75, 127, -32, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, 26, -44, 8, 127, 86, 87, 90, 127, -59, -13, 127, -109, 127, 127, 81, -96, 11, -128, -63, -128, 10, -128, -128, 127, -128, -128, 79, -128, -66, -11, -128, -39, 127, 93, -1, -42, -36, -43, -128, 127, -85, 127, 66, 127, 100, -36, 127, -121, 127, -128, -128, -128, -128, -128, -128, 49, 127, 127, 117, -128, -128, -128, -118, 106, 52, 31, 69, -21, -128, 127, 117, 127, 21, -128, -128, -55, 127, -38, 127, -128, 1, 127, 127, 127, 127, 127, -128, -128, 44, 42, -8, 47, -128, -128, -128, -128, 29, 127, 66, 127, 127, 48, 127, -128, 86, -65, 127, 66, 127, -93, -108, 127, 31, -3, 70, -128, -17, -32, 127, -65, 96, 118, 37, 5, 108, 127, -128, 101, -128, -128, -128, -128, -76, -128, -128, 127, 127, 26, 7, 90, -32, -128, 5, 23, 107, 127, 96, 127, -128, 116, 127, -57, -12, -128, 5, -128, -93, 107, -128, 47, 127, 127, 127, 127, -29, 127, 127, -128, 60, 68, 58, 127, 127, 127, 7, 127, -128, -128, 127, -28, 127, -87, -16, 127, -68, 127, 127, -117, 98, -128, -18, 127, 127, -45, 27, -128, -128, -128, -128, -128, -74, -71, 29, -128, -128, -109, -128, -53, -128, -128, -128, -128, 127, 127, 32, -128, -128, -128, -128, -128, -128, -128, -65, 55, -128, -128, -78, -128, 29, 90, 78, 127, 127, -5, 127, 127, -121, 127, -128, 27, -37, -50, 22, -128, -128, -128, -128, -39, 52, 127, 127, 127, 127, 127, 127, 127, 65, 6, -128, -128, 0, -128, 65, -128, 70, -121, -18, 127, 12, -58, 127, -128, -81, -128, -128, -128, -128, -128, -71, -103, 57, 63, 27, 127, 127, -128, 127, -128, 18, 52, -128, -34, 5, -57, -128, -128, -128, 15, -21, 127, 127, 127, 127, 127, 10, 127, -128, 33, 50, 53, 127, 12, -128, -128, -50, -78, -128, -31, 103, 127, -124, 127, 90, -128, 127, -128, -70, 42, 107, -55, 93, 127, -128, 116, -128, 34, 127, -87, 73, -102, -128, -47, -1, 127, 127, -57, -15, 127, -17, 127, 127, -128, 96, -128, -128, 127, 45, 127, 127, -55, 112, 88, 127, 127, 127, 127, -128, -128, 112, -96, -34, 127, -128, 127, -54, -128, -55, -128, 3, 127, 127, -128, 66, -128, -26, -60, 91, 127, -128, 127, -128, 117, 15, 108, 127, 127, 116, -128, -128, -116, 42, 37, 127, -28, 127, 127, 87, 127, 127, -128, -128, 39, -128, 102, -60, -128, -2, -128, -128, -34, 108, 127, 127, 116, -27, 127, -117, 127, -16, 127, 127, 127, 11, -128, -114, -27, -74, -11, 127, 65, 127, 127, 127, -27, 45, 127, 127, 124, 127, 42, -128, 127, 127, 5, 127, 127, -128, -79, -114, -128, -5, 127, -8, 127, 127, -98, 127, 127, -128, 127, -128, -128, 127, -128, -15, 127, -49, -128, -24, -128, 39, -21, -45, -8, -128, 49, -68, -29, -118, -128, -18, -128, 38, -13, 127, 50, 127, 86, 127, 122, 127, 16, 127, -58, -21, 127, 127, 127, 127, 127, 127, -39, 127, 60, -90, 27, 109, 32, 127, 73, 127, 118, -73, -128, -15, 39, -128, 127, -128, -128, 0, 17, 54, -128, -22, 65, 0, 127, 127, 127, 127, -98, -47, 127, -64, 43, -128, -128, -128, -64, 127, 127, 127, 127, -100, 127, 48, -1, 32, -1, 127, 127, 127, -65, -128, -10, 85, 33, 76, -128, -42, 127, 127, 127, -128, -128, 97, -15, 127, -18, -128, -103, 127, 3, 127, -33, -65, -128, 112, 88, -128, 86, -128, 95, -69, -33, 28, 102, -23, 127, 111, 127, 127, -7, 127, -116, 127, 44, -54, 127, 127, 127, 31, -28, -117, 38, 42, 127, 127, 52, 88, -55, -128, -128, -128, -71, 127, -118, 127, 127, -91, 75, 127, -128, -103, 127, -128, 116, -111, 26, -73, -128, -63, -128, -3, 103, 127, 11, 63, 92, 127, 127, -6, 127, -128, 24, -128, 37, -36, -24, -47, -53, -128, -128, -128, -128, -21, 103, 127, 127, 112, 127, 113, -31, 50, -128, -128, -128, -12, 119, 127, 87, 42, -16, -128, -128, -92, -73, -128, 103, 127, -80, -80, 127, 34, -23, -74, -128, -128, -98, 127, 33, -128, 22, -128, -128, 127, 12, -128, 127, 63, -12, -128, -3, -128, -124, -128, -128, -100, 127, 127, -86, -128, 79, -128, -128, 127, -70, 3, 127, 127, 127, 127, 66, 127, 127, 33, 127, -36, -15, -128, 29, -128, 127, 127, 97, -128, -44, -128, 117, 127, -128, 52, -123, -75, -108, -88, 127, 127, -128, 68, -128, 78, 127, 81, 101, 79, 127, 32, 127, 29, -128, -128, 1, 11, -93, -43, -47, -128, 107, -87, 97, -32, -128, -128, -128, 127, 33, 127, -128, 109, 29, -128, -43, -128, -128, -95, 71, 78, 127, 127, 91, -128, 70, -128, -36, 6, -128, 7, 28, -76, 127, 127, -128, 127, -128, -128, 127, 127, 127, 127, -128, -128, -128, -128, -70, -128, 127, 42, -95, 127, -117, -96, -128, -128, -128, 127, -15, -15, -79, -128, 54, -95, -128, -128, 21, -128, 127, 47, -128, 74, -10, 86, 50, -128, -128, -5, -15, 75, -128, -87, 58, 2, 127, 16, 18, 119, -32, 127, 49, 127, -53, -32, 127, -128, 127, 127, -128, 96, 127, -78, 127, -54, -128, 66, 107, 127, 127, 127, 127, 114, -42, -87, -42, 16, 127, 127, 93, 127, 85, -87, 55, 102, 92, -128, -96, -2, -128, 33, 127, 33, 96, 127, -22, -26, 21, -128, -85, -69, -76, -128, -128, -128, -128, -128, -128, -128, -128, 127, -128, 54, -85, -128, 97, -128, 127, 31, 34, 43, -128, -42, -128, -60, 45, -128, 127, -128, -65, 47, -128, 79, -128, 69, -128, 127, -128, 127, -128, -13, -23, 127, -108, 93, 127, 127, 100, 127, -128, -128, 12, -71, 127, 93, 69, -128, 112, 1, -128, -27, -128, -96, -128, -128, 88, -116, 127, 127, 127, 127, 127, 127, -70, 127, -96, -106, 81, -128, 127, -73, 7, 90, 90, 127, 54, -128, -128, -128, 33, 43, -124, 127, 18, -128, 127, 58, -128, -5, -128, 68, -18, 121, 127, -128, 122, -49, 28, 127, 127, 127, 127, 0, -6, -111, 127, 127, 127, -128, -128, 0, -128, -79, -128, -128, 15, -128, -128, 127, -128, -128, -128, -22, -5, -37, 127, -128, -128, 127, 34, -128, -49, 127, -43, 97, -128, -13, 122, -38, -128, -128, 47, 55, 127, 127, -36, 127, -101, -128, 7, -98, -128, 29, 101, 23, -58, -21, 31, 127, 127, -8, 86, 127, 0, 127, -128, -98, -128, -86, 127, -70, -128, -111, -128, -18, 64, 127, 127, 15, 0, -128, -128, -128, -128, 127, 127, -91, 124, -117, 0, 81, 113, -128, 54, 127, -128, 127, -73, 127, 127, -38, 18, -38, 76, 127, 127, -128, -43, 49, -128, -70, -128, -117, 127, -36, 31, -128, 53, 10, -87, -128, -128, -128, -73, -128, 127, -128, -128, -128, -21, -128, -22, 127, 127, 127, 127, 127, -128, -128, 127, -128, 127, -31, -15, 127, -128, 122, -87, -128, -128, -128, -128, -128, 127, -128, 127, 55, -128, -58, 10, -128, 106, -95, -128, 12, -128, 85, 127, -100, -128, -57, -128, -18, 127, -127, 127, 127, -128, 93, 95, 92, 127, 66, -48, -128, -111, -128, -63, 127, 95, 127, 127, 101, 112 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
