-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb2425 is
end tb2425;

architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 22533;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
            2, 9, -2, -15, -16, -4, 13, 14, 18, -7, 7, -12, -20, -6     -- C1-C14
                                                      );
    signal scenario_input : scenario_type := ( -61, -123, -69, -88, 28, -31, -70, -68, -84, 83, 105, 74, -76, 10, -108, 26, 73, 21, 24, -1, 40, -62, -74, -85, -75, -126, -69, 4, 59, 51, -72, 83, 45, -102, -86, -8, -46, -78, 70, 96, -100, -67, -11, 30, -74, 50, -126, -109, 29, -4, 111, -29, -46, 74, -117, -26, 86, -107, -90, -41, 71, -75, 112, 84, 14, 98, -27, 12, -86, -96, -49, 127, 64, -15, -105, -109, 127, 103, -103, -63, -64, 74, -44, -5, 58, -79, -104, 6, 12, 57, 32, 1, 55, 58, 77, 6, 33, 31, -13, 113, 71, -6, -104, -37, -119, -74, 1, 111, 80, 57, -38, 12, 103, 98, -5, -80, 36, 84, 4, 49, -69, 29, -31, -88, -108, 16, 63, 20, 75, -43, 105, -15, 126, -112, 78, 123, 0, 127, -40, 37, 91, 12, -127, -61, -17, 11, 12, -111, -94, -75, -32, -60, 6, 45, -56, 25, -28, -58, 56, 69, -47, 86, -127, -72, 86, 19, -75, -90, -107, 104, 112, 51, 39, 5, 37, 19, -49, 13, 37, -16, 55, -48, 23, 13, -40, -5, -62, 58, 98, 98, -49, -117, -29, 52, -1, -31, -76, 4, -6, -77, -51, -24, -23, 90, 2, 99, -83, -44, 98, -41, -116, 0, -90, -61, -98, -31, -88, -106, -3, 71, -15, -24, 68, -128, 12, -35, 8, 105, 101, -58, 90, -58, -96, -47, 32, 126, -10, 69, -36, -97, 125, 2, 68, -90, -3, 0, -45, 27, 101, 98, -88, -126, -49, -105, 119, 56, 116, -66, -97, -50, 88, -97, 32, 7, 126, 38, -22, 79, 6, 30, -31, -77, 72, 4, -77, 76, 81, 79, 85, -65, 2, -45, -85, 87, 85, 7, -103, -81, -72, 116, 114, 65, -98, 76, -49, 99, 25, -110, 79, 70, -45, 3, -78, -70, -7, 115, 106, 51, 7, 75, -107, -34, 96, 32, -85, 101, 93, 22, 11, -37, -110, 9, -101, -101, 81, 95, -61, 125, -50, 73, -63, 84, -84, -101, 111, 54, 86, -32, -88, -64, 55, -60, -63, -78, -118, 24, -76, -40, 120, -50, 12, -50, 30, 1, 11, 62, -87, -89, -14, -33, -17, 113, -98, 75, -31, 122, 88, -20, 3, -19, 79, -9, 124, -27, -3, -83, 104, -51, -30, 121, 112, 26, 98, -31, 59, 26, 72, 89, -76, 13, 38, -6, 96, -24, 25, 41, 24, 80, 42, -42, -15, -9, -44, -16, -103, 74, -51, -53, 62, 22, 68, -92, 126, -120, 39, 92, 35, 20, -13, 107, 55, 78, 17, 115, 116, 82, 49, -126, -85, 7, 44, 2, 113, -18, -39, -115, -76, -119, -5, 51, -33, 13, 79, -43, 124, -73, 22, -36, -50, -33, -111, -104, -76, 48, 1, -62, 90, -85, 87, -93, -103, 49, 50, 88, 63, -2, -41, 109, 84, -115, -58, -84, -109, 110, -58, -24, -56, 95, 20, -40, 120, -71, 15, -46, -108, 81, 72, -51, 85, 43, -84, 88, 84, 54, -53, -50, 56, -74, 73, 120, -52, 56, -55, -23, -40, -88, -88, -4, -98, 15, 120, 88, 108, 95, -67, -113, 3, 36, 127, -92, 87, 8, 65, 123, -98, -33, -104, -30, 95, 59, 61, 42, -4, -20, -46, -16, -62, -83, 53, -82, 58, -28, -86, -11, 38, 25, -67, -96, -73, 85, -97, 73, 31, 19, -34, 100, -33, -100, -107, 11, 17, 30, 119, 77, -56, -96, -85, 93, -70, 13, -37, 6, 110, -111, 127, -90, 65, 48, -1, -50, 64, 111, -56, 83, 87, 124, 21, -84, -26, -97, -30, 12, 94, -40, -56, 105, -16, 31, 26, -40, -85, -6, -100, -34, 94, 93, 59, -49, 11, 83, 95, -8, -49, -47, -105, 94, -111, 19, -56, 112, -64, -20, -64, 90, -33, 66, 127, 19, -97, -18, -37, 32, 63, -52, -87, -62, -107, 53, 83, -50, -61, -111, 126, -42, -16, -100, -119, -128, 77, 34, -74, 40, -118, 62, 70, 26, 104, 57, -30, 124, -37, -121, -30, -47, 34, -20, -97, 61, -113, -32, 32, -38, 126, -43, -7, -110, 68, 38, -41, -21, -75, 106, 65, -74, -39, -60, 48, 7, 110, -58, -11, -72, -13, 35, 52, -111, 48, 11, -12, -78, 82, 120, -43, 126, 15, 7, 65, 30, -11, 97, -122, 31, -63, 86, -66, -68, 23, 108, 100, -29, 36, -63, 14, 38, -70, -24, 99, -50, 30, -71, 70, -121, -51, 32, 82, -47, 107, -58, 121, -101, 100, -56, 95, -45, 42, 22, -40, -100, 105, 104, 127, -90, -75, -84, -67, 91, -116, -120, 82, -1, 7, -10, -110, -64, -92, 38, 19, -87, -16, -6, -2, -16, -63, 19, -48, -9, 11, 125, 121, -71, -127, 83, -102, -59, -121, -54, -91, -83, -35, 55, 110, -12, 16, 110, -101, 4, -34, 14, 22, 68, -109, 96, 15, 82, -85, 2, -47, 33, 91, -35, 120, -87, -115, 9, 16, 43, 14, 77, -75, 7, -109, -122, 123, 74, 28, -22, -86, -113, 125, -52, -23, -104, -126, -36, -11, 117, -80, -61, -91, 21, 39, 78, 17, 18, -18, 108, 66, -58, 109, -21, 40, -116, -20, 114, -13, 48, -104, 82, 89, -121, 31, 41, 119, -3, -41, 34, -75, -83, -64, -102, 32, -75, -24, 97, -35, -61, -4, 53, 57, 109, 59, 118, -90, 6, -85, 119, 21, -89, 79, -127, -18, -6, 127, -128, -25, -101, 33, -19, 97, -53, 118, -34, -59, 83, 37, -60, -39, -109, -41, 99, -45, -111, 69, 38, 70, -102, 43, 119, -105, 26, -8, -79, 113, 87, 72, -67, -26, 6, 3, -16, -43, -82, -113, -118, -39, -99, 109, -17, -104, 84, -58, -33, 119, 110, -22, 95, -124, 26, 100, -106, 123, 31, -49, -103, 54, -72, -114, 35, 106, 9, 121, -58, -51, 65, -55, -100, -127, -90, -106, -47, -66, 95, 88, -90, 89, 117, 98, 97, -28, -84, -61, 121, 52, -83, -123, -41, -34, 111, 43, -126, -54, -1, 85, 59, 94, -25, -92, 30, -88, -6, -22, -55, 115, 72, 92, -46, -9, -64, -110, -42, 80, 92, -76, -70, 22, 58, 47, -127, 63, 90, -43, -80, 51, 69, -8, 119, 98, -34, 62, 125, -22, 20, -64, -87, 48, 79, -27, 106, 79, 92, 56, -1, -7, 21, 110, 28, 76, 40, -16, -102, -89, -104, 59, 44, 52, -72, -111, 75, 0, -43, -122, -48, 66, 39, -59, -79, -124, -66, -86, -57, 69, 127, -74, 5, 45, -106, -63, -94, 109, -44, -69, -49, -6, -13, 82, 10, 43, -100, -82, -122, 124, -12, -22, -107, -24, 26, -19, -42, -106, -48, 73, 92, 33, -68, 84, 40, -8, -10, -53, 126, -44, -18, 101, 99, -88, -111, -37, 125, -124, 84, -84, -31, -117, -11, -36, 52, -121, 78, 35, -74, 126, -81, -96, -81, 100, 47, -110, -21, 58, 112, -107, 119, -124, -9, 27, 21, 83, 98, -126, 90, -22, 122, 74, 41, -30, -29, 12, 88, -3, -110, -18, 91, 30, 112, -105, -89, -33, -52, -126, -1, -27, -58, 70, 9, -126, 126, 74, 62, -1, -13, 45, -118, -28, -96, 62, 91, -8, -87, 119, 74, -127, -76, -80, 39, -12, 113, 90, -80, -125, -72, 72, -52, -67, -61, 14, 95, 84, -6, 64, 28, -41, 8, -99, -9, -123, -24, -15, 91, -77, -101, -50, 88, 60, -19, -54, 116, 99, -108, 120, -44, -56, -82, -45, 40, -107, 82, -67, 63, 93, -77, 1, 84, -98, 4, -50, 27, -24, 40, 11, 61, 10, 27, -2, 84, -120, -123, 108, -31, 115, 35, -118, 106, 104, 68, 85, 30, -1, -28, 72, -37, 14, 7, 52, 89, -5, -31, -84, -69, 14, -46, 50, -118, 62, 86, -59, 43, 2, -8, -47, -111, -38, -110, -47, 48, 111, -79, -50, -16, -121, -32, 34, 98, -70, -120, -69, -52, 7, 32, 112, -90, 76, -72, 7, -50, -43, -43, 82, -58, 51, 85, -18, 8, 71, 96, 103, -69, 50, 70, 45, 103, -27, -128, 32, -6, -43, -20, 10, 77, 75, 7, 84, 27, 13, 25, 35, 89, -57, 113, -44, 12, -28, -86, -61, 68, -60, -24, 37, 94, 41, 48, 96, -118, -119, -18, -42, -75, -105, 60, -109, 84, 102, -82, 45, -2, 26, 15, 40, -13, 64, 20, 66, -90, 69, 61, 2, -24, -66, -11, -59, 76, 28, 60, 92, 20, 57, 94, -102, 76, 58, 50, 126, 122, -110, -94, 78, 55, 117, 124, -17, -8, -56, 67, -70, 91, -111, 103, -81, 31, 100, 12, 52, 94, -110, 31, 5, -62, 120, -47, -76, -106, -109, -19, 123, -14, -88, 126, -10, -20, 56, 88, -97, 87, -30, 56, -87, -53, -113, 10, -29, 107, 115, 114, -91, -48, -117, -21, 117, 13, -42, 3, 108, 108, 119, 75, 83, -52, 6, -21, -116, 49, 34, 74, -48, 120, 113, 87, 88, 126, 36, -40, 98, -51, 63, 44, 68, 22, -124, 117, 29, -18, 104, -49, 103, -74, 9, -69, 59, 56, 19, 5, 75, -62, 29, -21, 39, -104, -19, 86, -2, -53, -86, -60, 125, -11, -94, 116, -87, -86, -112, -101, 45, -88, -31, -43, -41, 72, 20, 73, 33, -26, 25, -25, 63, 51, -26, -35, 19, 96, 109, 50, 127, -88, 88, 14, 124, -34, -54, 105, -56, -9, 88, -1, 41, 65, 9, 93, -121, 76, 54, -68, -85, 10, -70, 87, -62, 34, 68, 35, 27, 32, -91, 114, -100, -32, 21, 99, 106, 6, 61, -32, 67, -28, 6, 27, 18, -22, -26, -122, -86, -26, -125, 81, -123, -26, 39, -39, -48, 110, -64, 26, 124, -57, 28, -65, 111, 62, -19, -24, -56, 35, -123, -27, 50, -74, -6, 58, -18, -72, -126, -125, -2, 116, -89, 12, 71, -58, -26, 110, -50, -10, 77, -126, -39, 39, -125, 19, 111, -67, 74, -72, 102, -48, 75, -53, -52, 76, 18, 80, -3, 113, 13, -29, -35, -3, -58, 73, -27, -74, 38, -74, -71, -62, -59, 68, 58, -116, 26, -76, 53, -104, -113, 16, -95, -44, 72, -27, -40, 38, -23, -24, 40, -58, 120, -95, -115, 53, 82, 51, 42, 98, -61, -46, -42, 92, 68, 116, -23, 60, -123, 20, -117, 24, -64, -22, -82, -31, -74, -112, 29, -85, 79, -97, -66, -91, 34, -47, 0, -79, -36, -39, -4, 122, -90, 23, -110, -105, 93, 125, -104, 33, 22, 59, -110, 22, 118, -50, 92, -13, 77, -29, 29, -37, -71, 64, 49, 60, 123, -93, 20, 43, 109, 88, 112, 108, 50, 74, -48, -82, 19, 37, -78, 120, 34, -22, 85, -89, -32, 114, -59, 117, 122, 84, -21, -126, -92, 0, -67, -85, 86, -41, 11, -59, -77, 27, -127, -15, 47, -61, -107, 14, 0, -54, -73, 89, -107, -35, 78, -53, -39, 96, -1, 122, 2, 23, 84, 10, 28, -59, -96, 105, -6, 64, 71, -29, 73, 40, 113, 1, 13, 43, -25, 114, 11, -116, 119, 93, -13, 77, 110, -122, 2, -31, -92, 35, -59, -47, 38, -96, 1, 13, -70, 0, -122, 41, 114, -16, 49, 29, -117, -101, 82, -39, 105, -121, 52, 55, 97, 38, 98, 97, -24, 108, 12, 127, 47, -2, -58, -33, 26, 19, 69, 42, 101, -21, 63, -3, 94, -112, -122, -49, -90, 70, 52, -76, 78, 75, 79, 98, -8, 37, -13, 89, -27, -21, 111, -93, 36, -115, -105, 91, -45, -77, 113, -53, 47, -9, 103, 112, -26, -58, 71, 113, 95, -10, -90, -21, 11, -90, 104, -23, 44, -51, -82, -37, -71, -72, 65, -101, -16, -20, -44, -28, -92, -34, 116, -28, 47, 37, 31, 9, 106, 70, -89, -97, -37, 20, -9, -14, 107, 119, 88, -108, 75, -55, -113, -94, -6, 77, 24, 60, 16, 69, 53, 86, -72, -72, 12, 90, 93, 114, -52, 114, 63, 22, 100, -76, -117, -122, 58, -48, 103, -72, -14, 95, -41, -35, -90, 49, 22, -43, -104, 19, -54, -14, -60, -7, 35, 26, 82, -51, -121, -33, 121, 46, -50, -5, 13, 19, -54, -72, 104, -89, -43, -10, 72, 53, 41, 71, 3, -83, -11, -56, -123, -70, -112, 110, 107, 89, -39, -107, -5, -12, 66, 5, -28, 76, 30, 94, 43, -40, 78, 6, -107, 22, -76, -33, 62, 95, -55, 49, 115, -80, 38, -119, 127, -28, -84, -76, -75, 95, -119, -125, 45, 20, 118, 60, -54, -54, -65, -13, -47, 105, -117, 17, 106, 3, 38, 21, 102, -81, -69, 28, 7, 6, -128, -12, -44, -102, -114, 32, -17, 108, 81, 37, -127, 12, -24, -118, -64, 11, -1, -33, 125, 4, -105, -78, -69, -107, 85, -21, 9, 115, -30, -19, -73, -90, 18, -11, 122, 23, 54, 90, 41, 53, -78, -12, -32, -106, -89, -105, 51, 42, 30, -86, -87, 78, -121, 43, 52, 66, 119, -63, 64, 0, -101, 95, 64, -36, 91, 18, -36, -74, 19, 43, -61, 0, -113, 124, 77, -17, -119, -26, -80, -82, -3, 87, 51, -49, 60, 95, 10, 75, 24, -32, 50, -28, -4, 75, -113, -85, -126, -50, 104, 11, 94, -28, 112, 53, -63, 71, 28, 42, -37, 78, -62, 71, -31, -55, 52, -18, 90, -22, 18, 111, 66, -36, 6, -51, 64, -109, -25, 68, -65, 6, 56, -51, 97, -127, -59, 87, -59, -87, 23, -82, 38, -96, 48, -58, 126, 41, 11, 126, -51, -86, -29, -33, -26, 51, 64, 73, 6, -14, -69, 77, 39, 92, 111, 7, 81, 108, 1, 118, 5, -31, 95, 59, 98, -93, -42, 24, 59, 88, -21, 49, 77, 92, -117, 71, -88, 86, 80, -40, -54, 14, -119, 98, -24, -43, 62, -62, 45, 33, 14, 83, -19, 85, 15, 90, 119, -1, -22, 85, -89, 107, -51, -86, 65, -128, -48, -113, 54, 119, 113, 42, -1, 65, 52, -84, 0, 11, 99, -77, 66, -28, 95, 23, -118, -44, -50, -29, -121, 8, 122, 69, -37, 107, -67, 77, -1, 71, -17, 86, -4, -74, -51, -106, -16, -96, -52, 87, -97, -82, -57, 127, -49, 34, -86, 86, 43, 114, 50, 41, 79, 93, -106, 0, 1, -46, 85, 14, -114, 125, -8, -23, -28, -20, 74, -42, 67, 65, -116, -63, -61, 115, -126, 32, 57, 17, -19, -9, 81, -65, -44, -127, 73, 115, -112, -8, 90, -7, 81, 93, -42, -52, -101, 120, 28, 92, -74, -61, -126, 34, 58, -62, 74, 87, -105, 6, 105, -44, 44, -7, 64, -71, 47, -14, 77, 52, -39, -87, -8, 29, -70, -33, 90, -34, 82, 34, 1, 65, -126, -109, -57, -7, 56, -40, -72, 17, -33, -17, -127, -84, -27, -14, 61, 27, 97, 55, 38, -74, -101, 14, 108, 4, 73, 13, 44, -82, 4, 34, -33, 44, 94, 110, -24, -41, 119, 7, -75, 21, -12, -13, -57, -89, -86, 39, -26, 108, -11, -49, 11, 74, 36, -110, -128, 49, 30, -58, 20, -91, 4, 30, 65, -20, -77, 51, 41, -16, -107, 14, 9, -113, -42, 56, -12, -65, 32, -3, 26, -4, 70, 73, 75, -99, 73, -123, -77, -92, 5, -120, 96, 49, 113, 18, 46, 80, -91, -58, 81, 21, 81, 113, 15, 26, -30, -32, -77, 96, -19, 127, -58, 62, 94, 73, -5, 21, -30, 17, -12, 33, 100, -21, 72, 126, 49, 2, -111, -85, 38, -12, -23, 52, -85, 45, -38, 46, -15, 101, 11, -12, 100, -44, -59, 88, -18, 86, 51, -94, 71, 104, 90, 59, 71, -93, -28, 23, -16, -128, 3, -49, -123, -120, 26, -58, -128, -46, -94, 105, -99, -27, 13, 25, -33, 95, -58, 112, -100, -9, -36, 64, -61, -31, -56, 76, -17, -32, 19, 82, 127, -37, 117, 30, 53, -109, 64, -65, 46, 71, -75, 91, 76, -71, 5, -32, -116, -49, 121, 73, 109, 104, -78, 120, 96, 75, -12, 124, -124, -111, 118, 77, 118, -77, -36, 103, -19, 125, -119, 88, 11, 93, -113, -70, 116, -5, -116, -73, -80, 118, 29, -86, -97, 72, -101, -89, -103, 114, -105, -43, 3, -99, -11, 81, -40, 109, 23, 23, -108, -45, -116, -32, 31, -119, 116, -64, 20, 56, 67, -88, 72, 115, -7, 100, -31, -58, 105, -25, 14, -115, 25, 94, 81, -125, 121, -46, -5, 81, 67, -81, 13, -29, -37, 20, 119, -27, -20, -30, 46, -126, -85, 69, 91, 117, -37, -31, 51, 68, -98, 79, -121, -44, -110, 50, 88, -82, -25, 62, 49, -50, -44, 122, 36, 121, -45, -108, 102, -35, -3, -128, -89, 82, 28, 11, -9, -19, 115, 58, 56, 98, -9, 58, -24, -12, 20, 69, 69, 41, 89, 1, 22, 1, -87, 114, 12, -37, 116, -59, -78, 3, 66, 19, -61, -50, 51, -40, 34, 113, 5, -12, -94, -111, -91, -105, -122, -126, -75, 71, 102, 110, -39, 23, 8, -41, -105, 3, 58, -49, -53, -77, 9, 23, 45, -30, 11, -1, 42, -84, 87, 106, 126, -111, -123, 109, 38, -104, 12, 63, -52, 91, -41, 118, 22, -107, -120, 95, 104, -107, -65, 31, 59, -91, 108, 61, 94, 110, 74, -22, -127, -20, -81, 80, 77, -70, -66, 114, 10, 32, -82, -122, 85, -77, -42, -25, 121, -36, -56, 27, 117, -42, -57, 59, 117, -110, -15, -58, -69, -68, 125, -12, 105, -24, -72, -93, -55, -9, -75, -97, -114, 119, 29, 12, 34, 90, -98, -87, -37, 127, 42, -70, -126, -71, 49, 36, 21, -126, -126, -35, -125, -102, -52, -24, -103, -86, -25, 104, -52, -58, -112, -64, 111, 37, -88, -77, -77, 28, -109, 42, 114, 17, -7, 81, -9, -96, 94, -115, 6, -92, -9, 39, -62, -24, -3, -89, 70, -74, -48, 63, 5, 62, 39, 52, -72, 0, -6, 110, 57, -67, 70, 82, -41, 68, 120, 99, -32, -48, 78, 90, -2, -112, -76, 116, -92, 7, -81, -113, -47, 86, -7, -19, -15, 124, -33, 109, 59, -24, 38, -100, -94, -21, -37, 65, -104, -103, -59, 48, 94, 30, 18, 14, 92, 98, 115, -66, -20, 78, 78, 46, -23, -28, -18, 12, -126, -79, 30, -11, -101, 109, -101, 82, 26, 82, -57, -17, 71, 110, 4, -72, 109, -4, -78, -101, 59, -123, 103, -46, -71, -45, -15, 117, 126, -53, 4, 98, 10, -2, 45, -62, -55, 114, 34, -118, -90, -109, 114, 121, -38, 15, 61, -124, 122, 37, 81, -102, -71, -12, -53, 82, -115, 113, -8, 69, 21, 89, -47, -105, -75, -50, -51, -103, 14, -4, -38, -29, 11, -97, 101, 116, -26, -85, 45, 75, -122, -114, 10, 105, -12, -81, 35, 25, 106, 127, 77, -75, 98, 121, 24, 45, -50, 29, -87, -61, -65, -52, -103, 57, -75, 124, -87, -45, -92, -126, 7, -114, -64, 24, -107, 109, -69, -19, 28, -6, -42, 108, 100, -38, -48, -126, 120, 33, -88, 88, -7, -51, 99, -69, -118, 127, 1, -80, -58, 90, 11, 9, 95, -92, -85, -2, 61, 115, -14, 116, 31, 33, 22, 87, 34, -52, -21, 44, 75, -29, 28, -31, 121, -64, 18, 90, -100, 104, -90, 105, 32, -3, -71, -45, 21, -12, 5, -101, 53, -109, 47, 124, 124, 64, 13, -121, 80, 23, -117, -83, 26, 88, 70, 111, -121, -101, 45, -63, 87, -125, 14, 74, 56, -57, -27, -116, -107, -78, -24, 101, -3, -62, 69, 72, 67, -28, 26, -74, -113, 89, 45, -40, 4, 127, -68, 56, 0, 15, 92, 115, -88, 102, -94, 115, 88, 123, 17, 123, 123, 113, -124, 28, -104, 92, -67, 61, -128, 17, -86, 25, 17, 70, -38, 11, -12, 61, 87, -75, -88, -34, -102, 113, -72, -38, 33, -80, -103, -33, 122, -1, 101, 28, -110, 53, -101, 48, 70, 26, -86, -7, -78, 4, 96, -68, 105, -49, 89, -115, 126, 3, -30, -19, -19, 94, 73, -69, -2, -16, -122, 120, 69, -68, 19, 21, 46, 69, 50, 105, 76, -107, -127, -83, 104, 9, 79, -1, 0, -83, 104, 35, 117, 37, -114, -66, 117, -94, 68, 95, -88, -123, -119, -101, -79, -52, 0, -125, 3, 62, 18, -50, 27, 58, -61, -91, -25, -31, -73, -26, 100, -93, 29, -21, -67, 1, 77, 73, 112, 116, -113, -104, -15, -114, -41, -118, -52, -98, 7, -88, -1, -99, -64, -15, 126, -97, -76, 106, 66, 23, 86, 30, 54, 72, -62, -61, 65, 55, 26, 109, -5, -122, -92, -52, -43, 106, -8, -67, 15, 91, 90, -72, -92, 117, 49, -72, 3, 29, 27, -78, 22, 33, 90, 23, 49, 63, -62, 0, 11, 105, -90, 124, 20, -45, -82, 43, 65, -31, -65, -65, 122, -32, 33, 11, 22, 96, -120, 39, 72, 83, 120, 33, 92, -73, -115, 62, 105, -108, 11, -7, 19, -87, 10, 102, 17, -87, 6, 18, 122, -72, -112, 45, -50, 14, -124, 113, -81, 31, 12, 37, -113, 88, -46, -27, -103, 88, -14, 66, 48, -96, 49, 72, -37, -66, -115, 114, 82, -36, -78, -63, 124, 73, -4, 117, -6, 23, -58, -56, 54, 37, 60, 35, -108, 73, 46, 42, -89, 69, -18, 82, 96, -40, 123, -43, -118, -35, -109, 62, 126, 121, 7, 47, 38, 98, 114, -106, 4, -125, -14, 72, 119, 64, -49, -49, 39, -101, -106, 21, 54, 68, -58, 30, -35, 86, 105, 19, 72, 82, 69, -52, -106, -104, 123, 11, -119, -63, -74, -33, -109, 124, -78, -128, -99, -21, 60, 76, 13, 59, 74, -19, 81, -93, -2, -37, 118, -57, -15, 51, 28, -68, -110, 4, -59, 49, 79, 78, 82, 112, 54, 42, -50, -77, -85, 24, -10, -95, 80, -118, -111, 7, 92, -121, 12, -52, -7, 82, -54, 33, -117, -83, 2, -120, 102, 99, -18, 68, -15, -77, -47, 63, 26, 36, -66, -77, 82, -53, 103, 58, 92, -18, -84, -67, 94, 110, 115, 53, -4, 5, -58, 28, -92, 97, 109, -102, 78, -34, -111, -2, 86, 29, -64, -64, 116, 82, -58, 11, 34, -74, 88, -2, -86, 83, -128, -102, 97, -64, 27, -109, -89, -45, 64, 47, -62, 2, 70, -85, -17, -59, 88, 65, -3, -26, -5, 19, -116, -11, -65, -15, -95, 119, 97, 0, -125, -84, 56, 104, -30, -111, 114, -122, 58, -42, 8, 53, 0, 88, 51, -119, 55, 115, 109, 28, 9, 124, 125, -77, -113, -43, 88, -2, 15, 12, 80, -81, 36, 11, -107, 117, 89, -126, -80, 18, 103, -3, 16, -79, 51, -124, 13, -1, -84, -3, -36, -123, 115, -34, -60, 67, -76, 35, 39, 37, 37, 95, 25, 119, 119, -67, 28, 52, 7, 55, -62, 17, -90, 112, 49, -30, 84, -71, -74, -9, -30, -57, 109, 82, 74, -114, -91, -30, -14, -30, 38, 39, -112, -101, 9, 10, 78, -49, 51, 126, 121, 55, -28, -81, 36, -78, 53, 14, -54, -110, -127, 47, -3, 10, 57, 121, -15, 16, -93, 64, -75, 68, -31, 29, -44, -117, -96, -33, 36, -98, 7, 39, -88, 75, 49, 73, -125, -69, -67, -73, 60, -30, 98, 65, 29, -113, -24, 12, -24, 90, 89, -84, 117, 113, 70, 124, -71, 65, -99, -71, 0, 32, 27, 20, 53, 25, 125, -19, -105, -61, 60, -82, 77, -93, -98, 89, 24, 39, -121, -101, -44, -18, 48, 27, -116, -116, 43, 67, 57, 79, 48, 32, 32, -44, -61, 2, 68, -71, -110, 9, -89, -68, -115, 15, -4, -86, 99, -72, -99, -71, 88, -16, 126, 70, -127, 43, -29, 114, 106, 12, -82, 103, 38, 9, -85, 119, 9, -64, 58, 64, 20, 99, -89, 123, 41, -121, 64, -64, 57, 108, -69, 24, -29, 14, 74, 34, -96, 21, -17, -12, -84, -51, 35, -107, -90, -12, 20, -81, -120, 117, 68, 91, 7, 60, 89, -32, -111, 16, -8, 51, 29, -110, -52, -121, 39, 95, -29, 9, -45, -82, 64, -34, 3, 41, -94, -69, -72, 76, -120, -54, -28, 90, 24, 100, -52, 27, 5, -36, -97, 6, 47, -68, 62, -19, 68, -69, -75, 108, -61, -56, 57, -82, -35, 27, -54, 109, 118, -82, 41, -68, -127, 54, -68, 87, -43, 46, -7, -7, -74, 106, -124, -28, 20, -88, 0, -54, -59, -60, 7, -4, -107, -109, -125, 21, 34, -26, 82, -116, -91, -74, -76, 41, 117, 23, -20, 85, -121, -69, -74, 31, -42, -45, 2, -101, 12, -58, -24, -104, 117, -27, 112, -54, -21, 92, -110, 41, 40, -3, -20, 111, -26, 57, 52, 43, -98, -83, 95, -16, 95, 9, -48, -77, -125, 39, -104, 26, -43, 53, -94, -35, -32, 82, 107, 20, 80, -99, 91, -92, -114, -100, 43, 9, 9, 5, 46, 60, -58, -50, -58, 3, 37, -10, -16, -13, 79, 90, 91, -70, -124, 31, 116, 115, 111, -50, 80, -29, 89, 39, 8, -72, 54, -59, 37, -128, -2, 40, -95, 61, 41, -17, -112, 64, -113, -54, -13, -109, -50, 0, -77, -98, -60, -100, 10, -5, -53, 103, 15, -128, -93, 64, 32, 52, -11, 57, 69, 11, -36, -48, -82, -104, 32, 44, -31, 24, 56, 2, -118, 86, 13, -123, 119, 100, 33, 77, 117, 91, 78, -84, 126, -82, 2, -38, -17, -8, -76, -89, -35, -91, 104, -38, 8, 112, 57, 46, -80, -15, -45, 113, -28, 3, -88, -20, -68, -64, -77, -44, 28, 77, 34, 57, 28, -78, 71, 91, 102, 88, -125, 8, -71, -81, 91, 104, -102, -59, 96, 112, -24, -114, 92, -2, 0, -116, -86, 104, 49, -64, -48, 19, 22, -56, -8, 40, 125, 38, 80, -1, -101, 97, -119, 76, 96, 60, -50, -37, -57, 86, 106, -85, -76, 16, -97, 29, -13, 61, 22, -32, -120, -51, 20, 88, -13, 109, 7, 47, 106, -82, 64, -18, 67, -102, 44, 78, 113, 33, 22, -121, 109, 86, -42, -128, -5, -23, -54, 106, 97, -11, -33, 45, 13, -48, 92, -111, -43, 11, -9, -65, 84, -8, 116, 52, -66, 14, 48, -114, 103, -43, -7, -97, 83, -71, -21, -33, -53, 100, 18, 76, 124, -84, -109, -99, 66, -37, -80, -112, -125, -115, 46, 92, -35, 119, -29, 100, 83, 20, 123, -22, 0, 81, 115, -82, -45, 65, 105, -53, -31, -94, -44, 49, -40, -125, -62, 37, -33, -51, 17, 33, -108, -28, 103, -70, -14, 25, -40, 80, 100, -31, -105, -116, -13, 54, -23, 88, 93, 1, 7, -14, 61, 28, 39, -93, -39, 85, 122, -84, -101, 53, -5, 22, -27, -84, 64, -6, -116, -46, -100, 124, -87, -88, 13, -81, 60, -71, 30, 56, 85, -50, 67, 36, 0, -30, -48, 13, -30, -47, 27, 4, -25, -37, -105, -115, -12, 108, -121, -26, -53, 28, 69, -65, -72, 54, 2, 6, -122, 72, 64, -93, 127, 107, -51, -85, -79, 102, -102, -33, -55, 110, 101, 49, 84, 112, 19, -95, 70, -128, 66, -2, -39, 50, -3, -120, 99, 125, -30, 12, 119, 7, -78, 14, -66, -48, -41, 21, -2, -95, 82, 116, -48, -29, -108, -122, -21, 77, -16, -8, 45, -37, -30, -102, 27, -46, -9, -72, -36, -126, 107, 39, 45, 37, 94, -29, -122, 106, 65, 109, -112, 58, -4, 2, 60, -68, -122, -45, 7, 14, -80, 58, -108, -68, -36, -39, 124, -107, 61, -126, 71, -94, 108, -121, -52, -30, -77, 126, 61, -54, -60, -54, -81, 96, 61, -53, -115, -122, 94, 126, -8, 72, 60, 117, -119, -77, 16, 76, -38, -79, 22, 111, 119, 3, -62, 60, -76, 21, -85, 121, -103, 23, 26, -54, 7, -4, -30, -45, 127, -42, -90, 113, 22, -105, 82, -118, 105, -43, 102, 89, -1, -4, 11, 89, -27, 117, 77, 70, -123, -94, -88, 62, -108, -14, 119, 115, -5, -22, 14, -85, 31, 3, 111, -32, 120, -37, -127, 14, -16, -44, 120, 8, -21, -2, -108, 90, -124, -41, -93, -79, -82, -124, -92, 56, -87, -109, 32, 79, -54, 112, 59, -41, -97, -128, 20, 118, -54, -72, 8, -63, 64, 29, 120, -34, 110, -74, -4, 39, 91, -78, 42, -9, 74, -95, 64, -93, -9, -104, -10, 64, 28, 77, 28, 62, -15, -15, -59, 18, 16, -127, -119, 77, 102, -45, 110, -89, -102, -83, 103, -85, -52, 42, 90, 48, -89, -68, 54, -3, -108, 53, -121, 105, 124, 94, 37, -98, -84, -53, 71, 26, 114, -85, -69, 124, 23, -105, -31, 25, -67, -113, 15, 52, -45, 63, 58, 45, 84, -102, -90, -26, -19, 3, -24, -119, -25, 86, 36, 80, 113, -84, -64, -125, -81, 6, -111, -8, 7, -23, -40, 15, -53, -106, -82, 114, -83, -27, -15, 60, -75, 41, -117, -78, 12, -115, 44, 95, 41, -118, 79, -23, 1, -54, -52, -92, -45, -28, -10, -82, 60, -83, 43, 16, -80, -68, -66, 73, 103, -65, 116, 17, -95, 8, 91, 51, -36, -19, -38, -86, 33, 96, 109, -116, 9, -85, -35, -70, -38, -24, 98, -101, -15, 63, 100, -127, -128, -51, 62, 16, -40, -13, 55, 24, 72, 112, -118, 116, 101, -69, 65, 86, -24, -37, -36, 52, 118, 28, -37, -10, 51, 38, -104, -51, 61, 115, 104, 51, 0, -70, 48, -108, 64, -73, 31, -39, 89, -102, -74, 54, -15, 61, -50, 38, 57, -10, -54, 124, 101, 92, -52, -5, 101, 26, -90, -94, -16, 12, -121, 52, -118, 125, 115, -37, 33, 92, -49, 8, 13, 109, -82, 92, 48, 84, 2, -1, 101, 72, 0, -92, -115, 85, -116, 11, 56, 27, 19, 124, 57, -64, -117, 69, -73, 23, 121, -113, 53, 37, -87, 118, -97, 43, -113, -41, -2, -37, 116, 64, -80, 93, -101, 29, 16, -3, -68, -3, 90, 113, -56, -74, -102, 45, 113, 98, -111, -88, -78, 63, -51, 83, -22, 72, -121, -109, 33, -30, 95, 20, -66, -30, 108, 89, 43, 52, -95, -111, -118, 87, -1, -19, 107, 74, 108, 70, -6, 10, 107, 49, 124, -36, 28, -67, -89, 76, -123, 60, 53, -23, -104, -125, 77, -16, 19, -49, -69, -56, -8, 78, 70, 5, -60, -30, 101, 90, 108, 32, -108, 123, -72, 121, -109, -35, -7, 14, -126, 99, 26, -67, -73, 5, -18, 123, 71, -73, 73, -84, -90, -56, 73, -106, 96, -89, 80, -122, 64, -115, 13, 52, -100, -49, 37, 28, 22, -27, -4, 119, 57, -102, -105, 69, 101, 55, 39, -60, -35, -25, -111, -69, -121, -41, 88, -35, -83, 98, -13, -40, -46, -46, 111, 43, -2, 85, 59, -101, 62, 105, -74, -1, 96, 6, -124, -98, 30, 114, 65, 67, 122, 114, 11, -64, -98, 73, 76, 97, -24, -12, 69, 125, 50, 111, 6, 44, -75, -9, 73, -12, 41, -95, -124, 45, -93, -23, 27, 47, 86, -6, 78, -73, -30, -3, -27, -119, -96, -53, 41, 67, 86, -72, 75, -103, 117, -22, -95, -71, -2, -40, 65, 67, 67, -18, -83, 70, 123, -8, -83, 25, 90, -95, -94, -37, -110, -85, -110, 94, 28, -47, 45, -69, 98, -33, 9, 53, -3, 84, -31, -29, -92, 38, 49, 88, -121, 78, 66, -91, 107, -125, -106, 97, -37, 63, 42, 44, -21, -27, 103, -76, -61, 95, -45, -108, -25, 7, -18, -30, 17, -86, -36, 13, -112, -21, -98, -112, -49, 35, 37, 82, -16, 93, 123, 84, -90, -125, -124, 24, 76, -35, 99, 108, -24, -59, 121, -97, 0, -41, 101, 104, -100, -19, -45, -79, 123, 25, 39, -120, -91, 121, -62, 46, -61, -57, -32, -96, -28, -125, 20, -91, -94, 74, -64, -107, -76, -108, 118, 60, -101, -36, 36, 40, 73, 50, -92, 68, -22, 15, 124, -13, 32, -113, 82, -16, -72, -21, 87, -4, 91, 127, 38, -84, -116, -111, 62, -77, 62, -79, -110, 40, -48, 0, 20, 106, 40, 5, 97, 127, 53, -17, 96, -7, 70, 27, 65, 28, 37, -122, -58, 13, 72, 118, 58, 106, -31, -97, 122, 44, 57, -93, 54, -35, -19, 70, 100, -76, -18, 33, 15, 73, 53, -109, 71, -110, -26, 30, 38, 57, -39, -44, 68, 17, 39, 117, 118, 1, 84, 37, 120, 40, -3, 96, 2, 6, 122, 7, -115, 122, 76, 82, -77, -18, 94, 127, 67, -28, -89, -126, -121, 40, 61, 21, 39, -72, 12, 99, -39, -81, 98, 70, -20, -86, 96, -88, -57, -96, -51, -38, 107, -17, 38, -60, -57, -44, -80, 45, -88, -88, 17, -119, 61, 79, -56, -108, -80, 18, 82, 61, -124, -37, -124, -75, 73, -30, 51, 106, 124, -120, 44, -88, 97, -20, 117, 75, -93, 91, -94, 80, 3, -92, 75, -1, 82, -31, 1, 93, 69, -4, 76, 47, -109, 90, 87, 52, -128, -93, -86, -36, 41, -56, 30, 23, -44, 12, 20, 120, 11, -60, 75, -95, 64, -90, 16, 73, 14, 12, 21, 126, 100, -119, 83, 56, 81, 6, 42, 72, -97, 78, 75, -50, -58, 29, 44, -51, -98, -52, 39, -58, -24, -71, -3, -21, -79, -109, 55, 26, 124, 108, -100, 11, -111, -45, 109, 73, 8, -44, -63, -24, 55, -64, -119, -55, 90, 122, -122, 125, -6, -86, -67, -67, -23, -20, -1, 122, 91, 108, 122, -73, -53, -69, 99, -59, 42, -1, 13, -57, 59, -95, 11, 91, 8, 48, -45, 30, 73, 10, -37, 37, -63, -32, 3, -52, -43, -88, 85, -114, -86, 36, -90, -127, 35, -49, -51, -56, -41, 120, -18, -62, -53, -69, 55, 72, -106, 18, 104, 127, -44, 27, 30, -1, -99, 72, 83, 91, 27, 15, -119, 77, -128, -105, 95, -67, 31, -69, -47, 1, -19, -28, -23, 90, 120, -103, -95, -90, -120, -22, 13, -6, 61, -47, 115, -84, -64, 39, -86, 118, 115, 77, 111, -71, -26, -83, 63, 35, 8, 81, -98, -81, -91, -23, 23, -123, -87, 76, -11, -122, -9, 42, 9, -22, 23, -86, 26, 86, 52, 2, 28, 108, -87, 25, -121, 23, -89, -99, -101, -82, 101, -92, -78, -15, -107, -59, 109, 98, -123, -37, 86, 83, 124, 56, 90, -77, -34, 83, -23, -54, -124, -56, -38, -102, 90, 127, 6, 118, 73, 102, -85, 44, -23, -38, 121, 127, 106, 92, 101, -61, 40, -87, 113, 71, -56, -104, 19, -105, 32, -57, -70, 83, -114, 58, -85, -112, 16, 38, 123, -75, 7, 115, -44, -89, 118, -96, -54, -97, -100, 104, -11, -122, 121, -120, 53, 57, -102, -49, -11, 22, -4, -19, -34, -38, 109, -60, 57, -92, -76, -70, -116, -89, 127, 30, -65, -11, -97, -111, -97, 25, 13, -41, 63, 1, 62, 20, -117, -3, 75, -108, -19, 103, 57, -50, -99, 5, -54, 24, -37, 63, -125, 13, -62, -80, -82, 96, -18, -115, -80, 57, -46, 23, 124, 52, 41, 89, 60, 74, -97, -76, 108, 94, -27, -42, -10, -98, 45, -118, -27, -17, -11, 102, -22, -124, 124, -83, -106, 14, 104, 104, -21, -110, -111, -57, 78, 34, 45, -71, -87, 75, -100, 104, 82, 84, -4, 127, 96, 45, 31, 51, -87, 67, -91, 20, -59, 15, 85, 56, -79, -90, -49, 109, -123, -65, -124, 117, 107, -35, -13, -34, 58, -42, -17, 122, 17, 16, -7, 19, 11, 123, 115, 5, -54, 49, -99, 31, 117, 119, -8, 55, 76, -53, -112, 91, -104, 112, 25, 82, -128, -74, -61, -41, 12, 75, -13, 49, -59, 113, 22, 125, -15, 119, -39, 108, -19, -126, 126, -29, -105, 77, -75, -80, 54, -7, 58, -62, -84, 25, -69, 58, 1, 100, 30, -46, 4, -34, 112, 111, 8, 9, 61, -61, -15, -64, 15, 33, 120, -25, 81, -36, 126, -52, -39, 112, 22, 88, 102, 107, 52, -96, 62, 124, -97, 79, -96, 95, -68, 1, 112, -83, 98, -11, 63, -49, -32, 72, -75, -115, -109, -45, 126, 73, 28, -102, 30, 89, 32, 91, -81, -86, 34, 29, 111, 19, -107, 109, 90, -66, 126, 68, 43, 38, 42, 95, 79, 90, 90, -13, -120, 119, 13, 35, -61, -11, -5, 36, -99, -98, -33, -99, -55, -62, 61, -59, -45, 86, -67, -29, 6, 28, 124, 14, -44, 6, -46, 41, 116, 109, 99, 49, -120, -72, -14, 31, -78, -10, 35, -94, 106, 69, -126, 14, -28, 26, 36, -62, -119, 66, -68, -92, -48, -9, -50, -24, -116, -47, 121, 3, -81, -69, -62, 63, 67, -36, 117, -41, 126, 37, 78, -10, 55, -36, -106, -40, -54, -69, -124, 1, 44, 112, 3, -59, -126, 73, -43, -121, 82, 62, 125, -37, -8, 14, 118, 43, -29, -56, -117, 79, 56, 54, 83, 10, -14, 100, -8, -98, -8, 116, 91, 101, -33, 42, 127, -88, -87, -106, 65, -34, 61, -91, 6, -106, -109, -21, -50, -106, -37, 94, -10, 38, -93, -66, 49, 50, 124, 103, 52, 37, -114, -73, 24, -96, -7, -121, 103, 62, -55, 54, -77, 75, 61, -18, -63, 80, -63, -32, 16, 58, -48, -57, -49, 2, 46, 28, 11, -75, 122, 20, -55, 67, 7, 116, 119, -43, 113, 119, 72, 95, -87, -34, 42, -39, 63, 23, -18, 27, -38, -78, 43, 99, -89, -68, -16, -104, 27, 109, 118, 106, 71, 70, 30, -19, -124, -78, -79, -76, -55, 2, -78, 36, -12, -101, 83, 17, -44, -110, 73, 61, -34, -127, 78, -40, 83, 18, 49, -36, -85, -110, -33, 27, 101, 89, 60, -110, -121, 8, 2, 41, -19, 123, 124, 114, -39, 18, 88, 53, -29, -69, -32, 8, -5, 19, -74, 48, 11, 126, 71, -116, -23, -72, 87, 22, 48, -4, -102, -109, 123, -49, -76, 89, -108, 51, -78, 70, 25, 39, -109, 65, -104, -69, 88, 0, -50, 90, 15, 84, -99, 49, -106, -20, -117, 100, 100, -49, 50, -119, 108, -36, 31, 49, -105, 24, -48, -68, 123, 83, -28, 114, -44, -77, -13, 119, 17, -32, -82, 35, -124, -11, 93, -27, 111, 121, 23, -5, -15, 56, -74, 34, 120, -66, -38, 44, -124, 18, -100, -83, -107, 56, 89, 101, 2, 87, 16, 53, 53, -89, 37, -81, -14, -114, 120, 16, -121, 9, -34, -123, 52, 53, -105, -30, 32, -114, -42, -19, 121, 59, -94, 123, 58, -106, 67, -34, -30, 69, 52, -19, -75, 85, -95, -66, -96, 75, -79, -23, -15, 57, -20, -65, -65, -60, 113, -88, -66, 12, 123, 68, -31, 4, -23, 82, 102, 112, 65, 84, 109, 101, -75, -95, -28, 127, 56, -112, 2, -113, 89, -100, 70, 58, -76, -41, 68, -78, 56, -82, -29, 15, 12, 78, 101, 2, -57, -88, 5, 116, -63, -58, 126, -106, -127, 53, -91, -107, 37, -125, -112, -111, 48, 103, 48, 48, -90, -2, -8, -21, -87, -14, 13, -50, -90, -95, -126, -28, -28, -47, 43, -113, 108, -49, 76, -43, 94, 21, 104, 25, 60, -104, -23, 50, 36, 116, 45, -2, -92, -78, 127, -25, 65, 36, -13, -112, 32, -20, 59, 47, -33, 35, 28, 54, 81, -102, -10, 64, -14, 38, -27, -36, 40, -41, -32, -78, -6, 119, -97, -90, 97, 60, -96, -7, 114, -121, -8, -89, 85, 81, -104, -71, -85, -57, 18, -62, -25, -69, -116, -104, -73, -34, -11, -45, -56, -33, 68, -10, 63, 24, -40, 120, -68, -57, -45, -15, -63, -58, -69, -8, -107, 24, 63, -79, 47, 30, -101, -36, 83, 88, -35, 61, 29, -49, 111, 39, 51, 75, -59, -113, 111, -88, -81, 53, 24, 35, -94, -71, -72, 12, 48, -104, -67, -113, 17, -18, 14, 26, -115, -117, -10, -63, -78, 82, -89, -4, 76, 104, -16, 39, -51, -86, 37, -6, 117, -88, -56, -61, 110, -25, 6, 0, -124, 124, -40, -84, -52, -110, 63, 18, 47, -58, 95, -119, 118, 62, 91, -53, -107, -13, 56, 8, 110, -123, -16, 54, -84, -36, -37, 9, -57, 84, -23, 40, -25, -26, 37, -91, -120, -99, -46, -22, -21, 108, 45, -84, 119, 36, 89, -62, 1, 116, -91, -102, -22, -39, 4, 10, -48, 37, 86, 100, 13, 25, 95, -62, -99, 18, -119, 6, -68, 4, -88, 40, 106, -44, -35, -105, 21, -55, 7, -119, -70, 108, -43, 110, 75, -65, -70, 127, -97, 115, -69, 124, 107, -105, -33, -60, -45, 102, 7, 119, -11, -2, 102, 65, -16, 8, 112, 61, -2, -1, 64, 56, 91, 36, 70, 123, -48, 76, 12, -113, 43, -6, 27, -16, 56, 122, -16, -27, 116, 54, -12, -124, -26, 112, 17, 105, -58, 40, -41, -105, -128, -80, 27, 111, -28, -79, -109, -92, -31, -73, 81, 11, -30, 63, 111, -94, -4, -64, -48, 78, 36, 45, 64, 52, 119, -74, -16, -117, -85, -55, 113, 49, -21, 37, 57, 96, -30, -50, 9, -40, 65, -103, -94, -42, 48, -2, -67, 52, -21, -105, 64, 12, -40, 22, -122, -61, 33, 87, 99, -101, 94, -4, 22, -2, 2, -20, 59, -88, 34, -51, 6, -94, -114, -100, -21, 75, -86, 91, -60, -112, -113, -45, -29, -94, -38, 45, 113, -13, -30, 38, 1, 31, -84, -53, 42, -101, 78, -4, -2, 98, -105, 60, -50, -73, 69, 117, -51, 116, 76, -70, 59, 90, -115, -1, 20, -65, -38, -10, -128, 31, -16, -20, 41, -17, 58, 88, 119, 3, -119, -106, 83, -109, 127, 92, 24, -24, 110, 42, -114, 15, -54, -77, 43, 72, -55, 126, -64, 5, 15, 104, 61, -62, 115, 127, -93, -83, -116, 79, -127, 40, 7, 69, 79, 60, -59, -83, 14, -127, 68, 30, -64, 45, -40, -22, 34, 14, -44, -7, 107, -89, 100, 13, 72, -20, -123, 49, 102, -69, 116, -34, -110, -77, 105, 89, 101, -98, -16, 43, -94, 57, -75, 31, -77, 8, -70, 65, 72, -29, -37, 99, 29, 5, 4, 65, 112, 34, 46, 122, 94, -94, -56, 72, 75, -29, -24, 94, -57, 36, -78, 93, -21, 45, 84, -31, -40, -86, -117, -101, -64, -10, 14, -122, 103, 11, 70, 99, -75, 87, -126, -41, -17, -55, -15, -76, 91, 82, -60, -49, -42, 61, -46, 115, -57, -52, -51, 62, 45, -10, -28, -58, -78, -7, 88, -41, 101, -37, 16, 61, 54, -9, 103, -101, -36, 127, 126, 105, -52, 4, -119, 62, -73, -92, 55, 81, -58, 13, -119, 102, -33, 75, -26, -108, -18, 7, 74, -69, 102, 18, -96, 103, -102, 66, 30, -24, -55, 121, -115, -50, 43, -76, -79, -89, 18, 123, -72, -64, -119, 38, -71, 110, -102, 58, 108, -73, -40, -72, -74, -17, -34, -7, 82, -52, -89, -89, 109, 124, -52, 60, -7, 49, -17, 60, 107, 40, 9, 46, 57, -118, -112, 52, 89, -108, 96, -48, -15, 83, -92, -82, -31, -49, 106, 60, 114, -71, -83, 102, 46, 13, 82, 78, 15, 13, -122, -66, -88, -103, 9, 95, -21, -86, 85, -77, 83, -123, -36, 116, 60, -57, -118, -68, -37, -52, -70, -110, -112, 12, -95, -55, 97, -75, 105, -124, 103, 96, -43, 63, 38, -110, 15, -39, -33, 40, 10, -116, -81, 20, -68, 73, 23, -32, 83, 122, -56, 30, -108, 38, -103, -7, 34, 97, 53, -83, -4, -43, 50, 92, 104, 17, 106, -26, 52, -115, 81, 79, 87, 105, 59, 62, 110, 30, -104, 42, 124, -18, -86, 56, 125, -16, -52, -78, -128, 6, 16, 44, -74, -47, 20, -22, -1, 49, -53, -120, 63, 47, -12, 40, -107, -98, 90, -74, 20, -24, 91, -41, 88, 109, 77, -76, -48, 43, -35, 61, -68, 124, 18, -71, -118, 44, 111, 19, 40, -41, 117, 40, 8, -43, -104, 120, 26, -34, 103, 112, 42, -60, 86, 88, 14, -4, -84, 118, 40, -24, -66, -2, -47, -23, -44, 111, 86, 75, 111, -39, 32, 70, -62, 2, -4, 17, -59, 35, -79, -64, 41, 99, 124, 61, -102, -71, -76, 29, 90, -30, 59, 18, -39, -89, -67, -79, -116, -16, -76, 74, -51, 97, -70, -98, -10, 50, 95, 69, -128, -80, 94, 28, -78, -47, -18, -73, 124, 117, -96, -48, 100, 59, 46, 30, -11, -87, 63, -48, 125, -97, -46, -38, -38, -79, -111, -115, 25, 125, 60, -20, -39, -106, 84, 65, 47, 127, -13, -23, 6, 72, 108, 96, 25, -128, -98, 42, 30, -82, -25, -95, 55, 88, -6, 15, -80, 42, 25, -87, 81, 63, -85, 5, 56, -44, 4, -74, -116, 114, -36, -101, -39, -66, 63, -126, 23, 13, -45, 96, -2, -114, 50, -90, 98, -24, 71, -19, -110, -33, -32, -60, 125, -102, 123, -20, -79, 118, -10, 1, -109, -119, 109, 43, -16, -56, -10, -69, -38, -71, -34, -126, -111, -53, -43, 26, 1, -69, 115, -40, -108, -11, 63, 14, -24, -100, 84, 29, -120, 37, 35, -38, -67, 124, 49, 76, 31, 78, 57, -44, 73, 0, -94, -28, 9, -86, -91, 74, 79, -120, -108, -102, -69, 64, 3, -104, 92, -70, -59, -109, 76, -32, -87, -30, 67, -31, 86, -105, 5, -21, -112, 104, 74, -111, 5, 121, 3, -4, -13, 30, 7, -12, -65, 4, -107, -104, -98, 107, 55, -69, -96, 49, 83, -12, 69, 45, 112, 1, -49, -48, -39, -13, -77, 57, -85, 81, -12, -36, 97, -124, 85, 90, 98, -128, -23, 95, 107, 46, 28, 123, -98, -72, -64, -40, 7, -50, 41, -122, -99, 87, 126, -125, -4, 2, 66, 14, 56, 19, 53, -31, 55, -98, 13, 100, -69, 85, 0, 14, 116, -50, -13, 72, 11, 43, 90, -90, 84, -115, -49, -83, -89, -1, 111, 86, 73, 117, 53, 92, 77, 46, -51, -74, -125, 4, -38, 93, 56, -47, -80, -5, 77, 91, -81, -119, 59, 56, -41, -26, -108, 55, -58, 57, 20, 119, -32, -95, -118, -48, -102, -97, 45, 65, -110, 20, 80, 107, 47, -77, 16, 18, -70, -102, 23, -19, -99, -32, 115, 90, -72, -84, 24, 73, 43, -98, 41, 77, -1, 52, 66, 42, 0, 85, -40, -108, 16, -5, -1, 17, -65, 65, 97, 95, -30, -20, -13, 38, -65, -29, -39, 61, -45, 43, 2, 97, -62, 112, -64, 118, 107, 16, -79, 1, 41, 39, 20, 7, 103, -44, 115, -43, 36, -118, 38, -66, 32, -73, -38, -18, 69, -23, 28, -38, 91, 67, -32, -95, 48, -7, 18, 93, 40, -14, -13, -108, -21, 53, 57, -23, -123, -44, 73, 60, -13, -83, 47, 51, -96, 89, 50, -106, -40, -86, -98, 116, 107, -56, 35, -7, 91, 24, 10, -25, -29, 57, 55, 105, 90, 32, 72, -70, -83, 13, -59, 120, 121, 66, -10, -64, 79, 79, 28, -44, -108, -28, -30, -31, 98, -48, -21, -26, -35, 37, 76, -98, -111, 36, -11, -14, 78, -38, 93, 77, 92, -120, -24, -101, -123, 29, 44, 77, -57, -43, -26, -97, -81, -54, -67, -31, 85, 9, -18, -74, -58, -73, -77, -127, 89, 8, -99, -66, -86, -21, -85, -100, 5, -109, 13, -50, -9, 99, -27, 125, 58, 71, 66, -20, 109, -103, -85, 67, -7, -110, -46, 18, -44, -88, -115, -104, -12, -11, 85, 6, -7, -2, 78, -118, -102, -47, 22, -85, -39, 117, 10, 12, -97, 71, 123, 111, 4, -91, -30, -14, 50, 14, 12, -83, 8, -69, -115, 14, 119, -23, -128, 97, 6, -40, -6, -59, -126, 70, 82, 119, -38, -64, 20, 31, -42, 73, -44, -96, 98, 60, -85, -39, -24, -33, 26, -43, -54, 111, 122, 35, -86, 58, 123, -98, 56, 12, -98, 127, 115, -115, 72, 7, -121, 50, -46, -25, -30, 30, 76, 117, 48, -60, 74, 2, -97, -71, -60, -47, 41, 46, 97, 71, -67, -102, 101, 112, 71, 53, -2, 60, 91, -18, -79, 36, 31, -17, 39, -48, -91, -15, -91, -90, -107, 87, 126, 45, 13, -112, -72, -78, -40, 43, 8, -77, -81, 11, -89, 99, 23, -106, 77, 89, 120, -122, 1, 104, 75, 1, -6, 70, 39, -83, 79, 42, -62, -86, -47, 120, -67, 115, -22, 83, -124, 53, 91, 31, -62, -74, -4, -10, -90, 0, -76, 15, -35, 87, 11, 74, -67, -16, 127, -80, -57, -69, -99, 5, 15, -123, -45, 40, 105, 10, -13, 114, 117, 24, 37, 2, 111, 107, 102, -52, 51, -23, 34, 6, -90, -54, -96, -16, 104, -66, -22, 70, -125, 104, 62, 94, -5, 0, 70, -71, 104, -122, -66, -101, 50, -114, -54, 23, 86, 124, 45, -28, 44, -60, -87, 60, -61, -44, 43, -80, -60, 49, 11, -59, -21, -6, 79, 24, 29, -82, -32, -35, 87, 36, -82, -86, 4, 77, 82, -93, 35, -13, 71, -63, -35, 53, 36, -80, -125, -8, -84, -126, -81, 45, -100, 30, 58, 67, 72, -105, -54, 126, 54, 56, 4, 69, -16, -14, 4, -126, -68, -58, -25, -23, 65, 34, 79, 123, -75, -111, 7, -106, 57, 124, -26, -62, 124, -126, 10, -69, 13, -18, -22, 73, 66, -99, -86, 54, -9, 50, 118, 50, 114, 123, -32, 68, 2, 36, 38, 60, 79, 75, 75, -17, 115, -57, -65, 93, 109, -80, -75, 127, 86, 67, -20, -91, 72, -82, 24, -95, 105, 109, 25, -19, 111, 87, 82, 90, 117, 49, 58, 29, -59, 100, 5, -63, -122, -115, 1, 74, 17, -23, -118, -4, -93, -12, -18, 13, 116, -91, 14, -3, 100, 2, -90, -20, 79, 32, 35, 10, 110, 63, -94, 77, 63, 127, -20, 122, 70, -96, 43, 105, -3, -115, 116, -78, 120, -123, 109, -126, -111, 13, -49, -35, -70, 19, -13, 70, -49, -17, 61, -112, 42, 24, 4, 21, -28, 26, -77, -31, -104, 73, -1, -58, -49, 30, 125, -87, -69, -109, -83, 112, 48, 10, 64, 79, -62, -25, -5, -37, 0, 11, -25, -40, 47, 11, -24, -115, 48, 82, -112, 16, -48, -42, 18, 9, -74, -53, -20, -107, -43, 85, -58, 29, -85, 20, -121, -78, -90, -92, 47, 21, 34, -113, -68, -59, 103, 5, 30, -50, 61, -89, -39, 5, 118, 86, -43, 97, 9, -47, -41, -124, 81, -16, 79, 53, 43, 9, 113, -81, -55, -28, 66, 31, -82, 105, -2, 117, 21, -70, -113, 20, 11, 17, 88, 88, 37, -71, -122, 109, 15, -57, 99, 122, -65, -109, 18, -109, 90, -1, -94, -69, -37, 25, -113, 125, 11, -6, -125, 29, -124, -83, -30, -56, -89, 10, -10, 37, 112, 80, 1, -11, 4, 35, 80, 68, -82, -7, 87, 21, 57, -17, 71, 18, 103, -118, -109, -19, 5, 13, -119, -46, -40, 38, 1, -101, -37, 22, 19, 94, -29, -16, -68, 23, 76, -119, -46, -34, 1, 113, -26, -13, -79, -35, 19, -25, 81, -69, -123, -49, -7, -59, -111, -43, 49, -47, -88, 67, -100, 43, -86, -59, -5, 33, 92, 22, 9, -92, -46, -113, -12, 51, 61, 115, -41, 19, 15, 70, -12, -104, -35, 66, 79, -67, 24, 54, 72, -93, -16, -34, 57, 89, -120, -88, -60, 80, 36, 78, -89, 5, 51, 9, -50, -3, -18, -17, 8, -66, 23, 60, 126, -49, -53, -33, -89, -17, -53, 37, 94, -81, 2, 0, 25, 69, 75, -121, -18, 68, 88, 7, 37, -36, -107, 39, 102, 47, -103, -122, 15, 34, -58, -110, -103, -49, 94, -69, 48, -9, 26, 4, 127, 35, -53, -113, 114, -21, 15, 101, 69, 45, -127, -53, 122, -10, 38, -17, -79, 106, -80, 4, -52, -86, 45, -52, -10, 89, -37, 98, -70, 123, -57, -56, 116, 0, -66, -27, -69, 89, -128, 25, -106, -51, 52, -68, -92, 48, -128, 35, 37, 118, 124, -94, 85, 24, -29, 78, 69, 64, 33, 78, 77, 18, -11, 74, -35, -73, 10, 42, -13, -35, -6, 27, -30, 116, -45, 12, -8, -117, 19, 125, 32, 111, -35, -35, -111, 17, 13, -103, -93, 52, 38, 28, 105, 99, -68, -13, -115, -94, 76, -76, 2, -64, 81, 80, 86, 48, -6, -78, 13, -79, 44, -31, 59, 85, 21, 54, 117, 58, 31, -119, -43, -76, 72, -121, -55, -90, -18, -112, 37, -29, 75, 43, 55, -128, -74, 54, 116, 121, 98, 25, 49, 5, 42, -47, -1, 32, 14, -75, 17, 72, -19, -111, -79, 44, 110, -4, 85, 99, 41, 85, -112, -40, 73, -106, -123, -44, -64, -54, -22, -83, -27, 98, -33, -127, -118, 34, 31, -104, 7, -78, -50, 107, 9, -64, 23, 126, 83, 72, -77, 67, -52, 46, 68, 64, -60, -32, -14, -83, -29, -43, -71, 97, 122, -96, 86, 88, -20, 90, 33, -47, -23, 95, -123, -1, -42, 84, -64, 126, 108, 37, 72, -32, 9, 29, -82, 124, 124, -80, -73, -35, 34, 28, -36, -70, -45, -99, 69, 110, -33, -101, -105, -109, 34, 100, 114, 72, 1, 21, -52, 51, 17, 38, 24, 55, -76, -51, 39, -104, 88, 107, 10, 22, 72, 60, 42, -88, 48, -120, -2, -92, 2, -98, 58, 116, 29, -14, -88, 55, 49, 79, -9, -70, 120, 123, 1, 19, -94, -125, -117, -6, -113, 57, -109, -18, -62, 123, -108, -118, -12, -21, -26, 63, 84, -15, -7, -83, -18, -37, -127, -29, -58, 29, -25, -20, 38, 83, -83, 99, 17, 4, 115, 19, -47, 93, -36, -76, -61, 98, 51, -22, 50, 41, 37, 83, -126, -59, 90, 54, -25, 91, 106, 107, -74, -72, -123, -18, 88, -47, -99, -121, 26, -86, -106, -110, -14, -117, -66, 102, 82, 36, -12, -14, 51, -80, 41, 89, -83, 8, 52, -55, 100, -116, -6, 70, -92, -44, -39, -62, 122, -112, 91, 100, -20, 124, -84, -22, 59, 125, -58, 108, -32, -9, -68, -81, 102, -109, -63, 84, 47, 99, -78, -14, 84, 1, 36, -114, -29, 13, -2, -4, 4, -128, 72, 2, 119, 81, 120, 1, -90, 46, 53, 115, -38, -54, 69, -111, -47, 112, -111, 104, 26, 47, 62, 92, -8, 92, -47, 9, 2, -2, -13, -32, 76, 88, 15, 74, -51, -106, 12, -64, -33, 52, 35, -66, 120, -63, 79, 56, -105, 100, 27, -118, -42, -66, 23, -46, -100, 100, 14, -19, 121, 53, -83, 31, 6, -119, -84, -43, -128, 55, 55, 93, -56, -31, 59, 71, 37, -39, 117, 13, 78, 76, -113, -101, 19, 105, -35, 79, -85, 63, 127, 127, -121, 93, -122, -66, -49, -27, -4, 85, -26, 1, -14, 1, 73, -63, 55, -82, -87, 94, -96, -37, 47, -58, 33, -17, 10, 19, -76, 106, 111, 36, 103, 2, -65, -97, -70, -29, -60, -22, -115, 71, 78, 114, 124, -14, -54, -74, 39, 22, -110, 22, -48, 65, -78, -88, 120, 67, 72, -42, 9, -83, 13, 44, -81, 110, 98, 81, 28, -74, -41, 101, -17, 36, -93, 40, -94, 74, 98, -73, -103, -32, -123, -39, -49, 71, 26, 40, 54, -7, 104, 100, -117, 43, 15, -100, -41, -95, 15, 52, 44, -72, 46, -125, 56, 106, -82, -34, 37, 79, -117, 1, -93, -76, 75, -56, -119, -19, -99, -126, 70, -72, -43, -85, -17, -37, 14, -119, 110, 43, -14, -59, 90, 68, 111, -40, 45, 80, 99, 93, 75, 70, -74, 8, 12, -101, -65, 36, 74, -103, -41, -3, -74, 32, 62, -10, 81, 86, -54, -8, -106, -92, 109, -108, -31, -116, -17, -85, 74, 10, -9, -103, -86, -5, 110, 68, -63, -29, -85, 0, 106, 119, -107, -14, 20, 80, 109, 69, 106, 127, 52, -55, -12, 31, -106, -70, 0, -79, -10, -38, -105, -63, -94, -127, 82, -35, -11, 71, -86, -78, 81, -79, 68, 32, 61, 1, -107, -93, 26, -38, 127, 87, -82, -119, 94, 27, -86, 38, 49, -8, 62, -78, 76, 38, 71, -15, 55, 71, 18, -69, 14, -15, 127, 81, -117, 68, 73, 38, -18, 29, -40, -17, -68, 73, 12, -42, 27, -44, 4, -126, -14, -92, -60, 19, 2, -33, 22, 2, -81, 72, 17, -45, 78, -113, 60, 56, 87, -119, -64, 60, 80, 95, -89, -42, 99, -32, -29, 0, -7, 40, 48, -66, -78, -118, -112, -95, -62, 78, 96, -65, 61, -48, -91, -108, 18, -79, -65, 41, -26, 93, 112, 121, -20, 5, -21, -71, -125, -25, 19, 115, 9, 112, -125, -54, 62, -117, 38, -113, -25, 89, -50, -97, 70, 100, 109, -118, -57, 59, 21, 59, -125, -115, -7, 54, -100, 98, 82, -90, 94, 47, 2, 125, 24, 55, 34, -102, -51, 75, -94, -46, -27, -44, -43, -41, -121, -17, -32, -10, 68, 75, -8, -53, -36, -107, -13, -78, -36, -56, 1, 53, -100, -89, 39, 89, -1, -60, 115, -127, -75, -124, 65, 94, 47, -28, -121, -21, 92, 109, -64, 91, 99, -22, -22, 122, -91, -34, 114, 100, -113, 6, 120, 79, -10, -84, 102, 1, 52, 69, 114, 17, -28, -107, 126, 114, -77, 99, -82, 41, -22, 124, 7, 51, 14, -45, -85, -103, 95, -27, -77, 55, 17, 103, -114, -103, 115, 52, 67, -10, -83, -114, 11, 9, -17, 96, 50, 105, 5, -38, 100, -37, 85, 71, -79, 54, 92, -103, -102, -18, 3, 16, -105, -95, 115, -119, -99, -20, -85, 67, -58, 74, 46, -112, 74, 115, 1, -32, -70, -120, 85, -68, 20, -71, -42, -30, 114, -88, -117, -40, 103, -10, 72, -7, -3, 13, 97, 3, -50, -66, 57, -64, 40, 14, -62, -95, 108, -5, -106, -73, -48, -34, 65, -38, -45, 100, -42, -26, 44, 120, -89, 78, -101, 75, -46, -108, -81, -39, -31, 62, -15, 68, -94, -126, 84, 16, 28, 82, 81, 61, 37, 39, -80, -49, -104, -70, 75, -48, -104, 68, -47, 125, -17, 83, 23, 73, 59, 106, 52, -111, 124, -91, 75, -41, -67, -120, 116, 107, -1, -55, 45, -16, -102, 2, 42, 114, 13, 60, -2, -56, -65, 40, -29, 29, -70, 7, 104, -112, -47, 41, -22, -4, -79, -4, -49, 81, -7, 122, 44, 20, -98, 53, 104, 14, -14, 73, -128, -96, 98, -117, -125, -118, -24, -88, 19, 106, 77, 32, -116, 66, -86, 35, 125, 39, 35, 85, -1, -84, -87, 101, -84, 70, -27, 49, -30, -21, -74, 2, 93, 8, -116, 38, -86, 62, 60, 48, 93, -117, -123, 65, 8, -17, 43, 93, 62, -84, -7, 54, 106, -121, 84, -24, -101, -86, -74, 121, -17, -6, -75, 63, -8, 97, 101, -19, -5, 8, 90, -2, -4, -124, 58, 2, -48, 66, 4, -100, -13, 81, 43, -101, -50, 23, 64, -75, -85, 6, 11, 9, 117, -44, -74, -62, 47, -89, -117, 45, 84, -66, 16, 11, 31, 49, 40, -65, -55, 38, -45, -110, 3, -44, -93, 71, 5, -126, 62, 108, 6, -61, -50, 42, 122, 26, -4, -18, 88, -104, -38, -48, -19, 3, 90, 32, 119, 58, 33, 31, -76, 1, 15, 121, 27, -91, -28, -57, 76, 14, 30, 92, 112, 46, -113, -121, 116, -79, -26, -55, 58, 126, -113, 94, 68, -98, 83, 2, 37, 72, -73, -87, -22, 50, 89, -25, 61, 24, 95, 73, -14, 49, 124, -23, -17, 85, -55, -88, 58, -70, -88, 86, 70, 113, -93, -27, -75, 98, -69, 38, 16, 106, 22, -84, 47, -21, -101, 47, -125, -13, 82, 45, -11, 9, -116, -55, -96, 29, 24, -17, 88, 117, -74, 45, 15, 61, -73, 123, -88, 119, -43, 16, -87, 9, -22, 10, 102, -105, -106, 46, -37, -20, -30, 87, 109, -112, 51, -38, -117, -37, 92, -34, -75, -104, -20, 42, 70, -120, -95, -45, -69, 87, 5, -3, -95, -86, 84, -5, -14, 75, -74, 58, -10, -92, 57, 21, -30, -7, 87, -76, 12, -90, -90, -6, -25, -3, -113, 100, 24, -23, 92, -109, -100, 125, 31, -52, -50, -41, 57, -91, 119, -105, -10, -99, -84, 3, -97, 41, -36, 100, 21, 2, 24, 88, 99, -8, 123, -62, 63, -115, 95, 122, 10, -13, 0, -22, -4, -106, -109, -75, -28, -92, 95, 116, 10, -118, -20, -37, -80, 106, 116, -37, -43, 57, -81, -72, 8, -94, -47, 95, -1, 70, -119, -50, -90, 44, 44, 21, 127, -65, -66, 59, 1, 111, -127, -89, 96, -99, -92, 14, -99, 17, 31, -113, 109, -101, 111, -38, 55, -72, 50, 18, -82, -25, -6, -110, 26, -124, 34, 63, -98, 27, 14, 17, 30, 120, -64, 114, -66, 126, 38, 4, 50, 39, -109, 77, 88, -111, 86, -125, 62, -54, 107, -115, -112, -65, -103, -20, 82, -45, -3, 123, 4, -36, 24, 88, -33, -83, -34, -81, 88, 121, 110, -125, 38, 125, -58, 77, -40, -4, -21, -67, 78, -114, 66, -77, -70, 1, -57, 117, 126, -83, 103, -75, -84, 77, -80, 34, -36, -43, -58, 64, -86, 80, -30, -105, 69, -11, -80, -25, 5, -70, 48, -38, -41, -59, 77, -118, -88, 9, 111, -76, -49, 42, 36, -84, -128, 5, -37, 37, 118, -100, -79, -77, -5, -44, -10, -69, 106, -71, 126, -79, -74, -48, -23, -76, 37, -23, 61, 74, 31, 64, -21, 15, -86, 30, -24, 62, 36, -99, 40, -119, -128, 62, 1, 51, -23, -43, 25, 108, -23, 126, -32, 90, 59, 49, 118, 96, -93, 86, -114, -5, -26, 71, 7, 36, 5, -35, -14, -78, -20, -124, 84, 41, -125, -126, -63, 127, 106, -45, 74, 24, -49, -77, 57, -79, 126, 57, 92, -110, 123, -84, 41, -38, 42, -117, 67, 115, 23, -61, -23, -121, 103, 29, -48, 34, 36, 94, -70, -10, 52, -48, -53, 70, 11, 6, -99, 65, 123, -35, 41, -109, -95, 17, -40, -117, 119, 113, 95, 5, 45, -32, 83, 79, 116, 41, -26, -102, -127, 122, -9, -16, -119, 21, -56, 72, 19, -34, -93, -58, -88, -106, 41, -34, -1, -77, -101, 24, 17, 40, -48, -62, -46, 14, -56, -92, 80, 26, -85, -86, 78, -56, -38, -86, 50, 11, -59, 53, 42, -73, 122, 7, 86, -27, -61, -71, -110, 92, 55, 79, 8, 101, -8, -26, 40, -32, 50, -49, 23, 106, -49, -26, 11, -45, 126, 35, -93, 59, -115, 53, -123, -8, 37, -26, -21, -12, -122, 90, 104, -24, -75, 17, -93, -119, -10, 106, 66, -41, 51, 19, -11, 95, -35, -27, -40, 82, -48, -26, 36, -80, -80, -53, -27, -59, 15, 85, -48, 10, 0, 2, 111, -107, 127, 11, 40, -32, -120, -115, 28, 92, 21, -53, -11, 14, 49, 39, 114, -50, -43, 122, -68, 27, 23, 19, -53, 34, 87, 13, -83, -50, -42, -63, 35, -79, 91, -122, -82, 4, 16, 94, 92, -8, -105, 28, 32, 112, -121, -75, -73, -16, -127, 19, -85, -31, -3, -32, 123, 39, -125, 101, 61, 25, -124, -83, 94, -36, -107, 106, -119, -5, 1, 118, -53, 84, -29, 113, 39, 40, 5, -121, -121, 57, 119, -55, -125, 46, 2, 124, -60, 92, -71, -82, 34, -109, -93, -68, 90, -53, -72, 76, 104, -109, 9, 108, -18, 59, 20, -127, 90, -17, 90, -127, -31, -107, 61, -32, 47, 42, -38, 23, 88, -12, 124, -66, -12, 123, -14, 26, -37, 84, 45, -64, 118, -81, 90, 62, 91, -39, -8, 12, -109, 24, -39, -24, 83, -59, -45, 94, 15, -117, -45, -125, -121, 57, 87, 87, 125, -43, -52, -18, -49, -97, 119, -36, -120, -102, 93, 95, -100, 70, -7, 102, 102, 57, 75, 28, 35, -127, 36, 12, -37, 43, 20, -122, -9, 90, -61, -125, -7, -42, -36, 53, 21, 85, 78, -111, 45, -125, 2, 63, -16, 111, -68, 26, -9, -4, -45, -96, 5, -119, 109, 12, 34, -15, 115, 19, 25, 125, -56, 17, -62, -94, 52, -126, 2, -47, 14, -58, -91, 126, 27, -44, 26, -80, -91, 26, 36, -70, 33, -44, 89, -60, -90, -106, -11, -63, -117, 68, -14, 98, 34, 5, -125, -19, -123, 50, -99, 92, 48, -115, -73, 99, -5, -6, -82, 60, -99, 93, -45, -1, 47, -66, 109, -101, 89, 63, -97, -56, 49, -119, 108, 95, 119, 3, -81, 74, -61, 98, 43, -115, 67, 111, 44, -105, -58, 74, -47, 120, -34, 48, -79, 17, 68, -4, -93, -13, -17, 10, -120, -121, 21, 46, 66, -97, 44, 35, -106, 105, 33, -73, 75, 120, 74, -50, -56, -43, -84, -82, 122, -48, 44, 101, -97, 81, 72, -46, -95, 15, 66, -80, 83, 123, 11, 120, 14, -4, -26, -37, -56, -53, 30, 63, -7, -81, 103, -58, -74, 77, -87, 96, 18, -119, -60, 12, 4, -32, 34, 4, -57, -17, 109, -15, -127, -112, 6, -54, 70, 15, 67, -103, 101, -80, 41, -86, -91, 67, 3, -6, 61, -116, -44, 88, 99, -91, -68, 90, 87, -16, -58, -47, -125, 15, -60, 26, -94, 111, 73, -31, -77, -77, -89, 11, 55, 16, 100, -25, -94, -22, -17, -61, 50, -56, 78, -18, 19, 61, -56, 1, -44, -17, -75, 125, -73, 87, -87, -102, -27, -7, -107, 40, 113, -57, -102, -31, 127, 30, -22, -102, -12, 30, 107, 24, -21, 61, 86, 94, -84, 103, 90, 39, 109, 14, 65, 90, 79, 97, -109, 39, 56, -1, 17, 96, 51, -44, -21, -90, -6, 79, -43, -64, -2, -11, -8, 58, -22, 111, -66, -128, -66, -40, 28, -42, -12, -39, 58, 119, 114, 111, -114, 16, -46, 86, -128, -87, 124, -4, 78, 46, -81, 75, -74, -78, 66, -8, -94, 66, 68, 81, 48, -106, 58, -58, -49, 92, 112, 24, -121, -55, 84, -10, -120, -116, 84, 59, -42, -85, -111, 60, 13, 50, -4, -115, 8, -108, 78, -32, 107, -79, 27, -77, 126, 33, -16, -61, -83, 60, -29, -53, -54, -20, -80, -83, 33, -70, -40, 9, -96, -30, -95, 115, 117, -36, 88, 63, -125, -50, -72, 46, 62, 69, 42, -15, -34, -77, 124, -84, 123, -91, 103, -67, 61, -117, 8, -128, 84, -114, 24, 126, -72, -9, 23, -84, 107, 47, 60, -32, -63, -19, 25, -94, -56, 80, 66, -91, 9, -57, 81, -110, -58, 4, -94, -105, 0, -74, -116, -102, 26, -116, -65, -80, -16, 8, 127, 86, -80, 60, -128, -110, -126, 15, -73, -67, 109, 8, -126, -103, 37, 95, -39, -85, -56, -73, 105, -24, 76, 91, -45, -38, -102, 61, -87, -36, 39, -10, -82, 96, -87, -109, -50, 108, -107, -94, 67, -126, 102, 114, 36, -26, -60, -87, 46, -52, -60, -79, -79, 81, -7, 70, 90, -109, -105, -6, 100, 49, -75, -22, -117, 75, 66, 49, -106, 30, -103, -52, 87, 7, -82, -101, 99, -122, 36, 36, 70, 40, -93, -56, 6, 35, -4, -27, -120, -118, -44, 82, 95, -107, -112, -109, -114, 99, 94, -95, -30, -55, -17, -37, -97, -97, 101, 3, -31, 6, 45, -33, -94, -90, 110, 102, -84, 116, -113, 88, 19, -110, 125, -68, 58, -53, 118, 68, -58, -13, -123, 9, -82, -90, -117, 101, -73, -36, 34, -128, 104, -4, 108, -82, 110, -43, -114, -94, -93, -109, -29, -104, 50, 125, -128, -15, 19, 39, -123, -69, 94, -98, 90, 84, 11, 37, 74, 108, 113, -55, 51, 42, -117, -3, -6, -126, 51, 47, -31, 120, 11, 53, -28, -106, -108, -9, -107, 34, 114, -51, 124, -11, -16, -14, -42, 123, 42, 84, 41, -4, -85, -50, 33, 47, 2, 31, -13, -27, -92, -118, 96, 73, -120, 99, -31, 37, 109, -41, 30, -99, -126, 0, 68, 102, -95, 52, -9, -127, 98, -6, -15, 74, -26, -11, 31, 70, -81, 60, -20, 8, -27, 121, -112, -71, 114, 68, -117, 69, 108, 69, 7, -108, -45, -73, 116, 18, -30, 69, -98, -117, -57, -119, -33, 82, -20, 35, 37, 81, -99, -111, 97, 22, 45, -24, -55, 121, -32, -100, -79, -54, -126, -47, 113, -6, 1, -102, 111, -82, -19, -127, 99, -61, -52, 28, -1, 35, 9, 11, 90, 86, -124, -12, -84, 109, 42, 52, 1, 13, 64, -116, -57, 102, -79, 66, 44, 62, 117, -45, -128, -98, 102, 57, -125, -59, -85, 105, -121, -91, 92, 1, 95, -74, -57, 121, 53, -78, -56, -104, 8, -121, 68, 68, -52, 96, 101, 36, -108, 52, -125, -82, 96, -32, -91, 14, -24, 76, 45, -13, 29, 110, -60, 91, 68, 72, 57, 18, -84, -66, -124, 40, -5, 89, 8, 15, -45, -68, -61, -23, -62, 38, 100, -81, -58, 51, 9, 83, -89, -70, -2, 16, 88, -33, -120, -89, 118, -102, -127, -121, 102, 43, -53, -27, -54, -84, -40, -10, 70, -39, 60, 34, 16, -113, 10, -76, -88, 47, 115, 46, -53, -41, -84, -32, -58, -32, 90, -112, -66, -112, 84, 54, -124, -58, 82, -73, 38, -25, 5, 42, 66, 126, -93, -115, 107, -25, -37, -10, 6, 111, 73, 88, -38, 121, 21, -110, -78, -76, 44, -62, -46, -64, 31, -58, 49, -53, 115, 75, -85, -14, -125, -73, 31, 84, 103, -106, 20, 24, 47, 39, 10, -52, -49, -63, -46, -31, 14, -35, -112, 70, 8, -60, 6, 127, 102, -5, -102, -68, 39, 114, -54, 104, 115, 40, -55, 38, -76, 13, 26, -82, -68, -43, -85, -72, -45, -28, -14, 49, 20, -90, 51, -78, -62, 127, 122, 55, 90, -70, 30, 95, 32, -85, 18, -128, -113, -81, -110, -86, -30, 125, -127, -33, -65, 121, 22, -64, -82, -10, -66, -18, 80, 1, 107, 26, 57, -59, -112, -112, -15, 107, -109, -88, 73, 111, 126, 68, 44, 26, 123, -39, -113, -42, 1, 29, 43, 123, -79, -118, -93, -116, 77, 20, 35, 97, 63, -108, 79, -116, -57, -49, 49, -8, -55, -74, 70, 96, -85, 4, -112, 35, -79, 68, 95, -60, -102, -3, 69, 13, -62, -38, -13, 106, 2, 78, -119, -74, 6, 39, -54, -127, -10, -118, 4, -103, 22, 87, 68, -87, 45, 88, 110, -62, 111, -57, -48, -63, -27, -117, -4, -49, 20, 11, -126, -88, 68, -121, 82, 109, 3, -103, 36, 48, -44, 18, -15, 77, 31, 104, 57, -28, -83, 27, 11, -117, 98, -103, 30, -34, -56, -60, -113, 4, -97, -14, 109, 125, -121, 110, 21, 102, 118, 43, 22, 72, -64, -87, 33, 106, -11, -33, 32, -99, -88, -15, -95, -111, 34, -55, -89, -4, -76, 18, -77, -60, -25, 110, -70, 9, -81, 5, -35, 8, 2, 73, 75, -6, -67, 43, -109, 56, 45, 45, 62, -83, 125, 87, -111, 70, -115, -75, 107, 28, -112, 32, 95, 124, 35, 10, 107, -43, 97, -58, -45, -51, -23, -101, -35, -120, -26, 114, -35, 44, -23, -44, -83, 12, 107, 26, -28, 49, -90, 34, 7, -17, 117, -102, -90, 32, -31, 18, -100, -113, -88, -60, 58, 64, 38, 12, 119, 41, -56, 79, 21, 41, -72, -2, -119, 27, -10, 21, -11, 75, 105, 12, -68, -33, 46, -31, -49, 118, 47, -69, 5, -116, -116, -25, 68, 99, 82, 95, 95, 57, -125, -35, 93, 37, 104, -62, -59, -46, -105, 54, -120, -40, 124, -92, 126, -110, 2, -2, -90, 0, 124, 33, 33, 22, 66, -60, 44, -36, -7, 90, 125, -92, -71, 91, -20, 93, 34, -36, 41, -120, 19, 20, -112, 88, 100, -125, 122, -58, 4, 19, 52, 45, 89, -110, -118, 114, 55, -118, -36, 76, -85, -69, -73, 76, -19, -91, -36, 29, 0, -109, 82, 100, -37, 89, 82, 14, -115, 59, -52, -15, 64, -123, -33, 126, 102, 58, 12, -24, -17, 38, 99, -126, 68, 56, 95, -66, -61, -102, 107, 70, -108, 126, -75, -11, 94, 78, 3, -67, 81, 44, 109, 122, 35, 19, -91, 14, 63, 19, -115, 94, -91, 72, 53, 120, -2, -34, 1, 54, 119, -87, 116, 77, 93, -21, -24, -108, 99, -33, 85, -74, -121, 79, 75, -98, -23, 78, 101, 108, 41, -42, -46, 70, -59, -108, 16, 122, 80, -1, -104, -88, -5, -6, -17, 124, -126, -2, 95, 6, 68, 103, -57, -90, -41, -81, -51, -9, 39, -52, 19, 73, -97, 126, 9, -71, -25, 32, 34, -76, 72, 7, -89, -18, 61, -109, 63, -32, 92, 48, -122, 79, -54, 18, -38, 48, -3, 120, 40, -118, 44, 99, 67, 0, 30, -4, 126, 94, 82, 32, 38, 22, -115, 75, 83, 116, -111, 61, 54, 90, 78, 54, 29, 98, 25, 96, -124, 120, -36, -4, -96, -64, 88, -2, 40, 19, 115, -125, -21, 64, -125, 74, -91, 64, -107, 52, -30, 42, -123, -101, -4, -69, 32, -95, 108, 45, -97, -4, -115, -62, 56, -11, 4, -63, 60, 63, -123, 121, 115, 89, -30, 126, -99, -93, -45, -38, -98, -118, -35, 0, 66, 32, 60, -99, -2, 94, -127, -21, 91, -114, -15, -10, 13, -2, 22, -102, 113, 73, 127, 123, -54, -102, 81, -102, -88, 43, -78, -9, 38, 50, 86, 17, 56, -92, 33, -75, 127, -87, 48, 91, 108, -53, 114, 126, 65, -120, -41, -52, -85, 97, 85, -65, -43, -18, 12, 42, 113, 92, -58, -126, 30, 80, 58, -38, 76, 38, 42, 90, -45, -71, 35, 70, -83, -85, 42, 101, -12, -77, -107, 0, -93, -105, -120, 98, 1, -49, -127, -110, -85, 58, -3, -115, 44, -76, 52, 39, 78, -9, 101, 5, -92, -60, -30, -75, 9, -6, 28, -106, -14, -106, 59, 52, -27, 2, 68, -25, -100, 17, -50, -40, 112, -29, -88, -125, 102, -119, -4, 30, 116, -58, 110, 84, -85, 90, -102, 86, -21, 124, 38, -13, -103, 119, -60, 14, 27, 53, -43, -86, 80, 56, -128, 78, -100, 39, 77, 39, 127, -116, 81, -7, 50, 8, -52, 30, 126, 92, 72, -87, -95, 126, 122, 18, 119, -127, -45, -37, -2, 38, -35, -122, 25, 76, -25, 70, -115, -30, -8, 58, 66, -70, -26, 86, -75, -10, -40, -106, -82, -24, -126, -66, 42, 66, -14, -17, 47, 42, -117, 114, 97, -83, -35, -84, -57, -19, -116, 7, 101, 118, 125, -53, 108, -102, 81, 83, -58, -71, 68, 59, -58, -58, -120, 119, -107, -111, -11, 79, 76, 57, -36, 7, -118, -19, 28, -65, -15, 81, -68, -48, 66, -15, 87, -102, 85, -30, -126, 86, 125, 20, 4, -41, 14, 58, 10, -5, -103, 100, 54, -13, -53, -95, 18, 124, 12, -47, 47, 22, -67, -74, -112, 77, -99, 98, -108, -123, -30, 110, -97, 40, 84, 113, 34, -59, 48, -99, -87, 88, -110, 57, -10, -43, -122, 4, 123, -2, 87, 67, -115, -52, 51, -77, -113, -24, -114, -53, 111, 29, -107, 87, -57, 90, -112, -94, 76, 77, 69, 94, 82, -60, 87, -37, 84, 59, -24, 8, -84, -106, 43, 118, -61, -32, 7, -114, -127, 118, 117, -53, 12, -62, -48, 6, -6, 58, -81, -17, -16, 78, -59, 97, 29, -73, -124, -96, -116, -52, 121, 80, 74, -116, -15, 30, -27, -101, -7, -59, -25, -62, 90, -21, 67, 37, -85, 116, 32, 10, -125, -74, 10, -75, -18, -34, 74, -112, -15, 4, -121, 124, 111, 105, 111, -75, 72, -56, 59, -64, -24, -34, 68, 50, -58, 51, 28, 54, -122, -10, 33, -62, 2, 114, -54, -101, 68, 0, 44, 29, 21, 70, 58, 111, -91, 21, -107, 52, -108, -110, 37, 62, -70, -78, 126, 26, -120, -24, -67, 85, 38, -28, 78, -24, 13, 38, 40, 71, 49, -28, 14, -47, 111, 66, 70, -84, 39, 94, -108, 52, 24, 44, -7, 71, -55, 5, 121, 127, -13, 26, 10, -120, -85, 71, -13, -11, 119, -79, 52, 120, -9, 30, -94, -29, -8, 115, -128, 85, -9, -93, 9, 2, -12, 68, -58, 25, -66, 40, 58, 51, 39, 94, -43, -125, 116, -57, -128, -22, -3, -31, 21, 119, -97, -112, 85, -85, -30, -91, 60, 76, 24, -65, 118, 77, -84, -75, 58, -52, 10, -91, -122, 74, -106, -41, 119, 73, 114, 51, -42, 87, 85, -97, 24, 111, 47, 101, 102, -112, 54, -117, 4, 30, -63, 77, 21, 17, 27, -24, -127, -113, 56, -47, -128, -31, 23, -87, 50, -11, 112, -89, -5, 80, -104, -54, 17, 36, 43, -94, 110, -10, -36, -70, 120, 107, -4, -36, -6, 43, -29, -95, 113, 84, -30, -86, 118, 46, 20, -57, -48, 41, -15, 13, -62, 81, -105, 63, -12, -47, 70, -57, 30, 65, -128, 113, 34, 66, -127, 91, 124, -71, -111, -100, 90, 1, 44, -34, 38, -98, 110, -3, -122, -115, 98, -14, -61, 1, 113, 11, 11, 1, -10, -126, -95, -61, 39, -19, -42, -20, 33, 61, 127, -80, -24, -83, 56, 1, -58, 93, 88, -118, 33, 122, -58, -10, -94, -28, -4, -114, 68, 0, 51, -45, -52, -27, -117, 38, -47, -116, 37, 67, -79, 51, -59, 21, 41, -10, 126, -108, 122, 16, -107, 5, -119, 92, -19, 70, -107, -14, -55, -106, 45, -9, 35, -11, 108, 99, -91, -2, -72, 122, 5, -55, 98, -110, -32, 13, -83, 37, 113, 100, 54, 48, -123, 4, -124, 96, 41, 3, 121, -63, 86, 102, -100, -5, 65, 42, 104, 72, 58, -42, -126, 95, 41, -93, -55, 93, -66, 4, -49, 79, 117, 60, -110, 66, -66, 93, -30, 10, -23, -94, -69, -114, -62, 89, -77, 126, 110, 82, 12, 72, 84, 42, 59, 75, 58, -100, -123, -46, -70, 33, -2, 10, -16, 31, 12, 102, 43, -100, 114, 99, -74, -42, 68, 105, -68, 106, -104, -118, 25, 126, 11, -63, -30, 85, 64, -111, 45, -32, -85, 81, 8, -124, 38, 43, 98, -52, -37, -60, 122, 105, -110, 35, -127, 116, 55, 11, 7, -61, -100, -34, -11, 78, -111, 61, 123, 25, 84, 13, 109, -37, -111, 120, 57, -31, 77, -58, -58, 23, -46, -128, -18, 13, 63, 39, -83, -22, -61, -22, -124, -39, 107, -64, 126, 50, -28, -23, 22, -13, 109, 30, -8, -6, -14, -17, 1, 52, -122, -68, -126, -28, -24, 11, 12, 85, -105, -123, -44, 122, -31, -50, 85, 45, 93, -35, -114, 41, -49, 116, 118, 80, 49, -55, -44, 25, 27, 42, 6, -26, 75, -45, -96, -52, 110, -58, -37, -108, 8, -66, 122, -53, 82, -100, 69, 64, -35, 80, -53, 35, 54, -64, -96, 49, -56, 47, 8, -122, -42, 40, -95, 89, -126, 78, 116, -3, 11, -75, -37, 28, 117, -91, 54, 50, 36, -84, -3, -87, 119, -45, 116, 8, 6, -103, 8, 96, 101, 61, 56, 115, -114, -97, -69, -124, 23, -55, -25, 104, 102, -1, 37, -126, 74, 39, -8, 107, -74, -64, 75, 68, -83, -77, 63, -24, -40, 32, -86, 114, 82, 75, -114, -90, -112, -74, -112, 43, -75, -59, -31, 77, 10, 48, 31, -108, 71, 99, -125, -123, -12, 13, 5, -65, -42, -11, -29, -39, 127, -77, -27, -111, 3, -114, -51, 119, 72, 78, -102, -41, -26, -38, 91, 1, 5, 55, 108, 62, 87, -112, 76, -21, 115, -12, -62, 114, -36, -58, -26, -15, 56, 53, 119, -32, 108, 67, 42, -24, 126, 34, -35, -26, -104, 52, -102, 1, 1, 79, 26, -128, -81, -128, 57, 57, -31, -34, 120, 84, 50, 48, 55, -14, 88, 80, -82, -108, 121, -10, 108, -44, -12, -89, -7, 5, -23, -50, 68, 22, 80, -56, -114, 2, 12, -47, 13, -95, 38, -63, 90, -126, -1, -61, -62, -50, -38, -50, 104, -92, -46, -17, 127, -128, -51, 89, -51, 107, -68, 3, -50, 49, -91, -127, 37, -45, -29, 77, 19, 78, -73, 22, -118, 7, -3, -100, -106, -104, -53, 117, -122, -56, -117, 63, -77, -41, -63, -55, 58, -109, -29, 39, -73, -45, -92, 41, 10, -22, -122, 0, 22, 28, 36, -79, -40, 114, 37, 72, 67, -85, 34, 79, 47, 113, 19, 102, -127, -37, -55, -31, 14, -3, -76, 101, -57, 31, -8, 81, 60, -70, -113, 27, 16, -6, 108, -2, 113, -89, 125, 85, -89, -76, -76, -26, 72, -109, 79, -21, 46, -52, -121, 68, -67, -70, -94, 77, 118, 40, 117, -88, -77, 96, 88, 55, -112, 37, -1, -34, -106, 44, -100, -29, -114, -33, 113, -98, -115, -33, -57, 122, 9, 28, 55, 120, 89, 74, -22, -37, -88, 43, -69, -102, 35, 101, 7, -84, -71, -24, 35, -116, -69, -35, -44, 85, -110, -101, -70, 85, 10, 115, -86, -87, 2, 109, 36, -29, 37, 120, -98, -19, -87, 42, 64, -12, -79, -82, -89, -95, -72, 40, -106, -48, 60, 61, 90, 120, 65, -112, -92, -84, -16, -121, 48, -4, -5, -52, 106, -32, -76, 61, -41, 66, 99, -38, -108, 58, 79, 80, -45, 99, 35, -84, 89, 9, -119, -93, -43, -58, -3, -48, -23, -47, 69, -53, -101, -15, 80, -12, 125, 93, -113, -96, 110, 87, -86, 117, 92, 44, -45, 29, 115, 14, -64, 105, -94, -79, -51, 25, 68, 10, -128, 48, -7, -56, 93, 100, -38, -85, -53, 110, -8, -52, 117, 76, 89, -39, -78, 46, 86, 102, -34, 43, 51, 18, -126, 75, 2, 36, -27, -44, -67, -32, 96, -105, 111, -15, -112, -96, -102, 9, -6, -26, -43, -80, 103, -121, -113, 127, -118, -26, -53, 43, -27, 90, 24, 89, 90, 7, -128, 121, 29, -4, 118, -76, -21, 68, 122, -76, -64, -26, -78, -21, -118, 3, 46, 104, -104, -105, -77, -124, 100, 75, 83, -61, -125, 70, -33, 109, 64, 43, 22, 27, -124, 1, -90, -109, 19, -72, 48, -125, -126, 57, -63, 97, -28, 100, -92, -17, 79, -54, 92, 64, -16, 32, -72, 104, 36, -22, -67, 83, -58, -98, -112, 46, 69, 105, -101, 118, 10, -59, 77, 73, 26, 122, -81, -62, -40, -86, 103, 68, 25, -64, -24, 9, -3, 80, 44, -102, 67, 118, -25, 53, -96, 51, -71, 124, 32, 75, -91, -72, 84, 73, -96, -23, -125, 116, 69, 59, 107, 15, -64, -108, 85, -103, 6, -122, 53, -110, -24, -39, -104, -9, -56, 84, -127, -77, -17, 19, 27, -7, 103, -44, -37, 3, -72, -3, -80, 21, -111, 103, 112, -85, -125, -33, 106, 68, -28, -30, -29, -31, -3, 17, -11, 101, -85, 90, -104, 59, -111, 21, 97, -93, 105, 62, -90, -72, -108, 43, 123, -3, 12, -2, -107, -36, 126, -77, 67, -36, 16, -68, -41, 124, -67, 74, -46, -49, -117, -125, 65, -40, -22, 104, -99, -18, 57, -10, -17, 25, 65, -10, -14, 28, 23, -109, 117, 44, 104, 54, 116, 125, -13, -54, -121, 96, 99, -28, -102, 27, -126, 38, -44, 35, 54, -26, -115, 3, -81, -52, 112, -43, -39, 72, -84, 3, 20, 37, 92, -78, 7, 73, -93, -74, -9, 111, -65, 68, 4, 78, 67, -58, -104, -114, 15, -58, -94, -84, -74, 75, 45, 116, -103, 115, 85, 60, -102, -72, 78, 96, 55, -12, -10, -103, 72, -97, 101, -60, 111, 44, 14, -24, 104, -43, 61, -96, -55, 11, 85, -72, -82, 127, -81, 60, -30, -55, 52, -55, 36, -40, 0, 103, -92, 25, 89, -125, 23, -127, 45, 31, 73, -85, -125, -99, 83, -1, -64, -49, 24, -94, -52, -79, 102, 66, -126, -6, 94, -20, -48, -70, -95, -32, 28, -120, -18, -7, -91, -95, 71, -88, 119, -28, 60, 4, 18, -49, -105, -104, -94, 33, 56, 87, 30, 27, 72, -2, 84, -102, 58, 96, 34, -6, -21, 103, 81, -95, -123, 76, 90, 59, -106, 122, -116, -102, -44, -5, -79, 52, -107, 113, 114, 43, 71, 56, -128, 82, 127, -41, -92, 79, 77, -34, 124, 16, -99, -47, 80, 26, 97, 83, -87, 107, 39, 85, -120, -42, 103, -108, 4, 122, -102, -63, 85, -68, 46, 123, 27, 79, -17, 34, -122, -68, -2, -62, -115, 96, 99, -56, 83, 93, -119, -64, 30, -92, -53, 34, -41, 87, 45, -49, -26, -121, 121, 79, -14, -43, 71, 61, 56, -11, -93, 43, 121, 6, -72, -107, 114, -48, -33, -81, -8, -81, 8, -72, 18, 69, 14, 34, 8, -78, -101, 53, 77, -100, 113, -21, -68, -54, -14, 102, -65, 46, -92, -44, 61, -110, -123, 103, 38, -98, 107, 11, 65, 0, 10, -97, -125, -71, -110, -90, -14, -1, 6, 88, -17, -57, 40, 26, -26, -2, 34, 108, 6, -113, 44, -49, 54, 18, 61, -92, 125, -125, 117, -73, 61, 69, -21, 66, -41, 22, -87, -128, -104, 39, 72, -114, -42, 95, -93, 107, -100, 0, 77, 62, -102, -13, -67, 94, -19, -12, -123, -44, 24, 69, 37, 97, 72, 0, -95, 58, 116, 53, 66, -75, 55, -100, -7, 20, 123, -9, 113, -32, -13, 75, -63, 48, 55, 30, 39, 14, 17, -113, -57, -15, -10, 46, 123, -50, 71, -39, -84, -79, 74, -72, 52, 5, 75, -86, 96, -55, -49, 3, -3, 123, 28, -92, 84, -6, 3, -92, 13, 8, 120, 30, 94, 84, 123, -97, 13, -107, -5, -71, -57, 105, -125, 108, 98, 127, -79, 40, 111, -66, 22, -34, -89, -116, 15, -57, -26, 114, -80, -84, 99, -46, 101, 72, 53, 57, 96, -109, -64, 35, -30, -18, -86, 45, 126, -23, 115, -21, 14, -3, 71, 100, 80, 113, -9, 32, -53, 41, -123, 92, -113, 28, 116, 15, -94, 62, -113, -119, -93, 67, -50, 4, 59, -112, 41, 63, -116, 1, 63, 45, -41, -12, 18, 115, -72, 54, 33, -48, -74, 6, -74, -21, -97, 71, 103, -121, -67, -19, -15, 99, -91, 103, -74, 14, 110, -104, -58, 36, 10, -79, 37, -21, 5, 63, -3, 62, 6, -103, -14, 73, -128, 105, 17, 127, -45, 114, -36, -15, 102, -83, -94, 65, -97, 95, -55, -26, -68, 6, -34, -49, -126, -96, -40, 126, -107, 116, 76, 108, -111, 57, -115, -113, 70, 24, 124, 11, -71, -89, -3, -82, 56, -102, 122, -108, -75, -92, -58, 37, 31, 69, 101, 86, 71, 82, -38, 48, 71, -60, -72, 119, -18, -88, 106, -96, 89, -78, -90, -39, 14, 54, -94, 35, -128, -118, 15, 88, 19, 64, -64, -20, -61, 105, -65, -3, -96, 61, 87, -77, 22, 2, -96, -84, -52, -60, -33, 54, -98, 82, 18, -81, -54, 64, -114, -57, -42, 125, 79, 114, -92, -85, -28, -2, 5, -81, -126, -122, 5, -17, 83, 1, 43, -15, 64, 42, -99, 83, 37, -118, -41, -127, 85, -55, -43, 113, 6, 82, -29, 123, -18, -92, -119, -73, 121, 11, -111, -80, -72, -120, -28, -89, -94, 56, 1, 56, -101, 24, -107, 25, -128, -61, 18, -4, 55, 103, -43, -83, -105, 121, 76, 96, -5, -81, 46, -100, 67, 16, 59, -19, 60, -53, 112, -105, 110, 75, -119, 77, 36, -45, 64, -66, -100, -12, -73, -87, -121, 47, -92, 102, -16, -122, -21, 79, -43, 18, -18, -111, 106, -8, 34, 53, -112, -8, -85, -85, -5, -33, 83, 78, -56, 55, -8, -120, 60, -18, 91, 127, -126, 94, -90, -45, -17, -36, -68, -79, -77, -2, 5, 89, -55, -46, -61, -75, -20, 33, -23, -111, 2, 76, -125, 27, 44, -5, 3, 29, -86, 68, 1, 1, 38, -93, -125, -14, 47, 58, 24, 7, 121, -2, 115, -98, -17, -125, 107, 41, 31, -119, -74, -20, -65, 36, 73, 1, 93, -76, -76, 65, 7, 125, -65, 68, -7, -2, -62, 35, -48, 97, 15, 98, 109, -27, -127, 74, -37, -97, 22, 39, -108, -33, -124, 55, 64, 120, 89, 21, -95, -56, 33, -111, -9, -37, -92, -21, 90, 117, -124, 15, 110, 109, 24, 18, 115, -32, -127, 21, -87, -91, 100, 66, 105, -114, -63, 111, -20, -97, -99, 77, 80, -25, -46, 18, -119, -110, 59, -55, 55, -17, -104, 66, -84, 68, -68, 102, -82, -94, 32, 125, -37, 109, 77, 59, -128, -34, -45, 122, -38, -105, -101, -77, -2, -106, 17, -5, 19, -98, -40, -13, 18, 53, 105, -28, -31, -106, 50, 125, -67, -120, -111, 120, 81, 57, -85, 72, 53, 97, 65, 105, 85, -21, -42, 10, 61, -8, 46, -62, 78, 93, -125, -100, -41, 83, 2, 60, 6, 82, -75, 76, 51, -9, -95, -58, 8, 2, 52, -69, -59, -50, 67, 5, -25, 23, 23, 51, 70, -110, -47, 12, -83, 41, -3, 24, -78, 101, 13, 93, -89, -102, 36, -66, -2, 47, 7, -19, 78, 20, -47, -97, 72, 34, 102, 17, -78, 54, -80, 30, -120, 2, -5, 70, 44, 43, 0, 87, 13, -21, -11, 114, 127, -82, -121, -94, -106, -26, -110, 125, -123, -126, -67, 18, 53, 112, -63, -82, 106, 57, 57, -5, -75, 106, -40, 51, -9, -52, -15, 90, 30, -52, 55, 105, 114, -80, 119, 120, -78, -1, -74, 105, -81, 67, 101, 54, 106, -123, -77, 41, 18, 56, -81, 107, -121, -38, 61, -76, -48, 66, 110, 85, 72, 101, -71, -124, 110, 10, 84, 45, 122, 57, -9, 19, -32, 107, -61, 1, 95, 102, -95, 24, -115, -69, 53, 4, 80, 96, -31, -9, -69, 93, 42, -14, -125, -69, -95, 44, 40, -10, -25, -26, 86, 99, -86, 67, -114, -66, 23, 60, -58, -111, 112, 5, -54, 110, 87, 9, 20, 95, 23, -79, 47, 90, -88, -99, -84, -51, -7, -37, 8, -48, 99, 49, 57, 81, -7, -13, -45, -9, 74, -47, -83, -123, -23, -5, 108, 88, -49, 89, 109, 54, -119, -40, 38, -44, -82, -12, -50, 89, -39, -106, 102, -37, -6, 120, -88, -28, -30, -112, -115, 16, -96, 27, 39, -75, -128, 98, -77, -93, -41, 113, 38, -92, 79, -14, 95, 82, 25, 109, 72, -119, -125, -52, -21, -66, 59, -63, -95, -4, 87, 75, -20, 122, 105, 65, 116, 30, -30, 78, 94, 14, -25, -93, 113, -60, 17, -96, -104, 1, 92, 66, 27, 8, 113, 113, 17, -25, -95, 101, 99, -41, 38, 65, -15, 108, 54, -95, 114, 99, -16, 56, -113, 94, -108, 54, 28, 70, 92, 86, 82, -16, -92, -89, -1, 48, -47, 14, -49, 64, 80, 79, -11, 26, -95, -61, -31, 41, -99, -64, -99, -114, 78, 51, 9, -52, 42, 2, -54, 107, 32, -108, -48, -60, 35, 38, 6, -43, 75, -38, -54, 35, 12, -72, -6, 110, -83, 118, 45, -50, -2, 122, 127, 127, -53, 1, 121, -63, 123, -34, 21, -62, -11, -81, -96, -5, -70, 125, -50, -4, 114, 37, 126, -50, 95, -60, 75, -61, -10, 50, -123, -24, -100, 61, -20, 63, 68, 73, -71, -118, 30, -34, -38, -83, -48, -55, -125, -96, 86, -57, -44, -118, -115, -32, -95, -55, -82, -115, 4, 95, -54, 54, -16, -69, -102, 59, 79, 116, -72, 6, -78, -52, -35, -54, 6, -50, -12, -25, -42, -78, 119, -15, -70, -35, 74, 58, -41, -115, 49, 74, -29, 72, 119, -25, -58, 45, -52, 109, 86, 41, -49, -97, -115, 75, -76, -56, -20, 113, 22, -60, 121, -19, -29, 105, -14, -28, 48, -38, 36, 19, -14, 110, 45, 47, 33, 57, 86, -74, -21, -34, -10, -23, -112, 74, -115, 13, -102, -14, -127, 8, -65, 42, 81, 109, -35, 106, -9, 105, 74, -115, 52, 62, 17, -46, -45, -71, 20, 76, 52, -110, -123, 61, -21, -13, -76, 14, 1, -128, 109, 58, -64, -111, -71, 70, -115, 43, -38, -79, 49, 125, -49, -55, 121, -90, 59, 48, -9, -127, -37, 61, 49, 31, 79, 115, -86, -62, -71, -112, 32, 65, -68, -107, 39, 60, -86, -113, -51, -34, 115, 19, 83, 90, -87, -24, -81, -119, 115, 21, -91, -123, -102, -38, -115, -69, 2, 86, 6, 109, 25, 93, 38, 120, 50, 39, -119, 30, -45, -8, -125, -74, 8, -119, 11, 15, -41, -55, 49, -42, 15, -119, 111, -4, -84, -70, -123, 59, -2, -51, -102, -12, 39, -116, 29, -6, 121, -38, -59, -52, -50, 80, -13, -52, 52, -34, -81, -127, 38, 78, -97, 13, -55, -58, -85, -80, -24, 19, 50, 75, 73, 22, -49, -78, 84, -103, -48, -56, -88, 90, -95, 6, 67, -47, -7, 17, 118, -98, 119, 30, 109, 88, -101, -25, -110, 45, 39, -76, 43, 26, 46, 55, 48, -106, 95, 29, 11, -108, -15, 104, 101, -1, 122, -101, -115, -37, -128, 47, -41, -78, 112, 122, -83, -58, -76, -85, 98, 88, 31, 92, -118, 61, 12, 119, 9, 34, -15, -76, -119, 123, 36, -72, 122, 97, -58, 97, -40, 90, 12, 23, -2, 47, 88, -81, -8, -11, 44, 23, 89, 77, -52, 120, -75, 125, -100, -67, -108, -65, 79, 104, -95, -30, -113, 20, -19, -35, -25, -72, 65, -8, 111, -113, 32, 32, -84, -112, -56, -96, -11, -42, 59, -36, 127, -18, 6, 30, -128, 123, -85, -50, 33, -86, -35, -25, -77, 28, 90, 84, -69, -64, 35, 65, -90, -7, 71, 8, -105, -120, -86, 0, -69, -78, 46, -11, 79, 70, 49, 20, -1, -47, -73, 124, -121, -123, 95, 123, 101, -62, -11, 118, 29, -16, -76, -53, -17, -46, 29, 82, 56, 87, 96, -47, -21, -34, -67, 95, -12, 49, 23, 10, 113, 98, 6, 13, 22, -93, -74, 30, 118, -94, -2, 38, -60, -28, -3, 83, -25, 70, -121, 41, 100, 118, -95, 6, 35, 72, -98, -30, 13, 5, -40, -59, -23, 5, 27, 123, 60, -67, -94, 13, -71, 96, 30, -127, 46, 77, 124, -122, 3, 26, 120, -6, 37, 119, 59, -110, -11, -50, 120, -120, -5, -101, 36, 32, -1, 7, -81, 11, -122, -91, 47, 84, -40, 127, -87, 107, -4, -35, 108, -61, 10, 124, 18, -11, 29, 56, -124, -127, -42, -57, -110, -16, 20, 5, -28, -123, 67, -12, 97, -30, 124, 125, -60, -18, -117, 52, 73, 102, 64, 97, -85, 126, -31, 13, 32, 114, -44, 67, 4, 72, 67, 92, -52, 62, 23, -63, -84, 115, 68, 44, -113, -5, -64, -87, 56, -90, -15, -86, 5, -9, -2, -110, -19, 22, -4, 89, 43, 104, -73, -48, 126, -94, 77, 37, -59, -77, -66, 113, 97, 56, -127, 67, 36, -106, 15, 37, 77, 115, 124, 98, 70, 7, 0, -34, 93, -25, -64, -41, 18, 105, -127, 75, 56, 44, 9, 49, 83, -8, -22, 127, 69, -48, -108, -123, -101, 25, -17, 27, 74, 71, -39, -92, 108, 92, 12, -15, 41, 55, 38, -51, 122, 23, -21, -112, -68, 101, -36, -7, -127, -62, 127, 89, -37, 95, -105, -46, 26, 23, -108, -72, -95, -46, -96, -41, -28, -76, 22, 62, -70, -72, 90, -70, -52, 93, -55, 123, -53, -57, -28, 109, -117, 89, -62, 120, 59, 29, -6, -18, -116, 101, 8, 35, -89, -41, 33, -68, 19, 16, 114, -88, -57, -101, 18, 64, 117, -74, -10, -60, 107, 96, -72, -14, -7, 46, -38, -67, -109, -51, 118, -103, 14, 69, -59, 36, -87, 110, -109, 14, 62, 33, -97, 16, 21, -80, -79, -56, -128, 77, 99, -4, 105, -20, 95, -12, 88, 95, -117, -51, 23, 117, 85, -70, -78, 113, 104, -9, 10, -25, 108, -27, 23, -13, -63, 56, 24, -28, 11, -127, -54, -59, -100, -41, -46, 118, 1, 73, -9, 15, 61, 2, 37, 76, -120, 127, 121, 48, -34, 104, -79, -71, 118, -97, -8, 70, -100, -96, 0, -7, -17, 89, -123, 34, -118, -70, -103, 2, 39, -77, 90, 38, -24, 79, -13, 117, 91, -91, -53, -17, -5, -47, -7, -112, 60, -105, -87, 66, -7, 3, 63, 11, 38, -7, 86, 12, 71, -83, -55, -4, -104, -116, 38, -47, -127, -59, 0, 92, 24, 68, -91, -111, 84, 37, -92, -123, -92, 71, -116, -94, -70, 101, 95, -113, -81, -116, -48, 76, 41, 20, -100, 18, -125, 87, 120, 15, 50, -13, -73, 68, -125, -109, -100, -91, -82, -13, 86, -119, 77, -31, -97, 71, -96, 84, 126, -37, -22, 69, -59, 80, 122, -48, 51, -76, 59, 82, 37, -52, -84, 8, -10, -45, -128, -23, 75, -93, -47, 34, 3, 31, -34, 0, 32, -128, -25, 32, 61, -19, 42, 50, -41, 94, -93, 126, -22, 54, -55, 59, 79, -113, 89, -53, -85, 105, -25, 7, -76, -110, 101, 105, -125, 67, -128, -60, -111, 100, 53, -68, 111, -54, 113, 2, -28, -34, -96, 62, -46, 87, 78, 117, 76, -57, 7, 4, 80, -53, 123, 97, -114, 14, 97, -80, 56, 37, 48, -99, -22, 18, 109, 61, 104, -13, -44, 33, -32, -67, 105, 103, 43, -80, -49, -97, 72, 24, -79, -121, -63, -105, -13, 36, 107, -71, -99, -74, 101, 48, -60, 28, 4, -51, 3, -65, -97, 72, 11, -34, 30, -108, -68, 85, 17, -86, -65, 81, -42, -66, 52, 42, 99, -6, 39, -96, 49, -79, -2, -17, 29, -116, 72, -93, -14, 41, -76, 63, 87, 55, 16, -106, -57, -2, 12, 40, 47, -117, 58, 99, -118, -111, 92, -82, -49, 116, 115, -85, 110, -82, 40, 4, 57, 74, -93, -40, -56, -114, -96, 60, -14, 126, -13, -31, 51, -12, -107, 96, 55, 108, 96, -35, 77, 127, -63, -71, 96, 23, -107, -12, -52, -19, -67, -5, 105, 121, 60, -126, -95, -16, 70, 45, 54, -107, 7, -10, -124, 12, -121, -110, -95, 38, 31, -8, 48, 31, -75, -26, -123, -40, -33, 12, -127, -75, 80, 121, -20, -42, -70, -120, -72, -87, -36, 62, 87, 100, 82, 10, -96, -22, 102, 0, 63, 6, 81, -5, 89, -106, -47, -31, 82, -32, -72, -103, 76, 102, 59, 28, -47, 63, 118, 92, -30, -61, -74, 77, -43, -112, 41, -37, -50, -43, 111, 20, -98, 103, 15, -101, -54, 124, -126, -95, 67, -77, 14, 110, 22, -104, -65, -81, 117, -65, -34, -119, 49, 9, 62, 9, 19, 90, 24, -106, -13, -49, -93, -9, 84, -70, -116, 110, 53, 0, -40, 3, 42, -33, -52, 119, -71, 70, -78, -50, 25, -34, 110, 107, -103, 20, 32, -56, 90, -77, 11, 74, -18, -76, -17, -122, -114, 9, -96, 4, -118, 121, 37, -51, 71, 52, 75, 31, 30, -101, -90, 112, -37, 102, 59, -20, 41, 97, -50, -82, 13, -11, -95, 19, 67, 47, 118, 86, 103, 56, -8, -12, 71, 47, -23, -43, 100, -75, 107, 101, -98, 80, -38, 12, -124, 77, 26, 105, -40, -101, -124, 46, 96, -121, 90, -36, 113, 117, 125, 109, 107, 100, 66, 17, 31, 47, 83, -32, -51, 89, 70, -62, 33, -32, -7, 12, 31, 19, 6, 115, 100, -91, 37, -20, -38, -101, -51, -113, 69, -80, -35, 122, -66, 116, 90, -73, -61, -59, -62, 86, -67, -65, 37, 72, 109, -41, 65, -20, 12, -87, -41, -82, -36, -99, -43, -121, 19, 64, -101, 0, 59, 42, 77, -111, -60, 17, -52, 85, 78, -120, -52, -52, -35, -97, 112, -88, -106, 87, -7, -20, 52, 71, 27, 105, 89, 27, -26, -39, 30, -89, -55, 109, -30, -38, 119, 44, -16, 34, -26, -94, -13, -112, 116, 13, 29, 107, -98, -88, -1, -70, 92, 104, -89, -86, 56, -22, 122, 62, -5, 119, 67, -49, 115, 4, -109, 45, -27, -97, 5, -73, -117, 126, 120, 43, -59, -108, -11, -86, 38, -36, 25, -67, 11, 126, 65, -64, 48, -114, 1, 95, -81, 46, -45, -1, -124, 67, 55, -112, -46, -28, -62, 51, -94, 32, -6, -73, 95, 119, -120, -42, -90, 61, -117, -91, 61, 106, -128, 90, -72, -25, -41, 51, 59, 74, 111, 30, 127, 51, 35, 62, -10, -68, -117, -114, -121, -95, 47, 46, -71, -46, 93, -101, -93, 36, -55, -102, -99, -102, -120, 2, 75, -107, 45, -98, 10, 83, -104, -32, 39, 65, -17, 42, -114, 100, -112, 8, 89, 39, -57, 67, 79, -94, -69, -1, -77, -30, 16, 112, 55, -74, 126, 76, 85, -58, -4, 22, -72, 58, -42, -95, 8, -6, -105, -89, 32, 104, -109, 110, 8, -45, 96, 64, -100, -36, -86, -115, -37, 119, 2, -19, -106, 98, -89, -55, 62, 82, -44, 18, 69, 103, -100, 100, 39, -63, -97, -56, -118, -65, -29, 33, -113, -35, -104, -37, -99, -59, -83, 32, 88, 51, -89, -20, 75, 124, -119, 5, 124, 72, -76, -74, -91, 106, -58, -43, -97, -127, 75, -19, -47, -81, 77, -9, -125, -21, 80, -102, -120, 96, -81, -83, 72, 64, 19, 67, -51, -57, 106, -97, 112, 91, 62, 28, -5, 98, -63, -54, -115, 104, 111, 21, -54, -102, 26, 60, 95, 56, -43, 97, -4, 121, 76, 111, 111, 48, 29, -16, 108, 27, -48, -23, -111, -44, 11, -96, 45, -53, 36, -73, 1, 90, 5, 73, 44, -42, -126, 2, -31, -81, 12, -62, 64, 98, 85, -51, -26, 62, -13, -58, -37, -70, -7, -89, 10, -109, 91, 70, 116, 68, 17, 90, 99, -56, -17, 54, -42, -100, 85, 35, -10, 120, -117, 6, 32, 122, 126, -98, 22, 89, -81, 23, 58, 104, -126, 38, -59, 111, -52, 116, -116, 99, 35, -77, -10, -61, 102, -71, -39, 89, 85, 120, -70, 123, -99, -26, 68, 53, -68, 63, 9, 85, -45, 16, -17, -127, 122, -13, -4, -27, -54, 9, 67, -110, -9, 88, 62, -88, -16, 80, -20, 119, 110, -9, 49, 20, -31, -31, -12, 127, 30, 14, 18, -126, -50, -97, -92, 22, 52, -97, -101, 84, -49, 84, -37, -90, 45, -8, -42, -105, -80, -118, 5, 97, 39, 121, -34, 80, 24, 63, 23, 64, -50, 67, -117, -70, 76, 72, 17, -127, -114, 63, 116, -39, -43, -95, -113, -101, -85, 90, -10, 103, -44, -8, -9, 124, 71, 73, -60, 77, -83, 0, 104, 116, 81, -46, 8, 86, 44, -105, 15, 53, -63, -12, 14, 64, 111, -29, -43, -76, -78, -54, 97, 30, 90, -32, -6, 120, 119, -92, 22, 62, -95, 46, -55, 81, -16, -27, 53, 60, 86, -53, 107, -123, 33, -122, -123, -77, -98, 76, 5, -63, -109, -119, -106, -121, 120, -86, -9, 122, 51, -14, -32, -67, -39, -94, -6, -124, 87, 81, 42, -94, -36, 78, 109, 6, -121, -89, 109, -29, 8, 77, 104, 104, -13, -83, 89, -7, 4, 52, 17, -128, 76, -71, 48, -43, -100, 93, -43, -22, 76, -109, 100, -13, 64, -8, 92, -21, -109, -71, -124, -105, 19, 74, -117, -93, -97, -125, 96, -95, -122, -8, 118, 73, -47, 64, 59, -36, 40, 83, 50, -51, -16, -31, 49, 70, 33, -112, 85, 29, 26, -2, 7, -67, -122, 34, 88, -12, -65, -100, -1, -118, -112, -3, -37, -51, 35, 66, -11, -34, 19, 93, 47, -94, 61, 64, -92, 84, -75, 25, 90, -126, 60, -86, 60, 71, -42, -92, 73, 114, 66, -69, -17, -46, -67, -69, -45, 104, 72, -34, 33, -54, 104, -2, 62, 105, -76, 60, 114, 108, 45, -102, 22, 20, 34, -22, 79, 27, -82, 54, -52, 77, -119, -118, 88, -1, -85, 59, 24, 84, 52, 116, 6, -85, 68, -78, 112, -41, 34, 22, -62, -18, -103, -125, -73, -55, -15, -28, -3, -23, 52, 118, -114, 14, 69, 41, 12, -59, 78, -64, 86, 107, -118, 71, 75, -37, -57, -31, -107, -60, -17, -108, 31, 78, 91, -53, 112, -52, 86, -127, -81, 85, 81, -80, 62, 13, 7, -20, 38, -11, 75, -117, 7, -102, 94, 60, 8, -70, 1, -70, -93, 96, -35, 87, -26, -81, -14, -54, -67, -95, -32, 10, -124, 55, -19, 117, 79, 78, -107, 114, 4, -38, -107, -54, 85, 53, 97, 22, 5, -58, -95, 2, -40, -92, -124, -3, -128, 125, 55, -119, -110, -94, -90, -53, -116, -24, -2, 39, -35, 69, 5, 126, 85, 8, -38, -24, -84, 7, -109, -117, -16, -8, -51, 91, 18, 28, -16, 97, -109, -72, -15, 74, 76, 64, 36, 52, -122, -117, 49, -108, -102, 34, -66, -117, -41, -75, -36, 3, -99, -117, 79, -96, 65, 23, -95, -6, -42, 28, 13, 29, -95, -1, -20, 78, -91, -116, -66, -8, 82, 103, 105, -119, -59, 116, -98, 88, -1, -23, -51, -123, 99, 5, 33, 79, 50, -83, -84, -109, 123, -78, 29, 109, 34, 102, -62, 115, -34, 16, 32, 13, 40, 114, 23, -27, 96, -27, 22, 103, -68, -38, 49, -41, -81, -60, -43, 9, 25, 12, 75, 41, -75, -126, -30, -81, 8, -10, 77, 88, -116, -52, -57, -72, -105, 5, -84, 13, 3, -96, -100, -32, -4, 22, 44, -52, 48, -6, 30, 19, 75, -94, -94, -104, -46, -36, -87, -66, 59, -125, -34, 76, 34, 56, 67, 76, -64, 101, -75, 116, 20, 126, -88, -124, 43, 45, -3, -88, -6, 115, 75, -61, 56, -96, -44, -31, -60, 113, 84, -6, -127, -93, -81, -77, -52, 29, -35, 30, -40, -106, -6, 101, -115, -42, -21, 98, 126, 69, 47, 12, 72, -34, -89, 16, 88, -80, 58, -58, 31, -37, 122, 7, 98, 72, 104, -117, -66, 108, -4, 78, 49, 18, 51, -106, 117, -103, 110, -79, 93, 2, -99, -85, 93, 29, -109, -111, 56, 91, -48, 119, 58, -55, -58, 110, 46, 127, -66, 106, -9, 69, 0, -95, -35, 52, -79, 13, -14, 77, -13, -30, -30, 127, -107, 57, -52, 58, 67, -32, -57, 76, -46, -66, 92, -104, -99, 63, 53, -58, -50, -118, 54, -48, 27, 124, 36, -84, -111, -112, -22, -56, 120, -113, -102, -4, -44, -26, 49, 116, -107, 118, -26, -67, -87, -66, -68, 106, 88, -37, -57, -116, -76, 69, 28, 113, -107, -7, 103, 29, 94, 58, -94, 115, 25, 93, 3, 87, -20, -58, 79, 125, 110, -46, -72, 68, -99, 49, 40, 33, -108, 56, -81, 112, 29, -104, 7, -70, -34, -22, -60, -46, -2, 96, -125, 50, 110, -12, 8, 48, 112, 17, 109, -82, -66, -108, -124, -49, 73, 3, -14, -103, 110, 73, 39, 85, -45, -40, -7, -105, -116, 112, -49, -78, 63, 93, -49, 127, 33, -40, 71, 81, -119, 11, 26, -93, 71, -7, -26, -6, 71, 104, 116, -105, -43, -99, 61, -14, -98, 35, 102, -97, 89, -113, -48, 75, -110, 97, -11, -100, -104, -61, 40, 49, 34, -39, -97, -21, -28, 10, 127, 26, -61, -46, -20, 37, -108, 72, 10, 5, -49, 21, 2, -124, 21, 54, -111, -10, -42, -67, -93, 59, 33, -24, 107, -67, 108, 18, -72, -106, 71, -21, 73, 56, 78, -36, 70, 19, -99, -69, 9, 64, -17, 16, 43, -55, 89, 55, 117, -112, -29, 119, -105, 51, 15, 65, 28, 91, -74, 77, 94, 41, -90, -52, 117, 74, 74, -115, 62, -10, 28, -47, 82, 37, 114, 40, 35, 83, 106, 95, -65, -43, 101, -28, 95, -60, -69, -4, -25, 47, 9, -79, -100, 76, 74, 104, -72, -77, -65, -9, -10, 89, 64, -37, 48, -96, 16, 91, 14, 76, 42, 20, 124, 1, 98, 29, 84, 81, 43, -46, -88, -10, -50, -95, 48, 90, 59, 55, 70, -42, 18, -71, -40, 105, 121, -20, 26, -55, 118, 81, -113, -25, 37, -22, -10, 0, -64, -42, -22, -36, 120, -114, 70, -5, 92, -50, 35, 105, 117, 85, -47, -20, -57, 9, 52, -96, -100, 90, -117, -89, -73, 15, 6, 60, 89, 54, 127, 115, 112, -93, -58, -7, 64, 111, 116, 115, 101, 32, 125, 36, 63, -84, 68, 101, -124, 104, 20, -47, 57, 66, -32, -112, -77, -63, 2, 123, -75, 92, -8, 42, 83, -59, -15, -70, 41, -113, 33, 104, 42, -9, -65, 78, 92, 124, 64, 48, 94, -27, -63, 10, 82, 45, -105, 59, 99, 38, -63, -7, 99, 93, 38, 94, 95, 74, 59, -74, 67, 106, -70, -13, -39, 93, -22, 32, -96, -61, -123, 89, 85, 120, 118, 31, 95, 44, 53, 72, 40, -76, -111, -71, 53, -7, 62, -97, 77, 68, 11, -125, 25, 55, -63, -50, 109, 121, 122, 15, 26, 62, -100, 122, 127, 40, 86, 79, -50, 5, 31, 98, -35, 10, 6, -63, 43, -124, -77, -53, -105, -98, -70, -7, 26, -27, -64, 23, -9, -78, -7, -89, -80, 48, 12, -24, 37, -69, 112, 88, -47, 24, -14, -45, 79, -99, -74, -120, -73, 94, 24, 33, -17, 87, 61, -70, 54, 114, -32, -41, -86, 36, -109, -42, -107, 118, -47, 102, -88, -104, 56, 24, 21, 8, 76, 33, -84, 107, 74, 95, 85, -22, -76, 18, -82, 73, -14, 18, -52, -90, -67, -75, 46, -17, 60, 119, -5, -97, -37, 29, -82, 118, 122, 51, 37, -97, 63, -124, 26, -104, -4, -39, -111, -77, 81, 89, 91, 33, 73, 110, -70, 122, -102, 17, -109, -89, -4, 85, -12, 52, 40, -91, 101, -100, 61, 77, 7, 84, -11, -100, 21, -98, -36, -128, 60, -87, 26, 42, 32, -116, -69, 124, -79, -86, 99, -101, -51, 108, -88, 37, -119, -114, 39, 55, -57, 94, -105, 54, 109, 114, -16, -78, 12, 12, 37, -3, 97, -72, -76, 66, 24, 98, 66, 119, 35, 31, -116, 14, 104, 106, -35, -71, 6, -91, 85, 127, 126, -120, -27, 12, 56, -34, 77, -60, 70, -57, -15, 5, -48, 65, -76, 101, 99, 96, -65, -68, -87, 85, 15, -34, 106, -51, 44, -111, -111, -16, -119, 88, 95, 76, -112, -49, -19, 7, -39, -66, 121, 113, -25, -108, 86, 89, -21, -82, -126, -21, -27, 8, -37, -123, -64, -49, -30, 92, 78, 43, -116, -95, 81, 75, -114, -24, -72, -73, 107, -44, -49, 121, -22, 91, 100, -103, 117, -105, -16, 30, -72, -127, 122, 28, 76, 30, 62, 33, -27, 69, 79, 16, 9, -117, -23, -44, -123, -106, -115, 89, 50, -124, 104, -59, -26, -91, -124, 53, 31, 103, 14, 20, -103, 80, -79, 7, 122, 119, -126, 73, -71, -105, -10, 107, 67, 14, -111, -77, 100, -88, -16, -114, 118, 65, -32, -50, -68, 37, 118, -96, -103, -59, -2, -104, -128, -103, 104, -103, -100, -111, -59, -3, -13, -81, 17, -36, 14, -74, -40, -121, -15, -43, 28, 86, 53, 35, 53, 92, -108, 67, -77, -91, -79, -77, 29, 64, 30, -86, -28, 124, 19, -53, -54, -67, 94, -8, -18, 41, -87, -16, 114, 92, 70, 126, 37, -19, 60, -119, -36, -50, 27, 5, -82, 78, 97, -5, 13, -96, 84, 47, -21, -26, 125, -72, 29, 99, 97, -35, 11, 69, 77, -13, 10, 3, 54, -89, 43, 30, 117, 103, -20, -23, 67, 14, 65, -38, 72, -60, 73, 60, -23, 92, 19, 17, -63, 101, 42, -121, -121, 11, 46, 94, -20, 82, -42, 3, -90, -111, 39, -56, -17, 80, -71, 96, 6, 92, -99, 25, -20, 61, -25, 44, 107, -54, 114, 41, 34, 70, 45, 117, 127, -45, -4, 105, 3, 74, -1, -85, 24, 55, -4, 79, 101, -29, 10, 69, -113, -45, 104, -65, 51, -81, -48, -45, -78, -105, -18, 73, 11, 118, 73, -28, 18, 100, 28, 41, 47, -56, 64, 14, 100, 42, -89, -34, -17, -31, -42, -99, -85, 54, 29, -19, 15, -60, -122, 66, -29, 22, 34, -6, 5, -17, -42, -26, 80, 125, -60, 8, -92, 73, 121, 17, 60, 22, 93, 18, 40, -54, 19, -42, 103, -93, 41, 25, 37, -60, 57, -88, -99, 3, 55, -128, -16, -27, -120, -101, 47, 63, -14, 115, 39, -91, -69, 1, 100, -3, -58, 102, 103, -126, 126, 40, 11, 110, 115, 33, 47, -51, 27, -83, -127, -60, 16, -80, -46, 71, -54, 3, -96, -109, 69, -8, 53, 127, -5, 41, 33, 66, -75, 21, -48, 91, -108, 116, -9, -93, -34, -76, 64, 5, -101, 53, 88, 68, -61, 0, 84, 95, 25, 83, -1, 54, 88, -47, 100, -71, -87, 64, 65, 52, 66, 55, -24, -98, -38, -104, 76, -78, 55, 127, 117, 39, -87, 33, 82, -106, 41, -96, 3, 78, 112, -43, -28, -9, -122, 15, -82, -112, 117, 79, -64, 113, 97, -4, -39, 91, -99, -47, 11, 33, -43, -118, -107, 63, -8, -100, 86, 67, -47, 25, 74, -35, -94, 77, 52, -89, 76, 115, 26, 47, 77, -127, -108, 9, 126, -84, -58, 91, -55, -128, 83, 66, 75, -74, -119, -105, -25, -7, -69, 62, -125, 106, -112, 41, 4, -103, 50, 76, -98, 26, -84, -25, 39, -1, -84, -95, -46, -107, -92, -42, 100, 45, -109, -51, -68, 24, 14, 85, -60, -41, 93, -95, -105, -60, 54, -46, -116, -79, 50, -55, 114, 90, 67, -50, -121, -14, 88, -32, 59, 14, 108, -62, 59, 106, 3, 34, 35, -28, 49, 21, -51, 46, -10, -47, 35, -90, 58, 40, -18, 70, -80, -30, 97, -77, 77, 126, -34, -12, 43, -33, -116, 107, 47, -74, -80, 25, 65, -23, 58, -88, 54, 97, 69, 65, 22, 25, 18, -89, 125, 69, -17, 17, 101, -33, -41, 82, 23, -18, -104, -23, -14, -73, 17, 59, 92, 23, 80, -109, 33, -29, 84, -88, 23, 110, 96, -82, -28, -21, -1, -55, 39, -42, 111, -13, 63, 12, -107, 38, 78, 65, 91, -73, 110, 127, -57, -63, -59, -62, 108, -65, -105, 71, 4, 115, -116, 92, -100, -106, 103, -2, 60, 31, -25, -94, 81, -118, 75, 99, -18, -36, 70, 93, 63, 38, -109, 74, 94, 83, 61, -9, -107, -6, 14, 82, -65, -72, 8, -36, -100, 116, 81, -72, 68, 35, -11, -60, 108, -116, 54, -48, 124, -120, -12, 19, -126, -105, 84, 47, 73, 115, 39, 105, -22, -44, -86, 85, 89, 57, 39, 13, 82, -52, 94, -106, -93, -86, 68, 71, 10, 95, 85, 112, 107, 91, 64, 52, -101, -34, -26, 126, 49, 43, 122, 37, 55, 25, -128, -46, -100, -51, 44, 47, -58, 92, 17, 99, -88, -111, -51, -66, 41, 93, -9, -104, -119, 45, -36, -124, 110, -84, -10, 100, 116, -15, 20, -2, 18, 75, -74, 107, -89, 12, 125, 18, 92, 58, 23, 47, 70, 9, 60, -34, 21, -12, -105, 11, 99, 95, -27, -105, -99, -91, 66, 3, -88, -64, 94, 7, 61, -89, 16, -59, 60, 11, 37, -37, 82, 17, 15, 46, -14, 31, 33, -99, -94, 14, -91, 118, -108, -34, 13, 61, -20, 55, -97, 59, 66, -3, 8, 55, 67, 7, 119, 104, -121, -102, -13, -113, 17, -52, 25, -44, -123, -30, -67, 86, -80, 27, 121, -101, 6, 84, -11, -25, -113, -92, -80, 22, 26, -46, -21, 54, 13, -45, -18, -95, 47, 106, -81, 118, 35, 74, 88, 87, 17, 36, 39, 55, -33, -68, -50, 103, -103, -24, 123, -78, 114, 71, -36, 79, 35, -72, -62, -57, 18, 91, -43, -122, -46, -77, 27, 105, -6, 99, -42, -3, -94, 31, -65, 41, 27, -66, -127, -91, 10, 3, -65, 17, 68, -3, 85, 5, -1, -73, -97, 99, -62, -105, 17, 25, -81, -46, -110, -102, 86, 27, -34, -50, 124, -85, 52, -62, 51, -27, -24, -79, 19, -88, -44, 58, -111, 104, 116, -6, -29, 72, -94, 52, 84, -5, -71, 10, -119, -91, -11, 60, 74, 53, -27, 39, 106, -114, -91, -46, 67, -103, -127, 53, -78, -114, -103, 96, 90, 59, -86, -21, 41, 91, 67, 73, 58, -39, -80, 2, -38, 10, 11, -107, 58, -107, -50, -32, 126, -123, 95, -18, -37, -75, -28, -73, 37, 8, 64, 21, -37, 14, -32, -9, -28, -48, 14, -91, -30, 117, 47, -44, -87, -37, -21, -49, 99, -14, 37, -30, -87, -96, -32, -115, -83, 15, -42, 127, 101, 9, 57, 31, -29, 19, 52, -42, -89, -92, 70, 118, -42, 33, -90, -68, 104, -90, 94, -105, -38, 48, 57, 90, -31, 84, 67, 19, 78, 33, -18, -114, -69, 101, 113, 24, 5, 102, -26, -100, 117, 27, -113, -80, 73, -40, -60, 69, 120, -78, -23, -114, -9, -68, -123, 76, 39, -116, 41, -120, 119, -24, -2, -13, -28, -6, 70, -95, -122, -17, -117, 66, 19, -67, 99, -80, -69, -6, -20, -15, 43, 33, -32, 112, -25, -31, 84, 15, -96, -80, -60, 81, 26, -40, -58, -19, 20, 65, -57, 46, 46, -114, 73, 88, -96, -67, -19, -70, 54, 76, -107, -29, 97, -121, 113, -57, -69, 24, -67, -19, 55, -40, -29, 28, -112, 53, -89, 116, -21, -34, -50, -118, 65, -27, -89, 43, -102, 77, 117, 104, 102, 61, -101, 18, -74, -67, 31, 116, -89, 116, -62, -36, -38, 84, 111, 110, 90, 104, -104, 70, -92, 17, 54, 82, -70, 64, 82, -122, -38, 23, -15, -36, 36, 81, 122, 26, -7, 104, 108, -42, 12, -41, 32, 33, -104, 68, -95, -109, 32, 119, -20, 99, -70, 70, -45, 10, 80, 72, -14, 111, 44, 46, -74, -36, 119, 56, -38, 90, 75, -116, 99, -125, -54, 81, 41, -102, 60, 15, 67, -31, -94, 122, -17, 121, -8, -23, -42, -118, 111, -110, -118, -73, -47, 120, -79, -81, 64, 9, -62, 76, -59, -6, -60, -113, 19, -44, 2, -97, -80, -48, -84, -32, 38, -107, -75, -112, -98, -28, -3, 123, -112, -5, 79, 72, 97, 80, 65, -105, -18, -61, 44, -16, 75, -67, -2, -83, 13, -38, 122, -4, 73, -11, 76, -15, 27, 59, -82, 116, -48, -12, -111, 81, -27, 124, 106, -73, -110, 9, 74, -119, -95, -91, -42, 69, 61, -89, 80, 29, 95, -84, 83, -124, 112, -90, 43, -92, 68, -48, -94, 93, -13, 72, 6, 88, 112, -93, 58, 68, 2, 41, 47, -41, -13, 48, -6, -70, -48, -17, 6, 26, 113, -6, -113, -18, 0, 48, -19, -53, -79, 11, 33, 49, -104, -72, 42, 37, -55, 73, -17, 48, -16, 26, -79, 50, 33, -48, 108, -126, 118, -18, -2, -122, -68, 24, 32, -103, 36, 79, 65, 45, 103, -23, -43, -41, -57, -25, -34, 13, -86, 120, 89, 105, 63, 125, -53, 56, 40, 123, -8, -87, 59, 123, -19, -7, -108, 86, -49, 75, 110, -6, 3, 6, -13, 91, 80, 34, 41, 18, -2, 31, 89, -93, -103, 9, 72, 81, -34, 14, -64, -79, 43, -75, -84, -20, 55, 9, 80, -102, -17, 87, -45, -66, -15, 108, -47, 39, 85, 118, 76, -105, 76, -124, 73, 82, -126, -86, 29, -7, 108, 122, 51, -35, 83, -49, -115, -71, -113, -56, -38, 95, 110, -102, -125, -53, -8, -117, 102, 117, -7, 60, -35, -38, 105, -79, -110, 42, 91, -72, -37, 62, -76, 45, -98, 47, -88, -12, -70, 42, 17, 33, 92, -78, -81, 21, 57, 126, 5, 13, 27, -19, 22, 21, -56, 31, 21, 73, -122, 57, 71, -67, -110, 28, 27, -71, 126, -81, 121, 24, 79, 66, -101, -29, -94, 89, 54, 45, -64, 103, 110, 83, 59, -103, -106, -94, 8, 71, 44, 91, 66, -91, -57, -117, 9, -3, 109, -20, 64, -45, 32, -84, 48, 11, -44, -20, -75, -113, 87, 109, 113, -108, 118, 23, 55, 13, -44, 39, -91, 74, -54, -88, 74, -46, 2, -68, 43, 5, 97, -103, -25, -15, -81, 61, -24, 113, 14, 118, -90, -72, 34, -57, 57, 44, -31, -7, -11, 37, -119, 46, -45, -16, -84, 30, 33, -111, -99, 119, 81, 109, 114, -56, 117, -77, -120, 118, 114, 3, 107, 80, -128, 23, 69, -69, -50, -128, 10, 116, -49, 90, -2, 18, 126, -78, -27, 64, -38, 44, -124, 57, -124, 123, 8, -87, -97, 23, -25, 101, 123, -50, 85, 25, -68, 77, -111, -110, -42, -65, 104, -101, 12, 100, 127, -95, -26, -23, 98, -62, -91, 10, -43, -62, 32, 123, 89, -128, -128, 12, -88, 121, 64, -64, -66, -83, 105, 54, 21, -88, 60, 14, -27, 83, 19, 25, -70, -95, 95, 56, -45, 127, 61, 114, -100, -34, 81, -38, -29, -65, 104, -23, -107, -19, -51, -15, -5, -91, -78, 39, -79, 29, 61, 5, -69, 31, -37, -96, -13, 32, 123, 72, -62, -22, 40, -128, 119, 11, -120, 118, -10, -15, 63, 76, -9, -8, -116, -108, -3, -100, -16, -74, -3, 87, 125, 7, 40, 98, 55, 85, 83, -99, 99, 16, 1, 39, 6, 110, -104, 112, 77, 80, 109, 53, 124, -31, -50, -24, 125, 111, -58, -80, 43, 5, -73, 107, -58, 27, -18, -67, -58, -108, 81, 21, -108, 52, -90, 24, -25, 10, -107, -109, -56, 60, 35, 97, -106, 121, -68, -21, -72, -104, -47, 11, 68, -15, -88, -47, -117, -61, 27, -110, 86, -126, 59, -99, -34, 126, -11, -97, 49, -107, 62, 4, -86, -104, -54, 50, -7, 66, -25, 41, 92, -5, -5, -73, 35, 57, 126, 51, -52, 24, -29, -10, 24, -90, 72, 2, -50, 27, 64, -33, -110, 100, 109, -121, -90, 15, -125, -45, 100, -92, -52, 37, 49, 86, 86, 125, 27, 49, 110, -122, 102, -100, 59, -17, 90, 94, 43, 37, 64, 56, 86, -104, 110, 5, 55, 6, -76, 117, 46, 62, -106, 123, -77, -2, -54, 105, 96, 86, -10, -21, -75, 25, -80, 34, 119, -77, 68, 34, -69, 59, -51, 23, 118, 95, 73, -114, -7, 64, 23, 17, -101, -63, 23, -119, -110, -51, 21, 122, -90, 122, 94, -6, -61, 15, -28, -106, 99, -78, 61, -11, -47, 120, -53, 116, -14, 125, -54, 36, -63, 101, 12, 19, -111, -96, 58, -69, 73, -39, -47, -56, 34, 30, 1, -62, 76, 52, 89, 45, -54, -108, -63, -86, 83, -54, 79, -50, -50, 76, 9, -4, 71, -39, 5, 4, -32, -71, 4, -93, 95, -63, -116, 7, 52, 50, -57, -31, 24, 127, -56, -25, 60, -115, -65, 124, 67, -60, -96, -51, 59, 90, 103, -48, -81, 22, 124, -41, 126, 40, 12, -19, -96, 101, -45, -33, 108, -27, -57, 126, -67, -62, -16, -122, -31, -70, -105, 115, -102, 103, -11, 9, 7, -17, 6, -27, 79, -22, -97, -103, 83, 35, 81, -124, -108, 115, -36, 69, 102, -102, 88, -104, 86, 93, -128, -29, -87, 18, -39, -114, -35, 10, 125, 63, 99, -25, 50, 41, 85, 11, -39, 61, -88, -123, 124, 123, 2, -33, -37, 85, 20, 37, 126, -73, 88, 12, 86, -39, 105, 23, 60, -98, 31, -128, 34, 77, -106, -94, -64, 37, -33, -61, -32, -3, 24, -115, -5, -56, -100, 125, -66, -103, -12, -6, 27, 73, 93, -4, -90, -128, 85, 98, -115, 85, 69, 102, 94, 18, 105, -13, 72, -51, 47, 86, -126, 106, 78, -51, 66, -113, -99, -112, -79, -13, -14, -107, -95, 8, -116, -3, 104, 118, -77, 23, 5, -92, 126, -75, 99, -55, 14, -45, 42, 93, 62, 6, -28, 10, 123, -127, -31, -78, -22, -110, 85, 17, 93, 58, -94, -96, -15, -31, -55, -2, 14, -59, -5, -107, 67, -41, 22, 47, -38, 74, -58, 50, 17, -54, 61, 49, 13, 127, 55, -110, -87, 21, 125, 121, 78, -89, -53, 91, 120, 70, 32, -35, -99, 110, 28, 101, -40, -53, -4, 127, 16, 56, -111, 42, 41, 28, 77, 32, -89, 16, 82, 51, -23, 29, -64, -86, -115, 99, 42, -61, 47, -103, -74, 123, 66, 58, -111, 62, -7, -34, 40, 44, -96, -122, 97, -15, 123, -43, -46, -59, 92, -74, -86, -111, 7, 56, 17, -90, -49, -7, 70, -48, -48, -16, -74, -78, 37, 36, 45, -52, -117, 71, 107, 119, -77, 127, 21, -24, -48, 98, 42, -55, 124, -122, 49, 58, 25, 106, 73, 59, -108, -61, 113, 63, -95, 85, -23, -78, -15, -83, 85, -123, -21, 109, 94, -36, 53, 120, 56, -66, 29, -82, 8, 62, -57, 126, 26, -35, 91, 60, 47, -49, 109, -123, 6, -128, 74, 75, -15, -32, 88, 18, -125, 42, -9, -115, 9, 31, 29, -46, -44, 0, -89, -4, 13, 103, -43, 115, 84, 28, 41, 37, -77, 21, -110, 117, 6, 38, -78, 45, 34, 37, -27, -93, -28, 69, 111, -19, -110, 31, -32, 124, 42, -65, -53, -94, -34, -47, 2, -116, 104, -117, 11, -120, -56, -42, 47, 36, -67, -78, 55, -60, -34, -39, -50, 16, 84, 36, 97, -118, 1, -42, 42, 42, 59, -92, 46, -126, -24, -126, -73, -82, 54, -39, 49, 52, -109, -36, -10, -108, -76, 5, 93, 25, 67, 118, 77, 119, -42, -91, 75, 99, 28, 51, -105, 70, 113, 0, -125, -37, 2, 18, -21, -15, -37, 33, -4, 0, 73, 28, 89, -17, -124, -52, 56, -101, -5, 29, -69, 29, 19, -67, 51, -121, -35, 55, -34, 31, 32, -13, 107, 65, 71, -34, -1, 12, -48, 49, -127, -54, -48, 73, 101, -48, -43, 123, 22, 103, -123, 49, -40, -66, -108, -74, 57, 107, -101, -82, -47, -108, 48, 118, -37, 70, -5, 0, 17, -49, -86, 43, 94, 55, 80, 114, 6, -30, -46, -39, -91, 38, 50, -51, 81, -59, -77, 76, -87, -44, -36, -41, 22, 127, 38, 107, 121, 21, -71, -95, -78, 82, -26, 16, 33, -83, -125, 63, 30, 96, 57, -53, 81, 47, 49, 78, -111, 14, -70, -34, 65, 118, -32, 89, -107, -106, -46, -78, 58, 123, -1, 99, -30, -24, -58, -107, 123, 87, -122, 34, -112, 2, -115, 18, 84, -111, 116, -8, -36, -52, 51, 7, 96, -61, 21, 9, 45, 54, 75, -34, -87, -116, 14, -43, -41, -99, -23, 8, 124, -16, 114, -6, -128, 65, 55, -64, 55, 91, -102, 58, -88, 30, -7, 47, 46, -8, -19, -84, -84, 126, -19, -38, 41, 100, 109, -43, 25, -69, -111, 85, -97, 38, 26, -23, -84, 16, -56, -123, 75, 124, 117, -79, 105, -7, -58, 0, 53, 114, 2, -25, 20, 53, 113, -75, -3, -108, 117, -15, -49, -90, 0, 32, 33, 53, -49, 105, -72, 74, -86, 122, 103, -111, 79, 81, 111, 60, -46, -9, 50, -15, 0, 10, 46, -45, 55, -51, 94, -87, 53, -48, 52, -100, 57, 30, -28, -63, 71, 96, -87, 12, -92, 123, 42, -88, 38, 17, -69, -36, 114, -99, 26, 16, -16, -56, -112, 64, 117, -101, -29, -33, -105, 101, 19, 80, 51, -14, -114, 67, -86, 34, -99, -73, -88, -62, -37, 127, -114, 99, -104, -92, -80, -66, 22, -126, -8, -54, 27, 59, 55, -66, 104, 125, 45, -79, 92, -100, -123, -40, 73, -60, 120, -42, 3, 109, 15, -101, 29, 108, -66, -34, -45, -116, -93, 41, 1, 77, -16, -18, 85, -1, 20, -59, -106, -7, -60, 69, 122, 31, 16, 7, -15, -56, -12, -91, 98, -42, 113, -82, -98, 65, 106, -22, 78, -67, 93, 81, 115, 78, -67, -128, 110, -102, -76, 22, 27, 106, -11, -113, 51, -6, -91, -127, -112, 44, -2, 38, 87, 11, 116, 121, -80, 20, -84, 41, -12, 30, 111, 50, 94, 53, 111, -96, 115, -19, 19, 39, 46, 13, 98, -67, 48, -43, 66, 71, 104, -47, 10, 108, -57, -17, -19, 117, 108, 114, -17, 25, 56, 42, -120, -123, 54, -59, 22, 11, 54, -10, -70, 32, 107, -57, -116, -34, 76, -28, 3, -64, -29, 119, -59, 65, 39, 101, -72, 28, 23, 3, 47, 15, 75, 9, 84, -21, -96, 98, 110, 74, 43, 107, 23, 66, 28, 13, 84, -67, -41, -117, 109, -111, -118, 64, 33, 11, 51, 67, 21, 11, -109, 124, 22, -36, 83, 56, 16, 31, -111, -22, 106, -108, -81, -106, -88, 120, -24, -4, -69, -54, -77, 59, 111, -67, -26, -50, 71, -56, -112, -5, -105, -30, 44, 123, 12, 2, -86, -60, 104, -88, 109, -127, 103, 100, -31, 92, 59, 63, -93, -78, 43, -97, 0, -52, -11, -13, 59, 18, 78, -112, 37, 19, -3, 79, 69, -31, 74, 22, 92, -57, -113, 114, -119, -80, 31, -92, 18, -106, 29, -36, -8, -36, 31, -5, 39, -68, 90, 90, 114, 98, 87, 117, -18, -95, 39, -71, 94, 75, -6, -80, -123, -18, -126, -91, -47, 3, 71, -15, -87, 112, -83, 33, -22, -75, -66, 105, 84, 0, 80, -127, 93, -26, -42, -82, -84, 20, 62, 7, -10, 97, -33, -99, 2, 100, -86, 49, 108, -6, 113, -26, -89, -70, -85, -100, 47, 99, -108, 11, -26, 111, 79, 45, -10, -41, 102, 13, -6, 93, -79, -15, 54, 11, -125, -1, 93, -92, -115, -83, -70, -64, -104, -16, -12, -34, -74, -99, 97, 36, -59, -108, 62, -35, -37, -42, 14, -64, 42, -16, 110, -15, 86, -111, -95, -49, 7, 123, -38, -33, -126, 79, 114, 107, -1, 89, -112, -15, -87, -69, 60, -101, -89, -115, 97, 89, -9, -121, -119, 48, 16, 4, -27, 101, 112, -74, -49, 104, -6, -122, -36, 89, 51, 65, -72, 115, -78, 92, -24, -64, -34, 126, -1, 114, -53, -114, -108, 90, 33, 59, -9, -115, 125, -3, -68, 88, 11, 46, -100, -17, 85, 59, 109, 88, 55, 68, -41, -1, 72, 85, 13, 7, 14, -84, -121, 101, 55, -49, 55, 100, -50, 75, 70, 42, -126, 82, -125, -37, 10, -56, 62, -21, -3, -123, -100, 39, -38, -49, 12, 56, -11, 91, -114, 14, 74, 110, 124, -82, 60, 14, 3, 88, -126, 45, -91, -35, 111, 100, -51, 81, 41, -76, 18, -50, 114, -7, -127, 98, -33, -53, 22, 96, -101, -13, 28, -42, -100, 21, 104, 28, 100, -18, 26, -37, -36, 13, 102, 75, -87, 47, -76, 122, -57, 73, -86, -77, 58, -35, 24, -10, 59, 22, 6, -47, -122, 45, -66, 68, -121, -94, 38, -12, -69, 9, 14, 59, -98, 66, 36, -70, 39, 116, 72, 99, -106, -5, -60, -36, 103, -122, -44, -87, -35, -119, 115, -74, -70, 40, -15, 79, 89, -26, -67, -9, -88, 104, -128, 46, 97, 86, 24, 101, -75, 30, 84, 43, 78, 32, 99, -5, 90, -62, 31, -125, 0, 113, -126, 92, -71, 85, -83, -51, -108, -8, 35, 0, 56, -13, 26, 102, -34, -82, 93, -66, -57, -10, -18, -89, -110, -119, 117, 121, 32, -71, 68, -101, -99, 8, -39, -115, 120, -123, -38, 119, -73, 112, -11, 100, -32, 112, -3, 10, 20, -9, -121, -6, -105, -41, -84, 6, -93, -29, 35, 6, -3, 117, 95, -71, -126, -24, 89, -110, -72, 45, 82, 91, 11, -74, -107, 101, 2, -63, -23, 119, -84, 26, -98, 7, -127, -25, 11, 56, 32, -62, 62, 31, -31, -112, 60, 57, -45, 16, 3, -71, 63, 121, -122, 95, 112, -90, 31, -33, -91, -31, -97, -73, -52, -22, -87, 5, 0, -96, 123, -112, -76, 45, -74, 15, 74, 106, -109, -128, -91, -54, -30, 92, 67, 94, 52, -111, 7, 26, 94, -48, -47, 53, 83, 23, 13, -97, -89, -44, -56, -115, 122, 6, -88, 3, -87, -71, -96, -78, -121, -118, -118, 81, -20, -82, 29, 24, -33, -73, -38, 76, 58, -36, 31, -37, 38, -63, -121, -13, 58, -42, -117, -107, -20, 119, -19, 50, -59, 95, -46, -38, 104, -43, -58, -111, 67, -56, -42, 7, 50, -89, 33, -96, -93, 35, 114, 119, -110, -75, -128, -128, 35, 114, -102, -22, 88, 26, 98, -122, 57, 12, -40, -101, 48, -61, 113, 16, -84, -36, -63, 104, -33, -44, 66, -124, 3, 86, 110, 104, -121, 40, -73, 3, 6, 98, 110, 50, -114, 29, -56, 111, -50, -43, -26, -72, 108, 99, -46, -14, -59, -16, -106, 98, 61, -111, -108, 1, 40, -13, 123, 106, -124, 59, 81, -94, 116, 107, -97, -8, -22, 89, 101, -16, -32, -102, 29, -71, 91, 0, -8, -79, -55, -68, 60, 114, -126, 21, 113, -110, -17, -121, -83, -18, 23, 46, 86, -54, 117, 10, 55, 77, -71, -67, -116, -104, 117, 15, -105, 8, 15, -108, -85, 115, 76, 53, 60, -109, 38, 19, -50, -112, 7, 8, 107, -110, -27, 9, -98, 126, 108, 72, -122, 44, 22, -73, -117, -20, 26, -85, 49, 83, 70, 72, 114, 85, -28, -6, 122, 49, -63, 38, 79, -83, 4, -86, 105, 21, -113, -70, 54, 60, 37, 101, -67, -48, 35, 37, 29, 110, 121, -18, -73, 80, -56, -29, 85, 85, 52, 17, -126, 32, -118, 73, -77, -23, -83, 27, 98, -97, 95, -63, 75, -92, -66, 18, -120, 109, -49, 73, 113, 52, -17, -12, -127, -31, -93, 77, 85, 57, 112, -88, 46, 102, 26, 84, 35, -120, -119, -105, 53, -14, 83, -110, 43, -94, -64, 75, -48, -30, -102, -39, -58, 80, -76, -82, 120, -93, -102, 85, -121, 12, -84, -10, -11, -49, 93, 104, -8, -17, 28, 39, -32, 100, 99, 80, 72, -44, 20, 37, 7, -22, -28, 109, 88, 52, 66, -80, -69, 30, 40, -11, -88, -101, 97, -39, 33, -23, 89, 29, 37, -60, -71, 12, 72, 31, -41, 121, -82, -48, -1, 76, -18, -39, -23, 60, 30, -118, -99, 43, 127, 50, -51, -65, -82, -128, -76, 63, 22, -43, 66, -14, 112, 10, 81, 10, -93, -30, -36, 70, -10, -25, 8, 24, -82, 72, 115, 38, 11, 69, -102, -75, -23, 34, -72, 24, 97, 66, -123, -16, 43, 80, -41, -63, -58, -76, -64, -100, 68, -68, 79, -78, -39, 16, -19, 102, -56, -121, -39, -121, -7, 27, -83, 103, -79, -17, 87, 24, 51, -108, 55, 39, 64, 54, -110, -12, -87, -22, -39, -116, -116, -17, 123, -26, -34, -18, 111, -14, 74, 17, 95, 68, 14, 78, 61, -12, 19, 36, 24, -87, -78, 11, 15, -13, 41, -21, -29, -38, 31, -44, 95, -77, -86, 120, 104, 68, 61, 1, -71, -75, -35, -14, 32, 75, 27, 65, 3, -26, -23, -2, 106, 83, 38, 59, -37, 32, -53, -99, -26, 39, -90, 10, 53, -67, 75, 127, 89, -43, 96, 113, -86, 22, 116, 16, -9, 90, -97, 88, 96, 8, -69, 97, -19, 74, 73, 12, 68, 84, -23, 98, -26, 126, 34, 83, -78, 20, 120, -10, 93, -126, -102, -84, -121, -34, 62, 19, -33, -70, 10, -46, -6, 36, 18, -7, -44, -69, 123, 21, -67, -7, 24, 38, -53, -17, -14, -22, 76, 124, 107, 114, -74, 62, 13, 93, -59, 19, 25, 17, 119, -76, 103, 6, 8, 94, 120, -30, -61, -66, 28, 82, 7, -98, 59, -122, 39, 60, -91, 10, -4, -2, 127, -88, -114, 64, -113, 60, 2, -31, 40, 80, 3, -102, 114, -95, -95, 77, -43, -72, -75, 39, 82, 60, -69, -74, 99, -69, -103, -66, -71, -96, -14, 37, 16, -10, 114, 61, -97 );
    signal scenario_output : scenario_type :=( 48, 32, 0, -41, 0, -4, 15, -23, -88, -54, -28, 23, 63, 61, -49, -22, -36, -30, 21, 39, 61, 43, 63, 53, 11, -41, -60, -68, -37, -32, -17, 79, 35, 14, 58, 17, -70, -61, 22, 11, -5, 47, 11, -27, 11, 78, -22, -14, -42, -73, 9, -13, 56, 54, -55, 48, 49, -31, 12, -6, -69, -100, 2, -41, -3, 70, 44, 90, 25, -42, -61, -25, 4, 61, 7, -38, 11, -11, 14, 57, -6, -21, -57, 36, 60, -9, 2, -21, -70, -28, -21, -21, -8, -11, 3, 5, 25, -22, -39, 29, 37, 65, 90, 70, -38, -74, -89, -68, -20, 23, -7, -10, 2, 18, 17, 8, 11, -28, -6, 45, 20, 72, 35, -3, -30, -45, -71, -36, 3, -21, 15, -4, 21, -63, 18, -36, -31, 55, -28, 37, 69, 39, 36, 30, -24, 0, 41, 30, 39, -2, -42, -57, -11, -14, -12, 42, -25, -38, 3, -28, 21, 89, -38, 4, 29, -3, 40, 0, -82, -62, -75, -13, 40, 27, 38, 9, -8, 13, -17, -10, 22, -12, 31, 12, 5, -3, -69, -43, -6, 54, 53, 31, 10, -18, -10, 19, 14, 30, 3, -4, 5, -46, -60, -30, -9, 54, -19, 39, 60, -15, 45, 71, -6, 14, 13, 21, -34, -55, -27, -39, -40, 46, 46, -24, 24, -74, -69, -5, -18, 25, 119, 20, -4, -37, -61, -42, -8, 80, -7, -20, 17, -34, 40, 15, 42, -20, -75, -36, 17, 60, 65, 80, -18, -117, -60, -41, 68, 49, 34, 23, -20, -79, -17, -46, -6, -22, 10, 43, 5, 45, 3, -2, 31, -55, -55, -14, -58, 8, 58, 47, 79, -25, -64, -1, 4, 51, 60, -10, -94, -60, -27, 10, 32, 40, -45, 40, -15, -31, 53, -11, 15, 83, -1, -55, -77, -62, -39, 10, 76, 70, -35, 10, 11, -68, -45, 26, -22, 22, 92, 51, 41, 49, -70, -63, -17, -75, -32, 60, -18, 29, 19, 65, -42, -39, -17, -53, 55, 60, 31, 27, 20, -2, 53, 15, -12, -4, -91, -24, 11, -37, 32, -1, -8, -28, 23, 60, 11, 36, -1, -73, -20, 0, -53, 6, -65, 5, 8, 13, 35, -12, -28, -29, 48, 14, 24, 10, 22, -88, -48, -13, -56, 3, 53, -8, 7, -26, 21, 29, -5, 38, -26, -31, 18, -27, 8, -18, -25, 30, 25, 29, 52, 21, 11, -1, -17, 26, -60, -27, -2, -27, 0, 12, 52, -81, 2, -11, -32, -3, -19, -9, -37, -21, -35, -7, 3, 74, 109, 40, 21, -36, -86, -35, 55, 48, 91, 66, 8, -60, -36, -52, -62, 5, -14, -20, 56, -4, 64, 31, 41, 59, 8, -21, -40, -30, -60, -8, 25, -13, 79, -25, -29, -35, -90, -11, 26, -5, -3, 58, 34, 49, 98, -26, -46, 11, -57, -10, -17, -5, -55, 6, 59, -6, 73, -12, -53, 5, -65, -37, 65, -23, -51, 22, -3, 24, 30, 41, -11, -91, 9, -6, -5, 87, 25, 54, 41, 3, 13, -22, -108, -72, -80, -68, 55, 103, 51, 22, -24, -48, -25, -40, 30, -51, 22, 70, 39, 79, -40, -68, -59, -62, 15, 48, 46, 44, 37, 30, -15, -6, -6, -47, 47, -4, -21, 4, 0, 27, 32, 8, -3, -32, -91, 18, -15, -24, 20, 78, 32, 29, 1, -48, -107, -63, 29, 59, 64, 38, 5, -7, -57, 11, -30, -4, -6, -34, 53, -60, 25, 10, -28, -20, 11, -34, -69, 3, -12, 41, 68, 85, 69, -35, -48, -29, -5, -40, 9, 18, -49, 40, 55, 26, 46, 24, -78, -69, -48, -29, 13, -1, 0, -3, 14, 51, 77, 20, -6, 18, -61, 0, -18, 24, -15, 11, -11, -30, -94, 1, 47, 27, 52, 34, -48, -6, 32, 36, 63, -2, -75, -13, -1, 11, 20, -10, 21, -18, 86, 64, -20, -53, -20, -57, 5, 37, -70, -17, -70, -49, 29, -12, 26, 109, 23, 38, 27, -37, 2, -15, 18, 49, -54, -1, -41, -53, 42, 7, 27, -17, 15, -14, 3, 2, -44, 20, 1, 20, 42, -31, -47, -32, 34, 20, 54, -12, -22, 3, -12, -23, 51, -4, -37, -44, -4, -56, -42, 62, -23, 4, 27, -15, 34, 56, -14, 34, -12, 30, -34, -39, -40, -39, -9, 34, 65, -5, 30, 4, -45, 13, 8, -29, 36, 27, 51, -44, -15, -21, -57, -30, 30, -13, 34, -28, 29, -27, 15, -21, 43, 36, -29, -58, -36, -26, 61, 79, 93, -3, -8, 29, -65, -5, 8, -59, 41, 69, 29, 7, -43, -2, -21, -15, 25, -7, -2, 3, 5, 14, -44, -59, -64, 10, 47, 25, 81, 82, -18, 51, 30, 14, -30, -64, -79, -54, -37, -35, 59, 54, -12, 47, -25, -31, 4, -9, -42, 26, -13, 31, 19, 26, -44, -27, -30, 0, 107, 4, 12, -2, -74, -41, 11, 46, 42, 85, -41, -68, -23, -56, 46, 86, 4, -8, 24, -22, 79, 41, -22, -54, -48, 19, 5, 41, -24, -58, -61, -17, 1, -5, -18, 19, -27, -4, 65, 14, 43, -30, -4, -12, -30, 20, -28, 52, -8, -55, 15, -31, 0, 9, 66, 83, 22, 42, 4, -25, -9, -80, -9, 26, -30, -1, -21, -72, -66, -20, 28, 76, 32, 35, -30, 21, -30, 30, 85, -52, -11, 1, 23, 0, 59, -26, -44, -55, -24, -21, 61, -29, -2, 49, 4, 47, 57, -37, -10, 12, -58, -20, 9, -30, -6, -29, 54, 7, -30, 76, -37, -82, -8, -17, 34, 38, 45, 8, 1, 40, 63, 56, 25, -4, -57, -73, 13, -54, 4, 52, -94, -54, -3, -38, 31, 79, -34, 43, -28, -74, 82, 19, 11, 55, 59, -55, -55, -27, -78, -26, 74, 0, 54, 80, 27, 68, 53, 4, -40, -76, -93, -15, -54, -73, 3, -52, 1, 94, 65, 11, -15, 18, 14, 46, 46, -37, -78, 13, 14, 7, 12, -66, -75, -17, 61, 40, 57, 49, -32, 7, -55, -81, -27, -28, 41, 65, 100, 28, -45, -52, -19, 0, -4, 18, -4, -7, -14, -35, 53, 5, -34, 4, 0, -78, -64, 31, -14, -32, 47, 23, 19, 93, 5, -34, -15, -74, -74, -1, -28, 15, 43, 22, -5, -22, -26, -30, 49, 75, 82, 65, 2, -66, -49, -28, 37, 9, 9, 38, -4, 24, -7, -24, -12, 4, 60, 79, 32, -1, -81, -93, -26, -21, -21, 95, 62, 0, 6, -24, 15, -29, 20, 11, -51, -55, -7, 19, 83, 48, 1, -42, 1, -28, 34, 12, 5, -2, 10, 28, -30, -58, -48, -28, -13, 3, 43, -7, 10, 4, -6, 20, -77, -14, 49, 41, 25, 27, 12, -28, -51, 91, 18, 32, -6, -13, -22, -25, -53, 35, -47, -5, 107, -1, -2, -17, 2, -28, -32, 8, -10, -30, 5, 97, -42, 3, -45, -68, 25, 11, -18, 29, -80, -10, 12, 41, 35, -1, 0, 31, 4, -12, -8, -53, -15, 86, 38, 78, 53, -24, -23, 8, -64, -37, 34, -54, -63, 12, -52, 6, 42, 66, 62, 7, 9, -74, -23, -12, -44, -3, 77, 24, 29, 59, -36, -81, -91, 27, 66, 52, 42, 12, 0, -31, 1, -40, -69, -44, -34, 3, 61, 28, 41, 63, 26, 37, -39, -32, -20, 29, -1, -4, -30, -31, -30, -31, -10, 31, -36, -5, 117, 13, 36, 18, -3, -26, -49, 6, -75, 21, 8, -34, 65, 30, -25, 40, -17, -21, -37, -19, -22, 1, -6, 6, 48, 74, -25, 1, -24, -103, 41, -14, -52, 10, -71, -26, 54, 40, 22, 21, 20, -30, -6, -34, -11, 28, 46, 73, 26, -1, -18, -23, -5, -64, 22, -23, -34, 58, 25, 47, 51, 39, 24, -69, -68, -21, 1, 8, 93, 37, -59, -38, -15, 29, 35, 61, 11, -73, -75, -27, 0, -3, 76, 1, 39, 3, -26, -14, -23, -75, 14, 0, -44, -15, -24, -1, 13, -11, 27, -34, -2, 83, 29, 28, 51, -34, -30, -26, -51, -32, -32, -8, 36, -1, 0, -1, 1, -4, -9, 61, 0, 66, 38, -17, 5, 0, -69, -31, -31, -47, -29, 69, 104, 31, 63, 42, -21, -24, -4, -28, -110, 18, -14, -31, 54, -20, -17, -1, -9, -21, 7, 9, 9, -30, 31, 1, 20, 53, 23, -15, -60, -37, -70, -17, -2, -15, 53, 20, -40, 21, -74, -56, 64, 73, 9, 21, -45, -119, -9, 46, 44, 60, 18, 2, -25, 21, -25, 30, -73, -10, -21, -49, 56, 42, -6, 63, -36, -24, 74, 23, 76, 25, -69, -49, -20, -70, 3, 52, -68, -13, 40, -10, -22, 56, 0, 59, 41, 35, -22, -62, -121, -58, 6, 70, 85, 83, -44, -46, -18, -48, -23, -31, -64, -64, -2, 52, 71, 51, 86, 3, -48, -11, -51, -48, -62, -9, -56, -40, 28, 52, 15, 40, 40, -54, 0, -2, 34, 5, -17, 39, -68, -13, 32, -12, 62, 3, 17, -39, -17, -30, -22, 30, 30, -11, 35, 21, 19, -40, 5, 15, 4, 39, -12, -24, 5, -64, 27, 106, 9, 63, 11, -21, -4, -46, 10, -34, -57, -38, -51, 17, 17, 15, 11, -31, 12, 11, -4, -17, -48, -58, -43, 21, 49, -19, 28, -12, 31, -11, 36, 42, -69, 2, 0, -56, 3, 2, 19, 31, -32, 72, 23, 0, 43, -5, -49, -3, -68, -6, -12, -14, 39, 17, 14, 68, -54, -26, -52, -52, -18, 13, 47, 10, 31, -18, 6, 15, 19, 58, 65, 24, 29, -24, -38, 24, -70, 15, 2, -65, 1, 7, -83, 23, 25, -22, 22, -39, 11, -1, 27, 55, 41, 26, -43, 23, -8, -66, 18, 36, 40, 75, 14, -54, -34, -45, -73, 53, 15, -58, 23, 20, -49, 61, 54, -30, 61, -2, -93, 11, -21, -44, 38, -22, 15, -13, 47, -21, -17, -12, -60, -20, -9, 52, 23, 41, 41, -11, -21, 31, -19, 26, 65, 0, 19, -28, -58, 3, -10, 1, 57, 2, 52, -7, 29, 22, -82, -15, 3, -48, 11, 25, -27, 1, -8, -4, 78, -35, -22, -18, -86, -48, 40, 72, 19, 11, -46, -61, -46, 20, 52, 89, 30, 49, -19, 21, -5, 18, 21, 32, -12, -18, -11, -40, 51, 0, 18, -4, -9, -21, 25, 4, -8, -54, -21, 14, 7, 95, -36, -62, 1, -44, -42, 61, 19, -6, -43, 21, -26, -59, 36, -7, 25, 18, 51, -9, -36, -29, -74, 7, 43, -24, 9, -58, -73, -47, 0, 21, 56, 95, 31, 21, 20, -60, -59, 29, -39, 26, 66, -43, 11, -28, -122, -2, 11, 71, 106, 65, 47, 1, -71, -27, 9, -29, 45, 18, 29, 22, -60, 24, 21, -29, 7, 31, -21, -30, 22, 27, -70, 23, 14, -74, -13, -22, -61, 17, -24, 14, 29, 22, 64, -2, -18, -14, -88, 5, 0, -32, 2, -19, 13, 1, 31, -3, -18, 56, -35, -39, 35, -68, -42, 83, 47, 11, 97, -2, -17, 28, -38, 13, 17, -40, 31, 7, 4, 10, -75, -19, -43, -38, 93, 68, -8, 7, -21, -56, 19, -56, -4, -52, -57, -27, 26, 1, -13, 17, -36, 36, 41, 54, 32, -4, -41, -61, -32, -10, 14, -6, 29, 39, 92, 39, 58, -12, -90, -17, -58, -62, -1, -58, -13, 32, 15, 27, 7, 22, -31, 28, 45, 4, 91, -23, -4, 19, -90, -9, 25, -69, -15, -51, 6, 26, -9, -6, -19, -24, 39, 61, 54, 43, -39, -56, 15, -22, 58, 41, 41, 30, -37, -7, 12, -42, 32, 11, 7, 9, -53, -29, -29, -72, 15, -2, -36, -15, 54, 58, 44, 45, -2, -46, -80, -72, -25, 5, 26, 52, 127, 26, 3, -23, -64, -70, -53, -5, -19, -2, 30, 64, 14, -3, -51, -79, -28, -1, -15, 44, -24, 34, 120, 58, 39, -5, -48, -70, 15, -45, 24, 43, -4, 24, -8, 15, 2, 5, 25, 27, -25, -2, -29, -34, -43, -4, 68, 23, -14, -20, -21, -36, 11, 43, 19, 11, -17, 19, 41, -51, -7, -34, -54, -46, 10, 63, 41, 53, 83, 28, 9, -37, -120, -70, -43, 47, 65, 41, 0, -53, -15, -34, -21, -11, -41, 20, 2, 18, 79, 10, 24, 54, -64, -51, -11, -40, -45, 54, 27, -1, 43, -22, 61, 4, 34, 17, 1, 38, -56, -17, -42, -105, 6, 44, 59, 66, 4, -36, -19, 5, -80, 9, -14, -58, 9, 36, 57, -2, 27, 19, 0, 25, 20, 70, 13, -25, -28, -63, -114, -18, 31, 46, 46, 95, 9, -27, 3, -32, -82, -30, 61, 28, 65, 73, -34, -62, -26, -96, -6, 44, 17, 79, 24, -26, -54, -83, -30, -55, 0, 21, 31, 62, 41, 82, 47, 17, -9, -68, -42, -21, 27, 13, 38, 4, -100, -21, -62, -22, 22, 7, 89, -15, -43, 27, -58, -26, 71, 24, 15, 9, 14, -4, 1, -1, -69, 14, 5, 39, 79, 66, -36, -68, -49, -31, -43, -29, 18, -27, -22, 49, 11, 17, 32, -25, 40, 75, 34, 55, -46, -76, -69, -75, -7, -20, 49, -6, -13, 41, -14, -3, 12, 23, -14, 48, -15, -8, -4, -43, 2, -53, -12, 22, 4, 34, 49, 23, 29, -44, 24, -1, -62, 18, -6, 2, 71, -39, 35, 39, -45, 27, 27, -31, 9, -37, -24, -71, -10, -54, 20, 95, 21, 55, 29, -55, -65, -44, -28, 20, 40, 18, -24, -35, -83, -19, -6, -26, 28, -8, -8, 63, -18, -15, 8, 3, 55, 11, 14, -36, -44, -18, -32, 13, 30, 19, 15, 47, -71, 15, 13, 8, 69, 7, -47, 28, -52, 2, 21, -53, 1, -32, -21, 2, -30, -4, -51, 8, 26, 1, 55, 26, -22, 74, -15, 41, 79, -18, 1, -91, -89, -73, -24, 12, 34, 63, 23, -9, 12, -11, -12, -29, 20, -25, 54, 41, 32, 69, 13, -28, -83, -47, -41, -53, 19, 53, -37, 18, -21, -8, 0, 62, 42, 60, 57, 10, 5, -61, -1, 35, -36, -9, -18, -18, -42, 18, -41, -31, -65, -17, -18, 6, 61, 45, 13, 64, -29, -39, 37, -39, -19, 62, -29, 13, 9, -14, -22, -48, 61, 54, 9, 27, -3, -15, -87, 23, -3, -25, 1, 28, 48, 19, 13, -51, 9, -26, -61, 39, -29, -81, 35, 55, 38, 22, -38, -27, -40, 66, 66, 42, -27, -14, -69, -65, 57, 4, -45, 44, -4, -52, 29, 10, 10, -19, 3, -41, 19, 40, 25, 26, 29, -13, -53, -3, -23, -68, 19, -3, 52, 103, 26, 28, -28, -45, -4, -13, 20, 36, 17, 45, 7, -3, -55, -82, -61, -55, 6, 43, 79, 29, -17, -29, -62, -54, 34, 37, 37, -2, 25, -27, -76, -31, -5, 13, -8, 34, 57, -21, 17, 53, 5, 37, 38, -3, -28, -54, -65, 24, -12, -8, 12, 31, 46, 13, 11, 6, -51, 0, 42, -40, -21, -18, 8, -5, -2, 30, 8, 6, 18, 58, -5, -43, 12, 0, -43, -6, 12, -36, -31, -42, -13, 14, 27, 51, 117, 9, 31, 7, -53, -106, -43, -72, -18, 0, 68, 64, -19, 6, -34, -99, -11, 20, 25, 77, 45, -3, -32, -28, -55, 8, -55, 4, 0, 0, 37, 47, 6, -7, -44, -15, -23, -68, 6, 23, 52, 94, 36, 12, -12, -60, 3, 19, -25, 18, -37, -27, -29, 9, -29, 24, 58, -32, 4, -2, -64, 38, -3, -52, -1, -56, -27, 62, 77, 18, 55, 39, -4, 14, 77, 12, -15, 12, 26, -23, 1, -7, -42, 6, -63, 9, -3, -47, -19, 9, -9, 66, -11, 22, 3, 12, -9, 1, -11, 3, -42, -35, -36, -30, -30, -27, 61, 26, 35, 21, 32, -59, 7, -24, -54, 58, 7, 13, 102, 19, -61, -59, -82, -95, 21, 14, -34, 36, -24, -10, 73, 109, -39, -24, -27, -60, 30, 2, 30, -4, -36, 31, -40, 35, 9, 41, -23, 24, 55, -5, 34, 4, -60, 6, -8, 8, 62, 60, -27, -6, 1, 9, -58, 49, 14, -69, -11, -47, -71, 37, 31, 71, 66, 49, -26, -6, -45, -57, 28, -77, -7, 20, -24, -47, 20, -34, -15, 77, -10, 10, 44, -6, 27, -41, -18, -9, -30, 1, 76, -70, -18, 36, 0, 15, 64, -24, -56, -11, 8, -9, 43, 59, 42, -47, -43, -61, -59, 15, 7, 32, 36, -9, 17, 102, 3, 5, -56, -9, -20, -49, 20, 17, -14, -34, -18, -26, -32, 70, 10, 28, 59, -6, 55, -12, -30, -26, -59, -1, -14, -38, -24, -56, 6, 32, 14, 56, 0, -17, -29, -39, -34, 1, 34, 21, 55, -2, -25, 26, -62, 11, 85, -20, 0, 5, -7, 0, 7, 21, -15, -83, -10, 21, 32, 104, 80, 60, 44, 15, -11, -71, -113, -100, -58, 3, 25, 86, 54, 5, -13, 11, 0, 0, 27, -17, -32, -32, -9, -5, 18, 10, -21, -76, -19, 10, 60, 8, 36, 47, -59, -29, 45, -31, -49, 4, -36, 76, 48, -6, -9, 19, -19, -26, 40, 10, -64, -74, -5, -80, -28, 49, 86, 82, 57, 4, -83, -2, -4, -37, 12, 12, -14, 69, 19, 19, 38, -69, -29, -7, 9, -44, -11, 22, 6, -42, 0, 42, 11, 6, 100, 12, -57, -52, -41, -57, 72, 60, 60, 36, 12, 19, 0, -37, -60, -31, -89, -19, 61, 68, 7, -2, -34, -2, 21, 59, 29, -27, -41, -1, 65, 54, 72, 41, -37, -7, 7, -4, -32, -41, -26, 5, 8, 56, -24, -48, 2, -2, 41, 54, 8, -34, -104, -19, -26, -47, 37, 65, -8, 30, 68, -24, 37, -28, 0, 0, -20, 36, -4, -15, 36, -55, -17, -18, -68, -3, 26, 36, 2, -7, -43, 0, -25, -19, 48, -30, -71, 0, 8, 22, 10, 9, 21, 24, 37, 17, 30, 11, -36, 86, 18, -41, -27, -27, -54, -21, -5, -26, -65, 42, 14, 49, 103, 19, 15, -15, -21, 43, 0, -2, -54, -72, -48, -23, -4, -31, -28, 9, 44, 0, 15, -9, -19, 29, 43, 42, 52, 37, -20, 11, 2, -62, -15, 18, -89, 3, -6, 17, -20, -14, -3, -1, -15, 27, 83, 8, 19, 39, -10, -66, 57, -9, 1, -35, -88, -22, -13, -23, 47, 18, -28, 45, 49, -40, -7, 52, 23, 45, 11, -88, -40, -55, -20, 85, 2, -70, 25, -7, 57, 41, 47, -9, -38, -18, -68, 14, -58, -12, 26, 77, 56, 60, 46, 3, -29, -35, 2, -27, -11, 22, -32, -86, 12, 3, -13, 28, 71, 32, -20, -1, -12, -25, -35, 0, -18, -98, -41, 17, 1, -17, 35, -15, 5, 70, 53, 72, 20, 40, 19, -27, -38, -28, -48, 57, 18, 83, 30, 4, 18, -57, -1, -29, -57, 34, -51, 13, 13, -62, -51, 19, 20, 45, 35, -22, 19, -69, -17, 65, -44, 14, 75, -54, -5, 62, -39, -18, 9, -20, -69, 32, 80, -4, 0, -44, -69, -52, -32, 43, -9, -4, 10, 37, 20, 3, 3, -7, -14, -10, 10, -2, 17, -46, 42, 11, -31, 34, -62, 31, 17, 32, 28, 8, -3, -6, 10, 9, 9, -110, -61, -58, -15, 70, 54, 20, 83, 8, -21, -11, -68, -82, 13, 89, 25, 54, 2, -47, 20, -65, 0, 0, 4, 65, 103, 35, -6, -65, -64, -19, -54, -26, 3, -25, 9, 56, 86, -14, -31, 10, -61, -45, 30, 7, -42, 38, -41, -44, 18, 0, 6, 48, -86, -25, -48, -39, -35, 19, 48, 64, 57, 76, -27, 7, -13, 45, 1, 26, -53, -34, -24, -1, -5, 3, -30, 19, 48, 35, 68, -5, -45, 17, -55, 43, 65, -21, -35, -41, -66, -65, 65, 32, 31, 47, -78, -6, 8, 12, 45, 37, -53, -19, -29, -48, 40, -7, 11, -36, 54, -12, 7, -3, -43, 8, 3, 24, 82, -27, -68, 29, -40, -23, 31, -40, -47, -38, -18, 70, 98, 63, 25, -40, -68, -80, 27, 34, 4, -35, -27, -56, 57, 57, 8, 44, -17, -106, 60, 72, 51, 105, 46, -21, -38, -12, -22, -71, -9, -19, -37, -6, 45, 37, 11, 42, 35, -28, -52, -1, -3, -38, 63, -4, -51, -41, -78, -64, 52, 97, 60, 106, 51, -15, 29, -4, -4, -21, -2, -12, 31, -30, -45, -8, 7, -71, -8, -7, -85, -23, 20, -12, 45, 56, -6, 0, -17, -74, -5, 91, 66, 64, 40, -58, -65, 2, -38, -26, -8, 1, 21, -12, 12, 37, -41, -12, 43, 10, -10, -26, -11, -45, -31, -17, 44, 40, -8, 8, -5, -28, -45, 77, 17, 3, 3, 8, 1, 4, 1, -10, -9, -64, 9, -7, 20, 22, -55, -1, -69, -58, 4, 47, 108, 9, -5, 32, -27, -34, 62, 13, -14, -48, -1, 13, -12, 1, 2, -9, 40, -3, 41, 42, -34, -9, -19, 24, -70, 13, 20, -8, -5, 64, -9, -4, -21, -20, -68, 28, 9, -29, 51, 25, 19, 6, -45, 1, -13, 17, 9, -38, -34, -79, -9, 63, 21, 61, 5, -22, -29, -44, 26, 12, -23, 30, -12, -6, 0, 7, -70, -6, -15, 5, 116, 36, 55, 13, -120, -83, -63, -27, 6, 18, -17, 34, 56, 54, 91, -53, -70, -65, -19, 34, 45, 82, 62, -32, -28, -32, -47, -10, 3, 10, -62, -24, -36, -40, 23, 44, 79, 70, 11, -14, 25, -15, 37, 74, -3, -53, -30, 66, -3, 26, -13, -85, -74, -56, -28, 25, 8, 24, 70, -7, 3, -15, 6, -47, 18, 45, 28, 26, 28, -12, -98, -60, -66, -57, -8, 24, 51, 94, 72, 31, 1, 3, -42, 11, 81, -42, -17, 17, -24, -31, 48, -42, -20, 8, 9, 82, 12, 29, -37, -116, -12, -53, -11, 95, 31, -4, -9, -23, -13, 39, 3, 6, -21, -102, -14, -5, 60, 57, 4, -47, -75, -77, 3, 52, 68, 54, 18, -13, -75, 20, -21, -9, 119, -3, -40, 0, -8, -9, -19, -14, 9, -32, -2, 68, -9, -30, 52, -22, 35, 88, -55, 6, 18, -38, 71, 13, -21, -42, -27, -30, -19, 52, 28, -17, 5, -52, -17, -13, 9, 42, 52, 26, 1, 43, -13, -54, -87, -1, 14, 48, 29, -14, -20, -17, -21, 45, 49, -65, 28, -40, -24, -27, -36, 51, 1, -53, -5, -47, -31, -17, -1, 58, 65, 43, 41, -3, -41, -63, -2, 26, 14, -11, 61, -34, -61, 69, 17, -14, 21, -26, -39, -7, 47, 41, 39, -34, 40, -5, -9, 47, -39, -36, 36, -64, 10, 30, -65, -4, -35, -47, -19, -28, -44, 43, 27, -3, 55, -2, -4, 42, 14, 2, -53, 5, -44, 17, 93, 4, 35, 19, -73, -78, -21, 4, 73, 57, 57, 0, -61, -40, 36, 42, 2, 8, -34, -59, -31, -73, -32, -26, 9, 70, 66, 51, 13, -53, 32, 40, 48, 19, -23, -32, -102, -63, -4, 15, 24, 57, 15, 14, -45, 14, 1, 66, 56, 19, 0, -12, -34, -53, 28, -28, -73, 10, 12, 58, 52, 71, -22, -61, -53, -91, 4, 35, 46, 28, 29, -56, -76, 9, -37, -65, 12, -52, 2, 69, 51, 111, 0, -6, -23, -57, -40, -22, -24, 0, 76, 38, 32, 35, -21, -32, 63, -42, -25, 5, -15, 66, 45, 28, -35, -61, 14, 38, -4, -17, -49, -100, -49, 8, 15, 48, 60, 15, 0, 22, 28, -1, 49, 59, -9, -1, -22, -6, -60, -17, 77, -11, -6, -19, -73, -91, 49, 22, 0, 26, -88, -15, 14, -4, 12, 46, -13, -14, 3, 48, -48, -26, 14, -43, -4, 13, -26, 83, -3, 0, 44, -81, 3, 9, -14, 49, -31, -20, 26, 6, 12, 56, 9, 13, 0, 32, 34, -30, 4, 19, -3, -57, -55, -36, -86, -20, 0, 52, 68, 22, 25, 7, -52, 21, 49, 43, 28, -70, -31, -34, -8, 71, 5, -9, 6, -51, 34, 57, 6, 15, 10, 19, -48, -12, -51, -62, -32, 29, 6, 64, 43, 3, -8, 8, -37, -46, 18, -1, 40, -21, 19, 41, -57, 34, 44, -43, 10, -40, -91, 18, 0, 23, 124, 4, -9, 0, -75, -1, -28, 30, 15, -4, 23, 48, -42, 49, 15, -25, 45, 2, -10, -5, 24, 36, 37, 13, -46, -46, -71, 1, 88, 26, 56, -23, -103, -58, -37, -27, 69, 99, 10, 35, -4, -12, -27, 23, 21, -14, 32, -9, -30, -48, -21, -55, 35, -14, 44, 26, -62, 35, -14, -47, 0, 4, -55, 22, 48, 46, 0, 3, -27, -77, 43, 54, 70, 43, 5, 1, -68, -1, -5, 27, -13, -18, -69, -54, -35, 13, 56, 32, 115, 19, 6, -17, -43, -68, -31, -10, 21, 38, 29, 36, -15, -23, -15, -18, -21, -47, -37, 10, 72, 28, -13, -53, -97, -32, 27, 26, 46, -32, 22, 20, 18, 27, 38, 2, 31, -27, 28, -29, -69, 38, 12, 1, 44, 65, -31, 43, 23, -35, 25, 23, 0, 29, -1, -46, -19, -70, -38, 66, 22, -3, 3, -38, -73, -23, -18, 17, 24, 38, 75, 64, -6, -42, -20, -55, -46, 26, 34, -11, 0, 62, -68, -77, 12, -79, -63, 1, 1, 26, 34, 37, 88, -17, 41, 12, 19, 38, 15, 18, -30, -59, -13, -95, -29, 5, 5, 58, 35, 8, -29, 8, -2, 57, 39, 44, 10, 1, -34, -64, -61, -53, -19, 44, 7, -41, -21, -51, 26, 71, 56, 96, -49, -70, 19, -8, -46, 3, 8, -5, -7, 27, 54, -3, 42, -14, -26, 3, -31, 0, 35, 14, -18, -38, -36, -51, -39, -5, 75, 29, 32, 29, -108, -5, -2, 18, 51, 13, -46, 8, 17, 9, 78, 20, -62, -18, -45, 12, 48, 46, 4, -27, -58, -69, -45, 17, -30, 32, 30, -19, 51, 6, 7, -55, -23, -45, -7, 48, 29, -26, 49, 17, 18, 54, 32, -83, -86, -1, -13, -2, 42, 31, -25, 21, 65, -28, 30, 8, -54, -38, -24, -65, 34, 12, 11, 69, -10, -35, 62, -13, 6, 9, 32, -27, 21, -27, -58, -37, -80, 38, 96, 49, 53, 11, 11, -1, 66, 58, -35, -86, -62, -87, -51, 20, -55, 6, -25, -1, 56, -29, -2, 39, 23, -21, 14, 13, 2, 31, 76, -2, 0, 30, -3, -1, 14, -12, -54, -8, 38, 0, -44, 26, 6, -54, 30, -20, -73, 18, 47, 59, 61, 0, -38, -85, -88, 6, 4, 7, 28, -5, 1, 20, 38, -24, -24, 8, 15, -4, 42, 17, -42, 22, 1, 0, 58, 8, 15, 8, -28, 29, -43, 31, 17, -47, -1, -69, -23, -10, -19, -17, 47, 15, 24, 30, 18, 17, -25, -12, 13, 3, 46, 65, 1, -39, -6, -6, -36, 34, -36, -10, 13, -22, 13, 20, -9, -5, -27, 29, -70, -80, 64, 30, 30, 48, 26, 20, -53, -14, -69, -58, -73, -41, 40, 61, 34, 61, 54, -55, 29, -38, -10, 55, -39, -65, 19, -42, -58, 46, 55, 1, 52, 73, -9, -9, -9, 1, -45, -63, 20, 4, 36, 119, 26, -40, -36, -47, -54, 24, 46, 21, 27, 1, 15, -15, 26, 23, -23, -72, -26, -83, -31, 38, 64, -9, -27, 1, -38, 11, 7, 60, -28, 13, 77, 22, 17, 4, -27, -32, 11, 69, -9, 10, -37, -40, 5, -23, 57, -18, 10, -18, 59, -9, 37, -40, -88, 13, -1, 43, 74, -22, -66, 6, 19, 49, 13, -61, -51, -87, -61, 29, 48, 73, 9, 28, 7, -11, -28, -30, -43, -40, 2, 24, 64, 58, -21, 1, -12, 22, -54, 42, 6, -23, 35, -2, -41, -3, 36, -61, 2, 62, -41, 9, 46, -65, -7, -82, 3, 9, -1, 20, 1, -32, -66, 19, 43, 91, 69, 48, 4, -24, -115, -52, -21, -22, 26, 81, 35, -37, -21, -47, -27, -7, 98, 20, 24, 38, -81, -52, 22, -13, 48, 36, 9, 64, -10, 63, 32, 26, 11, -41, -9, 10, -69, -34, -5, -78, -68, 61, 48, 69, 43, -39, -19, -14, -25, 49, 8, -76, -41, -43, -6, 8, 71, -24, 2, 11, -9, -21, 36, 2, 10, 6, 70, 7, 24, -45, -42, -58, -61, -2, 10, 46, 37, 28, 8, 51, 35, -36, -34, -27, -80, -3, 125, 24, 11, 13, 0, -82, -27, -14, -2, 29, 15, 38, 29, -30, 6, 6, -124, -42, -42, 32, 107, 68, 18, -51, -68, -27, 45, -27, 19, 56, -23, 10, 72, 29, -31, -20, 0, -62, -69, -3, -27, 32, 89, 32, 47, 1, -29, 20, 8, -41, -31, -72, -85, 36, 85, 71, 105, 19, 2, -17, -64, 4, -12, -23, 23, 54, 11, -23, -1, 5, -66, 11, 11, -5, 11, 75, -3, 29, -15, -109, -15, -2, -20, 11, 65, -13, 36, 49, 30, -1, -5, -13, -27, -14, 7, -48, 43, 30, 9, -4, -61, -32, -58, -31, 95, 0, -29, 11, -10, -6, 43, 71, -4, -68, -45, -10, 19, 39, 104, 12, 9, -21, -43, -11, 5, -66, 0, 36, 48, 24, 31, -19, -42, -42, -17, -3, -39, -56, 23, 0, -48, 73, -26, -51, 66, 25, 4, 17, -39, -35, -3, 2, 20, 25, 34, 18, -24, -30, -71, -70, 1, 60, 60, 51, 32, -29, 25, -38, -5, 7, 45, -27, 8, -6, -53, 0, -29, 22, 8, -47, -45, -13, -21, 24, 6, 36, 52, 27, 38, 41, 20, -26, -25, -8, -111, 1, -36, -39, 68, 27, -31, 10, 3, -15, -58, 18, -21, 2, -13, -7, 26, 38, 69, 40, 34, 9, -102, -8, -32, -77, -18, 54, 48, 35, 47, 9, -98, 11, 6, -51, 70, -19, -20, 62, -8, 66, -6, 0, -56, -78, 11, -22, 21, 74, -41, 28, 12, -10, -36, -39, -6, 30, 49, 45, -49, -61, -12, 46, 56, 57, -12, -49, -73, 8, 23, 80, 3, 11, -29, -86, 19, 2, -26, -22, -36, -42, 52, 120, 69, 18, -31, -35, -109, -59, -22, -53, 18, 29, -1, -1, -21, -20, 46, 45, 90, 11, 17, 4, -92, 29, 30, 35, 21, -8, -10, -52, 36, 38, 5, -39, -64, -31, 5, 25, -4, -39, -58, -44, 42, 28, 23, 45, -31, 68, -11, 37, 27, -43, -47, 52, -5, 3, 22, -48, -80, 3, -10, 37, 117, 5, 1, 6, -32, -55, 35, -17, 37, -3, 38, -47, 32, 17, -45, 5, -17, -32, -5, -32, -15, 43, 32, 3, -7, -38, -69, 6, 70, 54, 75, 48, 23, 18, -61, -34, -11, -69, 0, 51, -17, 20, -12, -51, -20, -65, -8, 63, -4, -32, 59, -5, -57, 44, 62, 25, 10, -22, -71, -95, -83, -21, 31, 62, 77, 40, -23, -41, -53, 3, -6, -11, -27, -49, -19, 52, 47, 59, -7, 7, -4, 5, 80, 15, 29, 23, -83, -36, -47, -48, -9, 21, 71, 9, 47, 53, 31, 13, -14, -75, -79, -35, 1, 18, 41, -28, 73, 12, 21, 29, -45, -89, -38, -10, 34, 5, -25, 13, 3, -13, 18, 61, 34, 8, 85, 59, -13, -41, -66, -21, -58, -1, 24, -29, 20, -43, 0, -5, -14, 52, 29, 24, -28, -27, -18, -13, -28, 66, -21, 7, 110, -45, 0, -6, -106, -4, 9, 12, -1, 32, 44, -47, 32, 65, -22, 10, 25, -26, -26, 23, 28, -10, 40, 22, 2, 66, -4, -39, -54, -78, -60, -35, -59, 2, 42, 90, 100, 58, -32, -54, -96, -87, 36, 20, -11, 58, 61, -44, -1, -49, 7, 18, 23, 86, -36, -69, 0, -4, 61, 1, 11, 0, -59, 61, 28, 40, 36, 6, 11, -11, 27, -55, -5, 52, -7, 34, -21, -82, 3, -27, -17, 24, -44, -55, 19, 14, 6, 37, -69, -20, 24, 6, 42, 3, 57, -24, -31, -4, -54, -96, 2, 54, 81, 97, 45, -8, -30, -51, 56, -10, 4, 14, -78, -51, -37, -20, -46, -34, 5, 0, -5, 27, 32, -34, 3, -10, 17, 58, 68, 4, -12, -78, -91, -47, 15, 82, 3, -6, 22, -30, 19, 26, 49, -54, -42, 19, 7, -12, 34, -25, -45, 30, 18, 30, 80, -48, -18, -31, -25, 20, -7, 2, -12, -86, -48, -2, -15, -9, 20, -13, 18, -9, 18, 36, -44, 12, 60, -36, -34, 22, -26, 22, -7, -18, -35, -13, 63, 120, 103, 7, -62, -61, -72, -5, 29, -23, 26, 22, -52, -12, 32, -12, -5, 51, 76, -3, 52, 3, -58, -59, -23, -19, 63, 41, 38, 2, -5, 32, -25, 24, -7, -94, 19, 24, 20, 32, -31, -57, -8, 32, 62, 89, -38, -43, -49, -120, -36, 24, 27, 25, 68, -45, -35, -68, 30, 8, 14, 62, -39, 47, -22, -30, 14, -41, 6, -32, -12, 0, -38, 0, 69, -5, -47, 32, 19, 61, 76, 64, -25, -43, -39, -51, 22, -4, -31, -24, -27, 14, -6, 41, 53, -19, 31, -57, -10, -13, -44, -29, -23, 29, -3, -25, 43, -37, -21, 4, 51, 9, -40, 58, 12, -15, 23, 29, 20, 17, 17, 13, -3, -20, 20, 1, 27, 17, -22, -41, -65, -104, 12, 45, 57, 99, -53, -58, -25, -23, 45, 55, 9, 14, 37, -2, -26, -44, -29, -56, -27, 122, 22, 37, 52, -14, -42, -83, -85, -62, -62, 42, 95, 54, 49, 0, -14, -60, 26, 10, 1, 19, 22, -64, -8, -18, -25, 25, -18, 10, 8, -7, 39, 51, -9, 26, 26, -1, -4, 8, 42, -44, 43, 56, -47, 0, 31, -35, -6, -36, -36, 19, -4, 48, 11, -47, 3, -25, -70, -9, -18, -19, 0, 74, 42, -18, -46, -22, -56, 0, 62, 55, 51, 83, -59, -1, 12, -58, 44, 1, 4, 7, -27, -48, -52, 19, 51, 56, 116, 26, -54, -43, -66, -44, -13, 0, 69, -13, 34, -19, -122, -38, -61, 14, 96, 54, 47, -26, -24, -52, 20, 88, 38, 51, -2, 5, 4, -51, 6, 30, -41, -23, 18, -29, -28, 27, 17, -55, -19, -26, -36, -6, 42, 42, 18, 76, 15, 63, 18, 14, -28, -29, 12, -38, 56, 32, -89, -58, 8, -14, -36, 7, -62, -91, -10, 47, 78, 7, 40, 45, 17, 59, 37, 18, -69, -112, -40, -81, -68, 31, 28, 44, 29, 66, -54, -85, -47, -77, -20, 60, 69, 42, 35, -49, 35, 21, 23, 69, 29, -38, 23, -39, 0, 19, -28, 80, -18, -39, -37, -49, -9, -42, 55, 44, -45, 43, 83, -8, 61, -19, -43, 12, -69, 5, 48, -86, 55, 29, -19, 29, -13, -23, 1, 10, -20, -13, 4, -11, 87, 39, 65, 25, -76, -63, -8, -38, 51, 110, 28, -9, -35, -36, -68, -40, 0, -23, 51, 26, -10, 56, -3, -85, -2, 13, 5, 37, 48, 15, -46, -12, 5, 32, -1, 73, 2, -40, -17, 31, -11, 0, 22, -32, -112, -39, -21, -55, -3, 22, 45, 71, -10, -10, 3, -25, 21, 80, 32, 3, 37, -38, -1, -52, -35, 34, -29, 28, 95, -59, -41, -35, -42, 30, 83, 77, 0, -62, -57, -24, 46, 17, 26, -13, -119, -17, -42, -42, -22, 21, -9, 15, 68, 41, 18, 57, -18, 10, -57, -34, 19, 37, 36, 20, 19, 30, -19, 2, -73, -27, -38, -2, 53, 15, 0, -62, -19, 8, -29, 25, 10, -42, -61, -1, 18, 30, 75, 37, -88, -44, -34, -37, -3, 82, 65, 1, 32, 6, -106, 6, 12, 71, 47, 60, -20, -75, -44, -26, -17, 4, -40, -12, -47, 0, -4, 30, 3, 81, -11, 5, 80, -56, 17, 77, -56, -15, 0, -30, 42, 11, 24, 1, -72, -32, -45, 21, 15, 20, -3, -70, -18, -19, -2, 68, 57, 12, 29, -35, -53, -43, -18, -20, 25, 2, 48, -43, -7, -11, -95, -28, 4, 46, 29, -5, 57, -6, -22, 65, -15, 24, -57, 9, 0, -59, 40, -4, 30, -3, 39, 75, 25, 32, -44, -95, -52, -19, 23, -2, 3, -44, -3, 80, 12, 6, -32, -62, 20, -17, -19, 47, -64, -61, 42, -30, -10, 1, -24, -26, -26, 37, 75, 15, 3, 36, -36, 25, 20, 18, 25, 42, 20, 54, 29, -34, -28, -25, -6, -57, 12, 34, -43, -2, -43, -45, 17, 7, 46, 22, -73, -66, -62, -22, 79, 102, 51, 42, 2, -28, -32, 26, -34, -66, 57, 0, -8, 54, -37, 6, 40, -1, 28, 59, -29, 6, 20, -8, 7, 14, -58, -27, 11, -8, 42, 14, -53, -37, -61, -29, 14, -58, 12, -12, 20, 41, 85, 43, 38, 55, 12, -18, -57, -64, -64, 10, 46, 41, 30, 46, -73, -65, -22, -59, 11, 3, 8, -13, 7, 28, 72, 27, -44, -37, -89, -21, 30, -8, 26, 70, -3, -29, -31, -64, -40, 13, -2, 72, 79, 25, 49, -6, -30, -45, 31, 31, 80, 7, 10, 28, -36, -60, -30, -28, -17, 60, -4, -25, -66, -105, -32, 11, 79, 102, 37, 55, 19, -30, -14, -71, 2, -41, -3, 39, -49, 20, 4, -11, 38, 46, -43, -4, 14, 13, 11, 24, -18, -41, -24, -2, -14, -15, 39, -43, -15, -3, -76, 0, -22, -51, 23, -21, 30, 88, 24, 48, -9, -57, 14, -7, 19, 55, -15, -32, 25, 15, 1, 76, 3, -104, -76, -90, -65, -2, 34, 71, 93, 89, 61, 52, -7, -32, -17, -28, -36, 28, -37, -35, 47, -2, -13, -13, 23, -3, -10, 13, 6, -86, -7, 8, 64, 71, 42, -13, -72, -100, -53, 35, 93, 51, 30, -15, -76, -70, -80, -28, -7, 23, 9, 37, 28, 23, 43, 35, 5, -20, -10, -4, -36, -31, -58, 36, 45, 38, 43, -53, -35, -31, 57, 64, -5, 7, 21, -79, 21, 44, -47, 17, -52, 0, 4, 14, 34, 72, -58, -13, 9, -75, -26, 14, -11, 37, 30, 85, 4, -18, -79, -13, -34, 3, 55, -23, 21, -52, 35, 34, 0, 56, -63, -68, -4, -63, 7, 105, 0, -14, -5, -2, -3, 43, 61, 26, -75, -15, -59, -110, 9, 12, 14, 49, 43, 3, -60, 26, 21, -22, 77, 45, -7, 78, 5, -26, -78, -79, -76, -37, 0, 34, -3, 45, 38, 23, 74, 0, -20, -43, 39, -24, 14, 89, -35, -53, 39, -15, -24, 72, 26, -46, -30, -57, -14, -49, -19, 87, -19, -3, 75, -51, -32, 20, 1, 1, 45, 74, -9, 12, 1, 2, -57, -6, -3, 14, 21, 29, -8, -9, 23, -58, -26, -34, -30, -10, 26, 19, -57, -57, -55, -30, -18, 10, 61, 88, 46, 10, -23, -1, -5, 39, 61, -24, -10, -80, 37, 10, -24, 43, 8, -27, 49, -23, -9, -44, -76, -9, 36, 54, 45, -12, -2, -6, -58, 58, 87, -41, 51, 68, -57, 29, 74, -17, -15, -76, -85, -69, 2, 60, 26, 52, 17, -2, -6, 22, 21, 29, 59, 24, -22, -20, -53, -21, -12, -51, 15, -52, -3, -39, -13, -38, 12, 43, 62, -2, 0, -58, -70, 19, 52, 69, 5, -11, -23, -85, 38, 55, 21, 8, 0, -65, -8, -7, -17, 3, -26, 24, 36, -15, 35, -9, -29, 36, 1, 14, 36, 6, 9, -36, 6, 22, -64, 4, 40, -43, -34, 69, 34, -28, 26, -52, 14, 23, 30, 81, -2, -22, -5, -6, 58, 44, 20, 1, -31, -29, -11, -14, -26, -29, -36, -47, 17, -15, 12, 76, 0, 47, 38, 8, 2, 11, 10, -17, -62, 5, -31, -42, 70, 12, -47, -13, -21, -48, -13, 55, -24, -38, 8, -44, 38, 77, 2, 42, 64, -74, -13, 7, -15, 46, 40, 23, -27, -1, 20, 18, 39, -23, -31, -53, 26, 62, 15, 41, 13, -70, -18, 8, -92, -30, -17, -22, 25, 89, 13, -12, -20, -30, 46, 3, 14, -13, -13, -35, 51, 4, -21, 71, -10, 43, 19, -63, -27, -48, -10, 15, 13, -83, 4, -9, 57, 48, 18, -8, -61, -12, 49, -17, 66, 28, -30, 27, -3, -38, -39, 4, -24, 28, 6, 40, 76, 31, 38, 2, -49, -90, -63, 4, -44, -31, 30, -21, 22, -8, 59, 69, -6, 49, 13, -52, -14, -26, -59, -37, -32, -18, -5, 62, 78, 17, 64, 44, -38, 17, -14, -23, -68, -2, 12, 13, 60, 15, 13, -3, 24, -43, -22, -47, -106, 46, 30, -11, 42, 8, -74, 7, -70, 51, 41, 26, 85, -35, -66, -47, -57, 25, -28, -1, 27, -18, -23, 3, 10, -12, 1, 3, -23, -38, -19, -24, 27, 20, 1, 97, 14, -11, 32, -41, -36, -46, -1, 9, -41, 7, 45, 26, 42, -3, -17, -55, -53, 39, 27, 102, 68, 40, -9, -74, -54, -1, 34, 88, 48, -5, -56, -74, -10, -62, -37, 41, 25, 13, 78, -28, -53, -32, -69, -27, -10, 22, 69, 58, 110, 17, -48, -71, -39, -57, -22, 6, 3, 31, 21, 44, 15, 2, 58, -1, 3, -11, -23, -41, 3, 56, -29, -22, 34, -28, 30, 66, -32, -40, -59, -35, -12, -8, 65, -22, 8, 18, 0, 15, 20, -12, 44, 18, 62, 38, 6, -37, -41, -52, -35, 97, 38, 41, 30, 1, -30, -65, -57, -40, -15, -15, 30, 27, 10, 37, 2, 29, -11, -65, 11, -51, 8, 34, -12, 74, -40, -56, -2, -63, -56, 72, -6, -23, 85, 21, -22, 74, 14, -12, 49, 4, -38, 11, -53, -28, -14, -68, -40, -4, 65, 76, 45, 36, -42, -128, 3, -24, -30, 26, 71, 12, 30, 85, -38, -51, -6, -56, -23, 61, -37, -10, -23, -5, -37, -35, 76, 54, 41, 74, 20, -11, -94, -15, -69, -39, 27, 57, 49, 65, 6, -71, 18, -37, -12, 48, -29, -5, 17, -17, -26, 13, -12, -65, 27, -6, 55, 13, -23, 21, -56, -34, 113, 22, -18, -39, -60, -36, 35, 25, 76, 7, -32, 38, -13, 26, -6, -12, -58, 0, -9, -36, 5, 15, -34, -14, -21, -22, -25, -46, 3, 62, 47, 4, 24, 5, -32, -23, 36, 28, -21, 19, -24, -1, -61, 14, 47, 42, 99, 68, 19, -18, -40, -23, -49, -63, -6, -82, 5, 28, 30, 104, -4, 41, 8, -26, -32, -65, 9, 4, 10, 39, -6, -39, -35, 60, 1, 8, -15, -18, -11, 31, 63, 12, -36, -28, -46, -44, 36, -36, -2, 0, -26, 30, 62, -60, -40, -41, -38, 47, 80, 77, 14, 48, -57, -42, 10, -22, 5, 38, -29, 0, -43, 57, 28, 0, 0, -37, -43, -35, 61, -18, 7, 46, -68, 35, 0, -27, 39, 55, -45, 55, 54, -11, 0, -51, -22, 13, 9, 59, 5, -29, -56, -4, -76, 41, 35, 11, 89, 22, -12, -22, -60, -8, 44, 10, -11, -53, -28, -54, -22, 61, -4, -13, -46, -12, -3, -15, 25, 79, 68, -7, 0, 5, -61, -35, 68, -43, 28, 68, -4, 34, -32, -99, -52, -17, 57, 0, 9, 4, -85, -36, 23, 18, 63, 96, 59, 63, -27, -80, -31, -15, -37, 22, 35, -21, 48, -63, -20, 18, 10, 61, 68, 34, 0, 11, 28, 0, 1, -6, -85, -22, -14, -47, 18, -74, 28, -28, -27, 91, 26, 4, 55, -37, -19, 44, 25, 5, 27, -32, -79, 1, -54, -51, 27, 11, 22, 83, 22, 31, -60, -46, -45, -1, 25, 30, 29, -66, -63, -45, -28, 10, 61, 32, 31, -53, -22, -79, -47, 1, -12, 29, 71, 17, -15, 40, 11, -41, -11, 25, 5, 28, 103, 42, -35, -29, -34, 3, -2, 23, -4, -46, 17, 47, -18, -20, 7, -49, 21, 78, -11, 13, 9, -77, -5, -19, -29, -78, -2, 25, 39, 34, 47, 0, -42, -15, -38, 63, 29, 8, -18, -29, -56, -30, 10, -14, 27, 10, 52, 10, -24, 10, -90, -56, 21, 0, -9, -2, 32, 0, 19, 17, -18, 31, -7, 26, 52, 30, -22, -48, -74, -52, -69, 8, 45, 1, 64, 29, -14, 36, 9, -3, 15, 47, -37, -54, -70, -64, 28, 82, 77, 46, -48, -45, -46, -36, 61, 51, 51, 63, 49, 0, -23, -31, -66, -28, -26, 69, 0, -9, -36, -66, 15, 52, 0, 27, 22, -27, 19, 48, -51, -92, 19, -1, -34, 24, -13, -58, 23, 63, 23, 1, -1, -28, 56, 0, 59, 45, 27, 30, -21, -85, -77, -49, 0, 68, 30, -42, -35, -92, -20, 57, 7, 11, -29, -57, -13, 68, 94, 38, 22, 7, -25, 7, 17, -64, -25, -25, 2, 40, 0, 32, -37, -46, 51, -11, -27, 51, 9, 5, 64, -20, -13, 49, -28, 22, 27, -13, -3, -54, 23, -46, -36, 58, -6, 14, 27, -69, -6, -25, 62, 40, 27, 32, -56, -41, -13, -61, 68, -40, -13, 57, 4, 68, -4, -37, -3, -45, 19, 61, 43, 6, 25, 31, 43, 3, -2, -38, -59, -22, -47, -8, 72, -19, -9, 10, -17, -4, 0, -4, 47, -32, -29, 58, -11, -57, -31, -18, -70, -12, 7, 35, 8, 12, 81, 18, 11, 59, 15, -55, -32, 29, 22, 39, 78, -24, -59, -14, -54, 1, 82, -8, 4, -1, 25, -37, -21, 2, -34, -22, 47, 1, 61, -32, -66, 41, -32, -57, 35, 0, -35, 27, 20, 12, 15, 25, 47, 71, 7, -34, -62, -9, -18, -9, 1, -9, -64, -58, 0, -4, 45, 45, 61, 45, 8, -17, -21, -5, -51, 22, -35, 14, 18, -95, 6, 10, 20, -17, 3, -40, -65, -20, 66, 98, 32, 71, 10, -29, -21, 8, 51, -53, -42, 10, -26, -31, 47, -29, -45, -28, 6, 8, 21, 28, 35, -43, 15, -20, -56, 34, -43, 5, 38, -37, 19, -3, -52, 25, 26, 20, 104, 17, 57, -11, -87, -82, -85, -81, -18, 7, -13, 30, 56, 82, 88, 56, -7, -47, -91, 0, 21, 15, 0, -29, -4, 30, 0, 13, 22, -26, 13, 40, -5, -7, -80, -35, -11, 63, 63, 81, 68, 20, -64, -60, -3, -42, -70, -10, -39, -1, 29, 32, 78, 32, -8, 15, 37, -31, -65, -37, -2, 4, 9, 18, -6, -15, -17, -22, 25, -38, -55, 10, 2, -11, 34, 79, 11, 15, 21, -42, -7, -13, -64, -27, -18, 17, 34, 47, 30, 19, -7, 4, -12, -17, -48, -6, -13, -4, -20, 11, -76, 21, 27, 20, 29, 14, -29, -34, -20, 2, 1, -22, 58, 20, 49, 6, 28, -17, 23, -15, -18, -20, -19, -26, -6, -35, 24, 25, 9, 24, 8, -79, -35, 14, 14, 65, 56, -24, -23, -18, 18, 32, -3, -17, -27, -17, 0, 9, 37, -42, -45, 76, 21, 31, 80, -54, -90, -15, -49, -20, 38, -23, 3, 7, 31, 5, -31, -48, -68, -19, 4, 54, 95, 31, 31, -32, -120, -39, -17, 30, 32, -2, 7, -1, 49, 66, 37, 8, -63, -35, 18, -15, 38, -4, -40, 23, 40, -5, 27, 4, -79, -26, -14, -73, 1, 28, 61, 70, 113, -12, -64, -45, -49, 11, 30, 79, 54, 6, 20, -15, -71, -48, -7, 0, 56, 58, 51, 20, -39, -51, 22, -14, 27, 58, 11, 13, -19, 5, 4, -47, -4, -66, -39, -40, -79, 3, -26, 14, 23, 44, 92, -19, 29, 54, -22, -3, 40, 22, 19, 47, 12, -37, -70, -75, -14, -20, 7, 55, 70, 8, 35, 15, -30, -81, -26, 1, -20, 9, -47, -36, -34, 28, 70, 56, 18, -39, -20, 8, 31, 37, 66, -24, -61, -6, 0, -45, 8, 59, -38, 26, 74, -22, -71, -47, -54, 22, 25, 41, 26, -37, -7, 57, -38, -24, 45, -10, 8, 58, -7, -17, 5, -61, -66, -14, -8, -3, 5, 57, -9, -32, 85, -39, -70, 49, -28, -15, 119, -2, -11, 58, -32, -21, -44, -69, -42, 9, 8, 34, 95, 32, 35, 43, -35, -74, -72, -62, 25, 57, 0, -24, -30, -75, -13, 25, 0, 35, 41, 5, 18, 24, -32, 3, 64, 23, 44, 61, -2, -44, -95, -65, -49, 32, 107, 72, 42, -37, -45, 1, 6, 14, 28, -27, -70, 28, -45, -62, 5, -7, 14, -25, 24, -10, -36, -3, 26, 38, -18, -18, 66, 25, 12, 4, -17, -42, -78, 35, 10, 28, -46, 17, 7, 17, 45, 41, 28, -11, -3, 20, -37, -32, -56, -18, -6, 30, -23, 37, 55, 0, 82, 20, -31, 20, -8, -52, -28, -45, -42, -56, -25, 6, -18, 1, 14, -37, -20, 0, 28, 32, 59, 0, 43, 46, 37, 27, -54, -23, -12, -53, 48, 0, -94, 0, -42, 0, 14, 41, 20, 8, 96, 9, 35, 15, 7, -69, -46, -75, -71, -4, 18, 68, 85, -6, 15, 30, -51, 23, 36, -46, -2, 18, -21, -8, -7, -39, -15, 10, 53, 21, -5, -38, 13, 20, 11, -3, -38, -24, -9, -5, 42, -3, 17, -25, 6, 39, 30, 29, 59, 63, -17, -24, 0, -38, -102, -30, -42, 11, 51, -23, -5, -23, -68, 3, 31, 43, 18, 69, 65, 11, 26, -28, -65, -64, -55, -64, 29, 80, 38, 78, 9, -112, -13, -8, -40, 61, 71, -32, 48, -11, -12, -47, -38, 36, 30, -2, 24, -24, -109, -47, -41, -55, 32, 26, 9, 58, -13, -18, -28, -34, -15, 5, 7, 31, 78, -36, -17, 40, -2, -44, -5, -11, -42, 44, 46, 41, 45, -32, -13, -80, -15, -31, -41, -6, -5, -59, -32, 6, 15, 22, 60, 15, 3, 72, 42, 70, 32, -42, -55, -37, 10, 51, 43, 34, -43, -30, -60, -14, 17, -35, 17, -13, 25, 7, -6, 2, -32, -53, -24, -7, 40, -7, -31, 10, -45, -34, -18, 81, 11, -29, 56, 21, -29, 19, 38, -51, 30, 6, 105, -12, 22, 29, -40, -10, -21, -26, -28, 7, -18, 41, 15, -53, 23, -25, -12, 23, 24, 48, 17, 3, -32, 17, -21, -21, -20, 2, 34, 30, 83, -26, -76, -44, -88, -22, 53, 36, 14, 55, 7, -26, 6, 2, -21, -8, 22, 15, 0, -21, 32, -13, -17, 72, -20, -19, 23, 9, 13, 52, 10, -56, -10, -10, -32, 47, 32, 65, 19, 34, -31, -71, -32, -13, 44, 22, -2, -49, -32, -39, 18, 37, 53, -30, -36, -54, -30, -35, 3, 87, 31, 53, 24, -39, -27, -94, -19, -11, -11, 39, 74, 3, 19, -9, -12, -42, -30, 5, -52, 56, 61, 38, 19, -17, -92, -69, -6, 35, 68, 20, 4, 20, -96, -57, 55, 36, 20, 77, 14, -70, 41, 5, 13, 32, -4, -55, -70, 38, -1, 36, 61, 73, -24, 17, 14, -40, -34, -32, -93, -60, -6, 7, 29, 27, -19, -29, 18, 19, -14, 17, -19, -41, 6, -11, 5, 30, 88, 23, 36, 5, -14, 12, 0, 8, -28, 4, 3, -10, -3, -54, -41, 24, 19, 31, -10, 27, 24, -10, 30, -51, -48, 8, 8, 60, 13, -7, -35, -14, 69, 20, 29, 38, 4, -17, -22, 3, -4, -43, 14, 28, -29, 53, -19, -25, -47, -59, -6, 32, 77, 63, 34, -53, -64, -82, -39, 18, -3, 29, 13, 42, 24, -8, -11, -17, -32, -35, 23, 19, 20, 10, 21, -41, 14, 48, 13, 24, -46, -61, -29, 25, -8, 34, 11, -10, 17, 27, -6, 5, -3, -54, -39, -17, 29, 32, 88, 44, -15, -24, -68, -6, 2, -24, 30, -37, -41, 31, 30, -23, 6, -31, -40, 21, 83, 11, -41, -10, 3, 39, 37, 26, 19, 0, 25, 34, -22, -40, -40, -65, 22, -24, -43, -25, 41, 32, 14, 14, 7, -104, -35, 13, 34, 61, -4, 12, -15, -54, 47, 7, 6, 44, -23, 57, 1, -11, 5, -72, -15, -11, -37, 18, -9, 60, -45, 3, 55, -13, 32, 27, -2, 22, -15, 60, -32, 5, 24, -38, 29, 18, -94, -46, -81, -11, 7, -3, 81, -32, -46, 1, -35, -23, -7, 19, 17, 4, 41, 62, -4, 0, 14, -10, -13, 7, 2, -37, -25, 28, -8, 72, 14, -68, -29, -63, -39, 79, 63, 55, 8, 36, 4, -36, -15, -37, -103, -54, 36, 45, 68, 106, -7, -6, 3, -59, -11, -63, -48, -51, 9, 63, 56, 44, 23, -39, -21, -71, -23, -29, -52, -2, 22, 51, 89, 53, 34, 0, 27, -11, 45, 12, -22, -55, -31, -79, -15, 35, 61, -5, -27, -82, -103, -32, 22, 38, 49, 31, 30, -8, 14, 19, -10, -25, 24, 35, 20, 4, -29, -52, -78, -72, 10, 0, 41, 81, 6, 75, 64, -12, 45, 26, -37, -5, -9, -61, -8, 44, 18, 20, 6, 0, -38, -3, 51, -59, -36, 12, -51, -42, -21, -37, -7, 39, 35, 45, -57, -14, 12, 24, 35, 71, 28, -4, 17, -59, -80, 0, -45, -56, 59, -28, -32, 70, 14, -1, 55, 36, -37, 23, -26, -53, -94, -3, -29, 9, 65, 20, 43, -27, -75, 43, 25, 17, 59, -2, -18, 6, 32, 46, -14, -81, -10, 14, 46, 94, 14, -89, -103, -95, -29, 30, 56, 41, -10, 0, -35, -9, 34, 46, 7, 42, -18, -103, -4, -36, -42, 14, 15, 23, 37, 49, 75, -4, 34, -8, -28, -92, -32, -13, 10, 37, -7, -14, -35, 11, -20, -36, 10, -19, 44, 127, 79, 38, 9, -30, -48, 24, -42, -15, -1, 52, -19, 32, 14, -85, -70, -9, 3, 31, 65, 34, 54, 11, -12, 0, -44, -20, -46, -30, 6, -24, -38, 38, -55, -14, 42, -23, 27, 87, 0, -12, -21, -20, -57, -20, 17, -18, 40, 64, -26, 7, -11, -86, -59, 1, 17, 72, 88, 77, -23, -18, 12, 7, 39, 37, 39, -12, 14, 27, -5, -97, -74, -45, -51, 11, 36, 41, 5, -51, 35, 2, -39, 44, -9, -9, 53, -41, 49, 34, -19, 40, -27, -32, -18, -103, 19, -31, -6, 85, -34, -7, -3, -39, -18, 86, 27, 51, 1, 9, 32, -83, -24, -25, -40, 27, -11, 26, 9, 1, 56, 3, 19, -19, -24, 30, 4, -43, -24, -107, -49, -2, 64, 35, 5, 0, -29, 18, 7, 72, 55, -61, 19, -12, -98, 20, -55, -34, 8, 0, 13, 59, 0, 32, 13, -2, -25, -47, -21, -32, 19, 94, 32, 40, 34, -65, -31, -3, -46, -13, 24, -56, 49, -8, -26, 96, 17, 15, 49, -10, 2, -52, -37, 5, -91, -29, 57, -4, 19, 103, 40, 19, 58, -27, -100, -46, -44, 6, -8, 4, -6, -26, -25, -8, 9, -44, 65, 85, 7, 6, -19, -56, -27, 31, -72, -22, 5, 4, 52, 127, 0, 24, -13, -70, -35, -2, -15, 22, -7, -2, 6, 5, 71, -21, 17, 35, -69, 21, 4, -46, 13, -12, 9, -26, -73, -14, -58, -8, 95, 76, 76, 49, 11, -8, -10, -28, -86, -63, -100, -15, 69, 66, 58, 18, 23, -17, -14, 26, -13, 26, -54, -45, -17, -51, 28, 58, 49, -14, 10, -48, -92, -10, -32, 35, 66, 10, 12, 1, -23, 40, 19, 6, -74, 24, 35, 23, 93, 51, -40, -39, -71, -49, -53, -6, -17, -30, 52, 17, 0, 106, 27, 9, 29, -56, -40, -22, -6, 31, 34, -69, 26, 2, -46, 27, 30, 7, 18, 81, -30, -8, 42, -19, 45, 65, -47, -21, 25, -38, 21, 3, -6, -11, -35, -64, 23, -26, -25, -18, -22, -36, 3, -21, 0, -39, -43, 2, 55, 60, 30, 85, 31, -34, -11, 7, -3, -7, 59, -10, -70, -14, -52, -55, 37, 35, 51, 90, -13, 3, 32, -30, 56, 6, -30, -65, -2, 7, 48, 17, -40, -61, -25, 4, 49, 55, -56, -62, -6, 5, -6, 28, -58, -76, -55, -43, 18, 57, 49, 52, 85, 44, -9, 37, 6, -28, 40, 23, 26, 43, -41, -49, -14, -86, 19, 52, -32, 22, 0, -91, -3, -10, 48, 68, 26, 10, -60, -105, 26, 36, 0, 31, 39, -62, -35, 30, -28, -8, 18, -41, 4, -27, -13, -17, 24, 30, 17, 12, -14, -59, 20, -12, -29, 48, -19, -12, 39, 53, 13, -4, -24, 10, -26, 8, 47, 23, 42, 17, 39, -39, -30, -12, -41, -8, 29, -20, -25, 26, -35, 10, 32, -70, 4, 11, 34, -7, -2, -39, -28, 26, -4, 45, 27, -41, 18, 0, -34, 18, 48, 62, 91, 46, -5, -74, -97, -41, -40, 2, 111, 41, 21, 26, 8, -62, -26, -43, -112, -48, -13, 26, 51, 105, 76, 22, -23, -56, -85, -51, 11, 87, 3, 65, 23, -32, 45, -57, 2, 23, -63, -42, -19, -13, 35, 8, 38, -7, -7, 72, 18, 17, 1, -76, -83, 41, -36, -47, 45, -57, -36, 23, -11, 73, 62, 0, 48, 28, -35, 40, 18, -3, 30, 12, -17, -6, -75, -68, -10, 12, 41, 76, 49, 5, 20, -21, -18, -36, 8, 25, -34, -19, -13, -35, -32, 55, 103, 3, 20, -64, -60, -38, 32, 56, -11, -32, -38, -59, -45, 61, 6, -28, 59, 51, -76, -6, 35, -23, -46, 20, -1, -8, 9, 17, 11, -82, -36, 0, 37, 49, 12, -31, 14, -48, -5, 88, -29, -10, -40, -8, -20, 57, 73, 51, 2, -13, 11, -69, -27, 2, -5, 53, -29, -10, -15, -65, 52, 86, 41, 5, -18, -86, -72, -26, -26, 31, 3, 21, 13, -58, 41, 0, -30, 81, 53, 1, 40, 4, -10, 12, -24, 32, 55, -44, 39, 0, -65, -28, -62, 36, -18, -62, 31, 0, 23, 92, 24, -10, 8, -45, 38, -3, -28, 2, 47, -14, -1, -14, -59, -63, 31, -1, -14, 1, 29, 18, 25, 26, -1, -51, 40, 23, -27, 0, 51, -5, 31, 41, -40, -40, -6, -53, 6, 32, -59, -18, 15, -6, -6, 64, -7, 75, 25, 23, 18, -49, -61, -29, 2, 72, -12, -11, -8, -107, -52, -8, -15, 15, 63, 79, 61, 59, -26, -17, 11, -56, -10, -6, -82, -9, -45, 3, -27, -24, -2, 46, 18, 24, 63, -40, 72, 29, -26, -59, -17, -38, -7, 58, 72, -7, -34, -28, -61, -36, -4, 74, 51, 17, 10, -1, -23, 4, -35, 31, 30, -40, 39, 13, -19, 24, 3, -13, -55, -47, -65, 21, 30, 23, -18, 9, -23, -25, 77, 86, -25, 53, 77, -15, 45, 20, -52, -117, -71, -36, 6, 40, 41, 41, -96, -34, -27, -54, 36, 82, 44, 15, 19, -6, -76, 19, -9, 29, 26, 13, -35, -13, 15, -6, 27, 31, -83, -35, -45, 28, 94, 5, 23, 7, -90, -57, -5, 18, 18, -5, 14, 6, -15, -9, 114, 31, 17, -9, -52, -12, -38, 14, -4, -29, -82, 0, 17, 2, 22, 2, 17, 26, 32, 0, 27, -56, -21, 60, -4, -31, 5, 11, 2, 0, 19, 8, 8, -6, 17, -12, -77, -19, 56, 17, 38, 46, 31, -51, -32, 6, -43, -40, 27, -26, -24, 27, 37, 11, 42, 45, -14, 13, 40, -54, -32, 40, -51, -63, 22, -6, 1, 22, -22, -38, -21, -11, 26, 55, 55, -3, 44, -17, -64, -60, -57, -56, 11, 13, 58, 57, -5, -19, -37, 22, 26, 42, 27, -46, -35, -77, -47, 2, 54, 77, 29, 43, 34, -66, -7, -41, -9, -29, -54, 85, -14, -38, 42, -46, 24, 69, 13, 6, -34, -49, -39, -32, 4, -31, 5, -6, -24, 35, 22, -24, 58, 68, -21, 37, 54, -71, -56, -28, -32, 44, 37, 46, -7, -9, -71, -15, -20, 24, 6, 29, 78, -10, 18, 42, -83, -26, -21, -25, 56, 85, 31, 13, -48, -36, -78, -66, 22, 2, -19, 53, 1, -14, -7, 26, -42, 55, 7, 38, 6, -2, -51, 10, 57, -15, 37, 26, -59, -42, -43, 8, -1, 7, 121, 7, -39, 9, 12, -1, 37, -8, -39, -5, 32, 26, 56, -28, -77, -7, 0, 47, 0, -11, -10, -72, 7, 24, -21, 60, -14, -24, 34, -34, -29, 28, 26, 7, 82, 7, -4, 2, -21, -32, -46, 11, -57, 25, 86, -48, -6, 30, -35, 22, 36, 0, -25, -28, 65, 3, 72, 10, 1, -11, -65, -29, -63, -1, -26, -24, -17, -15, -23, 8, 68, 14, 27, -70, 2, -13, -6, 62, 48, 42, 63, 30, 26, -1, -76, -112, -18, 7, 27, 65, 63, -64, -93, 0, -14, -6, 80, 65, -15, 41, 22, -73, -34, -20, -15, 74, 35, 27, -48, -55, -77, -7, 63, -11, 19, 0, -11, 59, -17, 60, 57, -54, 37, 15, -65, 15, -27, -32, 25, -65, 26, -13, 15, -7, 47, 12, 4, 58, 7, -5, 14, -69, 17, -18, -48, 29, -41, -53, -1, 0, -21, 30, -49, 27, -24, 5, 65, -3, -34, 55, -15, -6, 76, -41, 7, -2, 74, 26, 68, 14, -82, -36, -36, -85, 2, 28, -34, 0, 38, 35, 20, 49, -8, -106, -57, -11, 5, -13, 65, -11, -40, 72, 11, 31, 2, 0, 18, -27, 66, -12, 1, -39, -102, -3, -25, 9, 121, -17, 18, 27, -51, 43, 6, -9, 3, -12, -39, 58, -24, -6, 60, -23, -1, 36, -20, -27, 36, -9, -4, 29, 45, -45, -18, 1, -13, -46, 25, 46, 25, 13, 22, -17, -98, -1, 53, 18, 66, 13, -19, -30, -29, -30, -11, -34, 82, 11, 45, 34, -31, -42, -27, -74, -27, -21, 0, 47, 38, 39, -6, -5, -42, 20, 14, 41, 100, -34, -29, -18, -71, 10, -4, -24, -12, -42, -40, 25, -42, 6, -41, -27, 48, 26, 45, 103, -25, -2, -36, -29, -21, 29, 34, 38, 46, 19, -12, -56, 45, 25, 9, -8, -76, -57, -68, -11, 93, 34, 7, 23, -24, -103, -7, -11, 12, 21, 74, -35, 30, 18, -7, -73, 0, -1, 13, 74, 24, -48, 11, -55, -34, 10, -1, 17, -10, 54, 27, -44, -5, 17, -8, -5, -42, 6, -17, 14, 111, 17, 26, 24, -87, -95, -35, -69, -6, 43, 29, -39, -29, -32, 31, 85, 94, 15, -20, 10, -36, 27, 20, -4, -64, 9, 24, 48, 65, 46, -27, -37, -7, -24, 37, 0, -24, -20, -34, 20, 26, 23, 21, 10, -46, -26, 37, -8, -12, 32, 31, -29, 4, -11, 3, -48, -29, 30, -42, -45, 20, -26, 60, 63, 64, -3, -73, -48, -81, -28, 13, 53, 2, 27, 23, -13, 6, -45, 12, 23, -15, 39, -21, -52, 35, -10, 32, 74, -8, 38, -48, 5, -5, -17, 43, -13, -74, 10, -9, 2, 85, 86, -23, -54, -49, -47, -45, 1, 44, -25, -2, 48, -3, 11, 11, 11, -31, 44, 59, 3, 29, 10, -40, -63, -12, -8, -26, 23, -22, -6, -6, -57, 47, -4, 73, 82, 8, -37, -45, -39, -12, 18, 9, -41, -52, -1, 38, -20, 39, 32, -60, 31, 17, -17, -31, 7, 24, 26, 52, 53, -11, -25, -14, -10, 65, -26, -1, -47, -99, -13, 38, 27, 10, 2, -6, 48, 29, 78, 32, -15, -24, 22, -42, -18, -55, -57, 32, -34, -31, 57, 10, 39, 12, 29, 21, -70, 19, 60, -77, -13, -24, -29, -38, 14, -40, 7, 4, 77, 92, 0, -34, -6, -8, -21, 18, -4, -69, -11, 3, 92, 7, 49, 72, -24, -18, -14, -7, -79, -29, 36, -22, -54, 40, -14, -42, 72, 11, -24, 30, -18, 55, 25, 38, -31, -31, -69, 4, -4, -35, 4, -25, -14, 52, -41, 18, 22, -35, 12, -7, 18, -27, -1, 34, -78, 1, -4, 20, 31, 76, 28, -14, 24, -53, -8, 23, -56, 8, 57, 13, 64, 93, -43, -88, -85, -115, -15, 71, 47, 85, 49, -45, -22, 62, -9, -15, -20, -13, -60, -39, 26, -76, -36, -24, -3, 51, 65, 47, 0, 41, -41, -26, 58, 6, -34, 43, 34, -17, 36, 30, -68, -56, -43, -55, 30, 37, 40, 78, -54, -14, -45, -39, 39, -11, 47, 26, 31, 27, 18, -15, -81, -6, -58, -28, -7, 3, -47, 23, 55, 17, 89, 17, 19, 30, -48, 18, -5, 7, -47, -39, 17, -43, 38, 88, -12, -13, 8, -37, -25, 13, -9, 60, 30, 43, 35, 13, -56, -52, -32, -90, 9, 45, 65, 57, 39, -34, -29, -80, 43, 13, -31, 22, 7, -37, 18, 23, 6, -47, 25, -40, 10, 0, -20, 18, -61, 63, 24, -8, 62, -23, -123, -29, -41, 25, 37, 43, 21, -60, 44, -17, -57, 29, 11, 18, 22, 32, -31, -72, 26, 0, 37, -22, 13, 25, 2, 20, 35, 20, 39, -10, -26, -38, -45, -18, -9, 63, -30, -49, 55, -54, -66, 7, -1, 32, 72, 93, 35, -52, -38, -25, -95, 31, 5, -56, 71, 31, -4, 17, 20, -56, -92, 1, -46, -34, 69, 31, 58, 60, 25, -15, -42, -17, -6, -23, 22, 61, -45, 13, 7, -66, 68, 24, 0, 34, -15, -51, -15, 30, -5, -35, 9, 54, 28, 40, 31, -41, -94, -24, -9, 8, 3, 57, -6, 60, -19, -20, -2, -61, 27, 53, -51, -15, 11, -6, -30, 7, 7, -13, 38, 91, 42, -14, 1, -41, -39, -71, 20, 12, 48, 86, 15, -53, -55, -72, -23, 66, 29, 41, 42, -31, -31, -9, -45, 7, -34, 20, 31, 3, 51, 7, -28, -28, 2, -27, 91, 17, 25, 35, -51, -82, 14, 22, -13, -1, -14, -13, -4, 45, 10, -32, -57, -21, -27, -15, 1, 1, -11, -35, 27, -49, -26, 25, -28, -5, -4, 34, 46, -5, 51, -22, -60, -3, 27, 23, 55, 52, -29, -1, 7, -22, 24, 11, -44, -29, -21, -1, 92, 37, 43, 15, -40, -24, -25, -20, -71, -74, -55, 21, 70, 38, 68, 18, 35, -57, -10, -23, -92, 36, 22, 24, 83, -36, 1, 38, -58, -52, -12, -51, 19, 39, 34, 70, -65, -63, -5, 14, 39, 21, 39, 38, -1, -10, -14, -4, -17, 34, 32, -22, -34, -55, 34, 42, 30, 23, -63, -23, -40, 28, -5, 6, -44, 18, 3, 46, 32, 3, 23, -18, 20, 43, 21, -22, 1, 10, -40, 26, 30, -13, -29, -91, -26, -62, -30, 109, 61, 24, 40, -61, -69, -57, -2, 47, 47, 8, -8, -5, -59, 32, -24, 43, 7, 57, 14, 25, -17, 1, -98, 10, 11, -39, 62, -11, -74, 0, -21, 42, 43, 29, 40, 7, -55, -21, 9, -19, 1, 44, 6, 38, -17, 57, 46, -25, 22, 47, -6, -5, 19, 14, -31, 9, -41, -90, -81, -5, 2, 61, 127, 36, 28, 1, -20, -96, -35, 52, 6, 0, -4, -17, -11, 13, 56, -3, -56, -44, -90, 26, 49, 36, 54, 20, 22, -60, 3, 15, -42, 14, 85, -20, -7, 25, 10, -55, 40, -7, -128, -6, -12, 25, 86, 40, 10, 28, -4, 25, -17, -49, -48, -85, 42, 75, 8, 6, -28, -26, 1, 48, 35, -63, -20, -18, 13, 52, 74, -54, -20, 27, -8, 2, 37, 8, -100, -9, -30, 13, 52, 19, 19, -13, -12, 40, 76, 25, -36, -70, -20, 29, 60, 95, -28, -99, -17, -25, 6, 78, 14, 22, 14, -39, -32, -5, -62, -8, 39, 42, 22, -20, -45, -15, -59, -3, 70, -40, 58, -27, -22, 52, -56, -8, -43, 27, 19, 49, 81, 19, 55, -3, -29, -17, 2, -66, 31, 1, -76, 1, -47, -1, 4, 109, 45, 65, 72, -2, -20, -47, -100, 2, 0, -45, 57, 34, 5, -23, 26, -26, -117, 9, -29, -46, -12, -25, 7, 20, 17, 100, 32, 0, 75, -21, -63, 6, -73, -55, 25, -1, 85, 78, 43, 37, -27, -107, -28, -54, -53, 71, 7, 28, -10, -57, -28, -54, 32, 70, 59, 15, -9, -29, -41, -5, 45, 53, 55, -19, -44, 6, -64, -34, 52, -73, -1, 29, 25, 110, 15, -36, -45, -45, -22, 2, 96, -18, -36, 34, -70, -5, 36, -31, 0, 21, -6, -15, 47, -21, -21, 23, 48, -63, 0, 34, -62, -59, 22, -19, 27, 83, 53, 0, -59, -17, -49, 42, 107, 29, 64, 20, -82, -46, -46, -76, -1, 40, 57, -13, 0, -3, -59, 15, -4, 10, 71, 11, 61, 77, -4, -81, -45, -20, -34, 14, 19, 58, -15, 14, -5, 27, -59, -7, 1, -43, -13, -37, -23, 44, 41, 24, 35, -65, -35, -46, 3, 19, 57, 49, -30, 27, -11, -98, -6, -48, 7, 95, 57, 19, -8, 9, -10, 15, 42, 1, 20, -77, -12, -13, -54, 38, -31, -3, 41, 2, 52, 76, 14, -26, -89, -5, -64, -77, 31, 23, 25, 74, 94, -56, -3, 29, -52, 0, 0, -66, -12, -25, -25, 24, -8, -61, 13, -29, 4, 70, 82, 72, 31, -42, -48, -78, -7, 17, 63, 52, 28, 11, -36, -71, 3, 12, -29, 19, -8, -20, 51, 7, 14, -27, -34, 46, 31, 8, 37, 54, -24, -2, -30, -23, -46, 22, 81, 21, -19, -34, -40, -37, -48, 28, 34, 32, 40, 65, -48, -76, -37, -23, 18, 72, 74, 18, -4, -49, 0, 44, -4, 13, -39, 12, -15, -29, 46, -3, -63, 22, -30, -44, -39, 14, 65, -5, 40, 44, -60, -6, -24, -69, -39, -21, 1, 12, 100, 52, 47, 44, -10, 0, -25, 5, -2, -15, -43, -27, -60, 35, 24, 54, 103, -24, -61, -68, -31, 6, -8, 40, -29, -21, 30, 48, 49, 42, 3, -19, -7, 13, -26, -22, 30, -51, -65, -31, -9, 26, 65, 37, -13, -34, -70, -86, 29, 18, 14, 63, 57, -23, 37, 30, 9, 56, 29, -11, -7, -26, -54, -35, 8, -4, 20, 56, -78, -74, -40, -70, 18, 63, -13, 29, 26, 8, 71, 113, 24, 47, 22, -52, -70, -24, 8, -41, 11, -37, 6, 2, 37, 57, 5, -68, -42, -48, -64, 13, 28, 95, 79, 32, -25, -11, -1, -73, -32, -59, -98, -27, 12, 18, 46, 89, 35, 39, 10, -70, -76, 5, 81, 61, 91, 3, -80, -57, -107, -30, 45, 17, 45, 109, -17, 0, -15, -5, -5, -20, -29, 6, -4, 14, 73, -3, -17, -83, 11, 32, -1, 14, 3, -13, -4, 11, -9, -41, -25, 6, 85, 10, 20, 13, 7, 13, 44, 38, -30, -12, -89, -42, -10, -25, -35, 7, -17, -22, 18, 106, 20, 52, 51, 5, -24, -7, -41, 27, 30, -13, 30, -30, -128, 10, 12, -11, 20, 44, -23, -29, 4, -41, -40, -41, 34, 52, 34, 37, 43, -31, -13, 47, -44, 48, 26, 30, 26, 1, -3, -105, -65, -8, -39, -38, 39, -80, -25, 10, 4, 71, 83, -3, -15, -2, -22, -18, 71, 78, 4, 47, 38, -41, -6, 25, -38, 4, 18, -19, 26, -24, -34, -13, -1, -17, 54, 3, 0, -36, -43, -47, -3, 21, 22, 54, 26, -69, -12, -44, -5, -4, -35, 64, -4, 26, 112, -57, -19, 30, -55, -51, -12, -56, -34, -7, 39, 31, -1, 81, 21, 47, 45, 19, 13, 9, -74, -38, -32, -48, 63, 42, 4, -41, -34, -24, -26, 44, 46, -25, 14, -43, 5, 72, -18, 34, 20, -17, 59, 41, 27, -36, -90, -64, -60, -44, -2, 40, -12, 0, 44, 1, 39, 47, 40, -28, -3, -47, -48, -51, -3, 27, 28, 32, 37, 2, -68, -27, 32, -6, 58, 113, 0, -41, -76, -106, -87, -43, 21, 80, 70, 1, 7, -44, -39, 63, 49, 78, 21, -5, 14, -86, -5, -15, -53, 74, -15, 59, 1, -78, -27, -31, -51, 15, 39, 23, 3, 37, -52, -46, 23, 25, -13, 39, -9, -80, 24, 13, 44, 56, -20, 43, -42, -75, 42, -37, -30, 87, -46, -10, -21, -35, 36, 74, -17, 6, 45, -39, -22, 72, 37, -25, 6, -7, 13, -21, -4, 23, 3, -49, -57, 11, -60, -62, 53, 40, 18, 37, 52, -49, 26, 29, -82, -38, -43, -54, 31, 60, 17, -9, 17, -6, -59, 24, -6, 38, 48, 19, -36, 0, -61, -10, 81, -75, -24, 8, -8, -1, -4, -20, -89, -21, 28, 57, 66, 0, 18, 7, -21, 10, 32, -94, -29, -26, 19, 19, 13, -9, -10, -28, -64, 26, -11, 38, 66, 37, -10, -2, -32, 64, -14, -18, 40, -34, -55, -9, -59, -57, 28, 56, 37, 53, 56, -34, -46, -37, -38, 18, 80, 59, 24, -26, -75, -5, 28, -66, 19, -30, -81, 42, 72, 42, 82, 45, -35, -35, -20, -30, -42, 22, -23, -46, 75, -5, -3, 26, -1, -32, -15, 63, -4, -12, 44, -11, -56, 4, -51, 30, 3, 0, 66, -36, -4, -24, -40, -38, 45, 0, -30, 15, -35, -26, 13, -3, -52, -24, -27, 13, 47, 73, 15, -51, -6, -20, -3, -22, 25, -55, -39, -1, -3, 3, 17, 22, 31, -6, 80, 5, 41, -9, -26, -26, -77, -12, 37, 47, -17, 72, 8, -47, 44, -23, 18, -34, 20, 14, 57, 11, 27, -2, -51, -34, -62, 40, 3, 38, 87, -36, -24, -13, -38, -9, -18, 28, -44, -89, 10, -42, -21, 64, 126, 22, 62, 56, 11, -6, -23, -53, -82, -45, 8, 34, -11, 61, 18, -63, 60, 25, -54, 30, -15, -24, 9, -19, -71, -37, -90, 19, 83, 37, 87, 78, -53, 20, 18, -79, -31, -47, -46, 0, 30, 56, 12, 15, -27, 4, -89, -11, -6, -43, -51, 37, 41, 56, 76, 86, -45, -85, 4, -9, 4, 45, -23, -78, -58, 20, 62, 32, 7, -8, -51, -43, -11, 18, -35, 18, 62, 1, 11, 41, 12, -30, -11, -2, 0, 29, 62, 57, 51, -9, -34, -43, 1, -8, 65, 57, -13, -44, -10, -41, -3, 24, -79, -30, -36, -29, 0, 79, 44, 45, 58, -9, -46, -10, 0, 25, 15, 13, -61, -10, -37, -36, 37, 47, 2, 28, 34, -69, -20, 53, 8, 20, 31, 14, -104, -23, -22, -52, -53, 62, 3, 6, 64, -49, -11, -57, 25, 27, 12, 24, 35, -71, 1, 23, 22, -13, -4, 41, -28, -3, 58, -82, -30, -45, -10, 38, -17, 53, -22, 15, 0, -49, -38, -35, 15, 78, 3, -24, -25, -78, 25, 121, 26, 53, -18, -22, 27, -8, -26, 1, -44, -5, 72, -7, 0, -41, -14, 5, -15, 46, 28, -15, 77, 44, 8, 41, 8, -68, -47, -37, -41, -27, 17, 37, -32, -54, 61, 8, 25, 97, 21, 14, -18, -93, -75, -87, -40, 17, 41, 68, -48, 51, 22, -29, 13, 30, 6, 29, 27, 11, 55, -57, -23, -39, -77, -28, 35, 69, 65, -10, 22, -18, -60, 20, 20, -46, 5, -3, -30, 14, -5, 82, -39, -69, 3, -40, -4, 53, 6, -2, 3, 13, 0, -30, 22, -7, 38, 35, -41, -28, -19, -37, 23, 68, 34, 36, 22, -10, -17, -42, 85, -11, -15, 7, -47, -108, -14, -25, 0, 30, 74, 88, -27, 14, 5, -75, 53, 27, -1, -39, -32, -66, -69, 77, 60, 5, 73, 47, -14, 46, 27, -90, -46, 0, -53, -2, 48, -12, 63, -34, -30, -40, -106, -39, 38, 23, 13, 36, -46, 21, 15, 43, 88, -8, -46, -5, -20, -17, 96, 65, -62, -63, -10, -51, 8, 96, 10, -11, -19, -12, 21, -14, 6, -15, -36, -45, 68, 57, 71, 87, 15, -93, -107, -64, -21, 47, 25, 64, 26, -9, 20, 35, -25, -36, -40, -24, -54, 31, -12, -32, 52, 20, 60, 39, 40, 0, -53, -13, 1, 15, -21, 52, -41, -116, -41, -86, 3, 58, 32, 72, 0, 41, -4, -10, -30, -5, -25, -24, 31, 22, 28, -2, 48, -18, -74, 20, 39, -35, 10, 11, -70, -17, -19, -31, -13, 17, 53, 36, 74, 20, 57, -41, -29, 14, -27, -58, 4, 54, -11, 20, 28, -60, -23, -48, -6, 39, -29, -6, -22, -28, 15, 23, 22, 1, -54, -11, -5, 17, 0, 61, 0, -53, 36, -26, -23, 15, 24, -59, -38, -9, -17, 24, 116, 68, -14, 4, -20, -92, 0, 13, -77, 23, 12, 9, 80, 7, -8, -7, -17, -41, 88, -6, -14, 25, -44, -17, 21, -4, 21, -43, -25, -43, -38, 32, 73, 0, 36, 92, -34, 5, 30, -61, -73, 19, 48, -23, 52, 57, -44, -3, -52, -27, -26, -42, -13, 65, 17, 2, 55, 23, -13, 57, -3, 11, 20, -116, -57, -53, -77, 25, 12, 4, 69, 0, -51, 11, -52, -64, 56, 55, 43, 91, -34, 10, -34, -60, 12, -27, 22, 82, 60, 8, 17, 30, -41, -11, 28, -40, -69, -9, -19, 20, -29, 63, 45, -41, 8, -15, -25, -23, -15, 64, -12, -27, -40, -6, -17, 10, 45, 37, 19, -44, -43, 26, -14, -27, 3, 23, -21, 35, 28, 12, 2, -23, 0, 8, 18, -40, 39, -28, -7, 19, -45, 38, -11, -66, 38, -11, -8, -37, 62, 41, 21, 42, -12, -38, -66, 11, 25, 4, -24, 79, 19, -11, 15, 9, -74, -41, -1, -13, -26, 48, 80, 66, 24, 1, -32, -25, -35, -18, -32, -56, -8, 44, 27, 56, -6, 0, -64, -44, 48, -17, -49, 60, 19, -2, 77, 19, 22, -26, -60, 0, -31, 27, 35, 54, 15, -15, 41, -46, -44, 20, -37, -25, 43, -37, -10, -31, -13, 11, -39, 93, 15, 25, 40, -61, -7, -23, 41, 26, 68, -12, -43, -10, -63, -48, -42, 31, 29, 19, 38, -31, 7, -45, 32, 78, -28, 46, -11, -100, -49, -55, -23, 66, 90, 49, 29, -73, -22, -76, -15, 21, -51, 66, 25, -36, 23, -47, -77, -3, 38, 79, 23, 0, 54, -25, -29, 41, 14, -48, -4, -64, -30, 8, 11, 32, 49, -43, 17, -3, 59, 61, 44, 31, -47, -40, -69, -128, -13, -30, -18, 7, 20, -10, -22, 19, 66, 90, 63, 60, -4, -69, -30, -35, -12, -15, -31, -28, 28, -23, -30, 70, 0, -32, 18, 4, -36, 14, 124, -17, -32, -11, -25, -19, 5, 8, 15, -14, 7, 82, -37, -24, 55, -32, -41, 3, -32, 17, 19, 1, -43, 9, -5, 20, 57, -69, -2, -35, 28, 91, 40, 2, -21, -25, -32, -88, 0, -41, -49, 22, 28, 73, -15, -11, 31, -62, 8, 85, -3, 38, 62, -8, -22, -22, -61, -6, 26, 34, 64, 28, 5, -56, -23, -58, -98, 45, 7, 11, 32, -27, -47, 11, -2, 31, 42, 1, -8, 32, 56, 34, 58, -18, -37, -66, -53, 15, 72, 10, -2, -10, -26, -81, -17, -1, -22, 59, 31, 25, -10, -122, -49, -30, 30, 80, 36, 15, -15, -32, 0, -5, 24, 69, 4, -9, 9, 13, -14, 47, 7, -32, -63, -7, -27, 26, -39, 22, -25, -15, 41, -28, 45, 44, -6, 24, 4, -55, 46, 23, -8, 37, -22, -39, 10, -97, 4, -7, 6, 78, 2, -27, -10, -22, -55, 44, 20, 19, 30, 13, -46, -26, -71, 40, 32, 31, -26, -41, -64, -62, -11, 76, 109, 58, 100, 18, -45, -17, -100, -72, -19, -19, 40, 55, -22, 18, -59, -2, 70, -32, 1, 40, -1, -12, 37, 21, -45, 9, -12, -88, -5, 9, 76, 91, 102, 27, -32, -36, 7, -49, -30, -31, -42, -39, 42, 6, -34, 74, 44, -2, 43, 0, -37, -4, 7, 22, -8, -56, -10, 42, 0, 66, 38, 14, -89, -72, -43, -24, 60, 47, 55, -32, -55, -9, -57, -34, -23, -21, 24, 46, 0, 28, -37, 23, -24, 18, 72, -17, 21, -1, -64, -59, -34, -14, -36, 38, 0, -18, 4, 52, 17, 58, 53, 11, 21, -62, -25, -29, 30, 59, 58, 31, -64, -29, -51, -63, -26, -15, -52, -2, 37, 0, -17, 60, 47, -12, 9, -8, -72, 45, 39, 53, 4, 6, -12, -40, -31, -17, -10, 63, 26, 22, 26, -30, -7, 23, -19, 3, -12, 38, -7, 63, 8, -2, -3, -45, -15, 29, -43, -1, 22, 14, -59, 30, -10, -59, 49, -3, 30, 30, 53, -12, 8, 13, -89, -45, -14, -19, 41, 39, 59, -9, 47, 34, 23, 26, -45, -25, 18, -23, 40, 0, 10, -28, 20, -7, -1, 11, -49, 34, 26, -10, 11, -26, 2, 3, 8, -8, -6, -47, -4, 24, -32, -20, -35, -66, 39, 34, -24, 7, -53, -52, 13, 46, 96, 34, 64, -13, -31, -3, -36, -14, 24, -53, -8, -26, 28, 51, 19, 21, -2, -85, -52, -3, -15, 11, -42, 77, 44, 39, 72, -13, -23, -30, -59, 30, -6, 48, 8, 15, 62, -25, -26, -64, -64, -77, 5, 95, -9, -7, -3, -21, 17, 25, 75, 11, -2, 26, 47, -8, 19, -49, 0, 36, -21, 37, -23, -89, -31, -73, -34, -26, -21, 14, 72, 75, 51, 28, 42, -48, -52, -8, -4, 18, 45, 30, 20, 14, -10, 23, -30, -18, 49, -8, 0, -40, -69, -38, 66, 4, -3, -19, -34, -45, -11, 54, 43, 7, 49, -37, -13, 8, 35, 75, 66, 10, -31, -10, -4, -76, -38, -63, -103, -23, 69, 95, 83, 82, 20, -36, -65, 2, -37, -35, 1, 41, -32, 8, 6, -83, 15, 42, -10, -8, -6, -48, -34, 0, 70, -15, -3, 99, 31, 29, 54, -9, -38, -5, -19, -19, -3, 40, -15, -18, -13, -79, -82, 64, 54, -14, 15, 10, -88, -66, 45, -4, -2, 0, 21, 13, -25, 49, 99, -8, 12, -28, -40, 6, 0, 7, 49, -71, -68, 26, 23, 22, 20, 1, -7, -85, -41, 1, -19, 53, 26, -7, -23, -40, -14, -6, 55, 44, 1, -10, 30, -35, 23, 44, 23, -17, -10, -29, -54, 95, 40, 48, 40, -34, -27, -26, 1, -7, 17, 51, -66, 28, 52, -71, 21, -17, -49, -63, -28, -53, 20, 56, 4, -1, 35, -77, 6, 65, -46, -5, 22, 21, 21, 86, 43, 0, 1, -65, -43, -10, 42, 48, 88, -19, -113, -57, -41, 47, 32, 20, -11, -110, -20, -17, 21, 77, 61, 39, 79, -18, -14, 0, -19, 55, -24, -2, -21, -99, -11, -7, 44, -25, 24, -19, -79, 25, -1, 12, 22, -31, 32, -3, 0, 41, 74, 9, 4, -41, -62, -52, -27, -12, 81, -39, -38, 10, -53, 11, 91, 35, 70, -17, -88, -19, -20, 25, 35, 19, -39, -43, 24, -15, -43, 30, -17, -3, 69, 3, -2, -73, -6, 2, 58, -1, 0, 27, -4, 22, 28, -75, -44, -96, -14, 81, 62, 39, 40, 37, -34, 29, 2, 31, -25, 40, 6, -27, -9, -11, 41, -23, 11, -23, -61, -49, -4, 45, 0, 53, 38, -4, 20, -6, -28, -88, 30, 34, 6, 17, -28, -41, -24, 30, 60, 12, -19, -21, -36, -11, 13, -9, 59, -1, 30, -56, 9, -32, -73, 80, 41, 37, 39, -64, -48, -42, -17, 87, 46, -36, 3, -15, -61, 54, 17, 22, -30, -9, -3, -44, 80, 55, 63, 2, -23, -19, -96, 6, 37, -53, 28, 7, -46, -12, 6, 1, -13, 22, 36, -27, -58, -8, -85, -44, -28, 32, 73, 72, 41, -30, 5, -10, 9, 75, 45, -51, -4, -62, 0, 40, 20, 44, 40, -72, -26, 9, -59, 35, 39, -49, -2, -36, -9, 18, -20, 69, 48, -27, -2, -9, -39, -62, 12, -32, 29, 72, 65, 56, 22, 21, -11, 7, -26, -81, -65, -44, -11, -51, 43, 21, 43, 11, -11, -35, -48, 17, 68, 44, 5, 5, -63, -8, -69, 15, -6, -9, 21, 26, 3, 73, -7, -9, 7, -1, -44, 22, 21, -61, 54, -5, 0, 20, -28, 10, -37, 9, 8, -53, 64, 32, -5, 56, -60, -23, -7, 56, 49, 15, -14, -9, -41, 5, 52, 32, -15, -23, -55, 12, -21, -37, 49, 15, -1, 71, 39, -12, 10, -6, -32, 53, 13, -38, -3, -28, -88, 7, -41, 23, 35, 68, 71, 47, -7, -74, -82, -78, -29, -10, 15, 17, 17, 28, -52, 12, -8, -14, 0, -6, 47, 41, -3, -5, -12, -45, -17, 48, 125, -9, 30, 22, -43, -30, -23, -107, -21, -57, -19, 86, 22, -43, 54, 10, -39, 12, 20, -72, -30, 93, 22, -3, 5, -56, -80, 22, 2, -26, 45, 11, 44, -2, 58, 8, -95, 48, 37, -58, 42, 1, -112, -17, -21, -26, 57, 65, 82, 14, 44, 19, -74, -68, -3, -73, -51, 94, 48, 0, 82, 28, -57, -3, -35, -73, 22, 20, 38, 11, -63, 2, -36, -23, 7, -2, -14, 39, 19, -27, 6, 11, 15, 24, 22, 34, -32, 37, 34, 7, -19, -8, -62, -27, -27, -19, 60, 60, -1, -18, 2, -60, -36, 91, 5, 9, -2, -23, -10, -9, 66, -11, 40, 47, -66, -15, 21, -86, -44, 35, -44, 21, 62, 90, 61, 58, 31, -41, -44, -51, -78, -29, 23, -14, 8, 29, -19, -28, -22, -9, 32, 10, 27, 35, -65, -14, -2, 0, 4, 40, -46, 30, -62, 7, -6, -10, 54, 34, 91, 45, -6, -38, -13, -29, -47, 39, -7, -48, 53, -60, -3, 26, 5, 19, 29, -32, 10, 10, 49, -2, -29, -66, -82, -49, 27, 49, 17, -22, -12, -45, -5, 55, 48, 66, -42, -34, -45, -45, -21, 58, -6, 35, 18, -57, 7, -20, -17, 30, 58, 61, 14, 15, -49, -87, -25, -6, -1, 104, 36, 2, 8, -19, -78, 0, -5, -2, -1, 71, -15, -2, -30, -52, 20, -20, 6, 65, -2, 17, -9, -31, -70, -49, -63, -2, 41, 64, 54, 98, 14, 14, -46, -14, -23, -126, -8, -17, -1, -7, 71, 23, -10, 99, 54, 8, 9, -10, -88, -6, 36, -54, 12, -7, -109, -9, -32, -14, 68, 76, 9, 51, 21, -23, -12, -56, -25, -51, -40, 63, -2, 0, -36, -48, -46, -4, 45, 39, 65, 37, 23, -10, 26, -95, -3, 19, -20, 64, 120, 2, -2, -12, -40, -77, 25, 8, -47, 61, 0, -59, 18, -6, -18, -5, -2, -2, -8, -35, 69, 36, 9, 44, 34, -12, -23, -64, 22, 18, -5, 52, -26, -46, -15, -27, 46, -53, 38, 48, -38, 38, 25, -38, -13, 20, -48, -21, -10, -14, 61, 24, -3, 43, -29, -90, 4, -53, -10, 0, 61, -23, 42, 70, -26, 35, 10, -63, 45, -3, 23, 14, 23, 29, 44, 2, -41, -43, -62, -120, 13, 2, 27, 61, 122, -30, -42, -46, -86, 36, 54, 59, 52, 0, -41, -14, -24, 78, 6, 49, -9, -68, -72, -94, -53, -26, -10, 35, 34, 0, 63, 34, -32, 21, 42, -58, 11, 41, -36, 81, 5, 0, -7, -21, -7, 24, 96, -24, -43, -44, -74, -20, 59, 24, 11, -7, 21, -15, 13, -38, 7, -18, -18, 91, 46, 17, 40, -6, -48, -18, -28, -55, 57, 3, -8, 57, 39, -42, -27, -79, -68, -13, 80, 54, 58, 11, -4, 42, 47, 19, -25, -65, -89, -27, -23, 3, -3, 38, -8, -17, 83, 24, 25, 41, -30, 0, -92, -35, -3, -56, 0, 5, 89, 58, 56, -6, -42, 7, -6, 56, 91, 11, -10, 13, -59, -53, -23, -35, 23, 22, 56, 10, 42, -37, -17, -49, -91, 0, 54, 37, 11, -49, -54, -64, 37, 48, 54, 30, -65, -6, -36, -8, 5, 13, -3, 9, -61, 62, -13, -36, 71, -27, 4, 88, 10, 39, 60, 0, -10, -17, -37, -74, 54, -6, -20, 26, -23, -35, 55, -10, -37, 8, -63, 37, 57, 26, 80, -7, -24, -45, -85, -9, -17, 4, 90, 0, -24, -7, -93, 9, 14, 8, 119, -10, 25, 35, 10, 21, 0, -38, -55, -35, 23, 20, 66, 20, -31, -9, 10, -15, -18, 37, -18, -68, 32, -20, -27, 36, 5, -26, 22, -29, 35, 81, 9, -10, -36, -71, -51, -34, -8, 5, 4, 88, 36, 27, -52, -7, -7, 51, 46, 45, -27, -86, -35, -42, 1, 74, -8, 0, -20, -56, 6, -14, 61, 18, 10, 5, -14, -62, -32, -68, 26, 68, 21, 49, 77, -48, -20, 51, 8, 8, 25, -77, -75, -98, -20, 60, 76, 52, 61, 14, -31, 47, -11, -71, -48, -6, -14, -56, 10, -29, -45, -11, 57, 89, 20, 60, 71, -78, -75, -35, -27, 45, -4, 46, 56, -15, -3, -19, -15, -32, 2, 86, 72, -27, -3, -17, -68, 36, -3, 1, 27, -53, 1, -8, 64, -29, -30, -9, -72, -83, 39, 47, 62, 36, 18, -26, 31, 21, 63, 43, -3, -29, -61, 0, -1, 17, 0, 2, -53, -73, -17, 34, 40, 35, -37, 10, 34, 15, 17, -45, -51, -55, -4, -5, 4, -64, -48, -18, 39, 56, 32, 25, 5, -18, -10, 3, -34, 60, 55, 8, 28, -31, -64, -66, 1, 13, 11, -32, 45, 31, 35, 30, 5, -32, -21, 32, 9, 4, -19, -14, -40, -11, -5, -28, 30, 49, 12, 60, -6, -59, 7, -15, -22, -36, 2, -6, 69, 20, 43, 20, -78, -14, -8, -44, -6, 44, 23, 2, -17, -31, -61, 23, 22, 39, 61, -1, 34, -34, -21, -61, -41, -21, -9, 4, 38, -1, -25, -30, 24, 58, 72, 115, 47, -26, -54, -34, 66, -21, 12, -32, -97, -38, 25, -24, -2, 0, -46, 27, 18, 8, 24, -42, 44, 11, -28, -8, 0, -41, -42, -7, -10, -29, -34, 82, 25, 7, 59, -4, -12, -95, -17, -28, 22, 97, 12, 29, -11, -48, -8, 21, 73, -42, 40, 24, -78, -44, -52, -77, -35, 61, 97, 7, 6, -4, -108, -41, -18, 25, 23, 35, 25, 3, 21, -65, -10, 25, 8, 45, 106, -24, -28, -51, -97, 0, 30, 25, 27, -24, 17, 22, 61, 61, 11, -63, -35, -31, -9, -12, -35, 5, -5, 28, 109, -23, -12, 9, -4, -37, -1, 27, -93, -49, 23, -35, -25, 34, 47, -8, -8, 63, 44, 27, 70, 11, -32, -32, -32, -36, -60, -25, -55, 6, 49, 36, 40, -4, 7, 41, 31, 47, -5, -66, -98, -31, -39, -43, 39, 40, 41, 31, 64, 22, -23, 7, -11, -32, 25, -41, 0, 29, -86, 17, 56, -7, 95, 59, -10, 9, -18, -83, 21, 23, -26, 26, 62, -54, -35, -19, -11, -48, -10, 20, -77, -20, -35, -14, 93, 92, 59, 69, 9, -60, -30, 40, -26, -36, -34, -52, -71, -51, 4, -44, -2, 61, 4, -5, 26, 13, 30, 27, 13, 35, -13, 74, 6, -46, -55, -64, -45, -26, -22, 9, 22, 49, 29, -25, 8, -44, -35, 42, -23, -37, 51, -23, -42, 44, -21, 14, 65, 9, 37, -71, -17, -65, -58, -19, 24, 85, 82, 48, 3, -15, -31, -24, 1, -57, -34, -23, 10, 60, 88, 19, 10, 11, 18, 17, 58, -31, -76, -29, -48, -11, 22, 31, -45, -26, 62, 18, 28, 37, -45, -32, -22, -19, 15, 45, -26, 6, 38, -21, -38, 12, -31, -74, 61, -8, -47, -31, -52, -19, 34, 10, 57, 2, -47, 63, 8, 52, 46, 52, 5, -7, -38, -62, -1, -82, -20, -15, -39, 27, 10, 55, 2, 42, -13, 46, 47, -5, 25, -45, -40, -87, -25, 28, 64, 35, 40, 40, -19, 18, 30, 46, 12, -44, -17, 8, -14, 69, 37, 17, 8, -19, 22, -26, -69, -29, -47, -40, 77, 39, -9, -44, -52, -43, 18, 44, 97, 22, 11, -5, -19, 0, -14, 20, 6, -39, -25, 34, -29, -11, -2, 1, 12, 1, -5, 7, -70, -74, 35, 32, 0, 45, -2, -88, -6, 9, 68, 90, 31, 8, 17, -66, -37, -24, -14, -55, 4, 56, -56, 7, 44, -32, 22, 22, -32, 5, -40, -42, 0, -32, -3, 4, 36, 48, 22, 57, 17, 12, -6, 0, 40, -27, 47, 12, 15, -24, -21, -95, -62, -32, -26, -10, 26, -31, 54, 17, -24, 52, 0, 13, 53, 19, -46, -34, 12, 42, 14, 27, 15, -44, 0, 9, 32, -43, -62, 51, 11, 26, 39, 18, -19, -56, 51, -40, -64, 9, -7, -43, 47, 27, -78, 46, 46, 21, -3, -11, -56, -85, -37, 45, 69, 54, 103, 4, -63, 1, 0, -28, 3, 39, 13, 11, 32, -37, -89, -63, -70, 46, 65, 52, 96, -27, -52, 35, 3, 55, 73, 31, -4, -62, -58, -64, -76, -63, -1, -30, -9, -17, 31, 53, 61, 34, 63, 14, 34, 3, 29, -10, -68, 15, -10, -31, 7, 18, -10, -4, -28, 56, 6, 44, 30, -37, 7, -14, 3, 7, 22, -22, -60, -8, -35, 28, 20, 51, 2, -31, 0, -40, 15, 72, 25, 2, -26, 2, -30, -17, 82, 28, 26, 5, -35, -59, -80, -62, -13, 38, 55, 28, 41, 51, -19, 44, -14, -28, 2, -78, 20, 9, -48, -6, 1, -23, -65, 12, -52, 40, 73, 54, 62, -32, 0, -40, -46, 9, -47, -18, 34, 5, -20, 51, 6, 17, -24, -32, -47, -59, 36, 127, 44, 79, 20, -56, 5, -90, -74, 29, 11, 36, 98, -22, -89, -51, -69, 17, 57, -22, 11, -48, -7, 10, 80, 66, -14, -30, 6, -98, -53, 52, -31, -12, 52, -34, 20, -6, -4, -8, 25, 28, -4, 30, -28, -56, -45, 7, -5, 5, 46, -5, 99, 34, 58, -28, -78, -17, -1, 26, 74, -7, 2, -22, 0, -5, -41, -23, -23, 24, -21, 80, 51, 20, 57, 14, -46, -40, -57, -46, -45, 24, -11, 56, 19, -11, 69, -47, 36, 43, -25, 31, -19, -79, -41, -8, 21, 9, 26, 27, -18, -44, 30, 42, 38, 58, 40, 4, -14, -59, -34, -37, -89, -25, -9, 19, 58, 48, -2, 28, 63, -79, -49, -32, -59, 1, 0, 32, 26, 5, 61, 48, 20, -30, -75, -52, -60, -48, 32, 56, 43, 71, -9, -40, -11, -58, 0, -32, -44, 6, -1, 24, 89, 64, -14, -23, -2, -17, -38, 68, 25, -35, -9, -21, -18, 2, 35, -62, -14, -5, 0, -5, 48, 23, 11, -6, 37, 9, -2, 9, 2, -28, -75, -55, 26, 44, 48, 54, -13, -69, 32, -23, -53, 6, -11, 9, -15, 24, -29, -39, -58, 13, 60, 32, 30, 38, -6, 25, -13, 42, -36, -20, -25, 7, 42, 43, 61, -43, -44, -32, -76, -27, 37, -32, 52, -31, 5, 36, -75, 2, 17, -36, 23, 80, 74, 29, 60, 35, -42, -52, -18, -21, 7, 1, -23, -11, -73, -42, -62, 40, 42, 45, 69, -44, -54, -87, -44, 25, 28, 5, 66, -44, -15, 7, -7, -26, 22, -39, -20, 8, 12, 5, 80, 29, -30, -30, -6, -15, 42, 59, 77, -22, -9, 27, -26, 21, -19, -1, 7, 7, -17, -3, -60, -76, -22, 6, 49, -9, 41, 11, -77, 65, 40, 15, -6, -68, -40, -14, 12, 19, 88, -15, -48, -3, -86, -89, -44, -10, 32, 61, 52, 21, 9, 45, 0, 6, -8, -4, -21, -68, 31, -31, -34, -6, 19, 12, -38, -8, 46, 42, 91, 97, 12, -42, -59, -99, -44, 13, 30, -10, -20, 6, -39, -13, 19, 12, -2, -25, -13, 57, 29, 54, 7, -3, 3, -11, 49, -39, -53, -31, -65, 28, 104, -14, 24, 37, 15, 31, 60, 14, -5, -25, 0, -36, -57, 10, 4, -34, 32, 34, -71, 0, -7, -49, 68, -5, 4, 23, -12, -56, 15, -73, 0, -6, 36, 73, 9, -31, 13, -22, 34, 14, 31, -3, -64, -21, 0, 46, 28, 48, -40, -66, -35, 11, 11, 23, -45, 5, -1, 0, 49, 11, 25, 39, 35, -23, -12, -19, -86, 38, 10, -23, 26, -2, 30, -69, 12, 22, -11, 4, 66, 26, 17, 55, -25, -97, -39, -80, -41, 32, -15, 7, -30, 59, 56, -9, 4, -47, -17, 19, -9, -4, 2, -39, -1, 30, 2, 14, -13, 49, 4, -21, 18, -10, 40, 73, 21, 54, 2, -38, -53, -74, -39, -48, 23, -4, 7, 0, -24, 37, -10, -80, 22, -26, -18, 68, 86, -35, 32, 37, -75, 57, 58, -24, 23, -4, -65, -3, 35, 7, 97, 13, 2, -36, -26, -60, -64, 23, -39, -21, -1, -53, 49, 48, 26, 68, 14, -11, 9, 11, 3, 49, -57, -17, -5, -80, -19, 5, -20, -5, -14, 6, 17, 65, 27, 73, 52, -31, 5, 42, -23, -21, -29, -74, -54, 5, 78, 0, 3, 45, 8, 31, 32, 18, 21, -45, -26, -55, -8, 17, 48, 86, -35, -72, -43, -17, 35, 44, 12, -99, -26, -46, -12, 79, 28, 49, 94, 15, 62, 25, -47, -68, -27, -31, -41, 76, -22, -2, 6, -109, 8, 0, -28, 56, 1, -80, 18, 3, 0, 53, -42, -3, 9, 31, 42, 31, 32, 13, 4, -21, 17, -6, -57, 10, -7, -34, 5, 3, 52, 30, -37, -3, -34, -48, -25, 26, -4, -2, 19, -44, 35, -21, 7, -15, 37, -3, -8, 88, -46, -15, 36, -17, 56, -13, -49, 17, -34, 12, 127, 3, -17, -58, -21, -70, -24, 31, -46, 48, 22, 49, 28, -20, -25, -103, -49, -42, 22, 46, 26, 35, -9, -41, -57, 61, 7, -26, 73, -7, -70, 34, 21, 24, -5, -13, -65, -63, -17, 55, 30, 52, 46, -55, -63, -8, -4, 49, 75, 32, -32, 19, 15, 41, 66, 9, -78, -71, -27, 34, 21, 12, -23, -18, -48, -1, 63, 5, 18, 51, -27, -28, 6, -43, 29, 62, -39, -7, 23, -22, -11, 30, 20, -61, -27, -20, -52, 4, 30, 55, 21, 44, -30, 6, 10, -4, -4, 44, -49, 13, -18, -86, -11, -15, 35, 75, 32, 14, -41, -51, 12, -1, -36, 73, 31, -35, 57, 31, -120, -46, 9, -44, 1, 86, -35, 0, -29, 19, 48, 36, 99, 36, -39, -43, -65, -80, 19, -15, 36, 62, -35, -51, -24, -89, -4, 5, -21, 69, 43, -26, 38, 61, -13, 18, 62, -4, -19, -69, -77, -42, 23, 80, 55, 24, -47, -63, -5, 37, 24, 81, 10, 11, 83, -4, -20, -47, -53, -71, -27, 45, 38, 49, 66, -8, 0, 4, 6, -58, -52, -29, -21, 32, 112, 74, 23, -1, -75, -94, -89, -75, 1, 70, 57, 5, 3, -32, -62, 4, -5, 8, 27, 75, 5, 13, -7, 14, 7, -2, -48, -49, -60, -2, 20, -27, -15, -3, 38, 63, 44, 20, 34, -37, 6, 51, -39, -44, -19, 11, -51, -5, 90, -8, -22, 59, 43, -63, 38, 9, -115, -9, 39, 25, 48, 20, -25, 14, -18, 25, -20, -28, -64, -23, -27, 6, 56, 29, 43, 79, -17, -52, 9, 12, -60, -21, 18, -43, 2, 25, 24, 4, -38, 3, 18, -27, 69, -5, 2, -38, -86, 23, 5, -7, 74, -14, -21, 35, -53, 22, 35, 7, 72, 79, -9, 7, 3, -47, -31, -71, 8, -61, -39, 14, -36, 5, 62, 72, -3, -2, -31, -105, 19, -8, -22, 53, 49, 3, 44, 49, -32, -55, -27, -81, -80, -23, -11, 40, 45, 17, 12, 22, 0, -6, 22, -9, -82, 44, -2, -12, 91, 10, 3, -42, -17, -37, 56, 64, 29, -19, -7, -56, -57, 21, -102, -59, -60, -40, -1, 20, 38, 34, 18, 10, 21, 30, -18, -1, 28, -20, 3, 59, -14, -15, -12, -24, -47, -36, 31, 11, 15, 97, 35, 36, 35, -2, -29, -2, -89, -13, -23, -95, 61, 45, 38, 78, -9, -23, 15, -56, -29, -34, -44, -10, 4, 70, 32, 52, 36, 41, 15, 18, 5, -11, -61, 1, -26, -64, 1, -30, 1, 61, 14, 43, -31, -81, 36, 32, 21, 81, 9, -49, -17, 45, -66, -3, 24, -82, -36, -6, -54, -46, 18, 29, 44, 51, 55, 30, -53, -3, 5, -89, -17, 27, -31, 30, 83, 31, 26, -7, -75, -21, -79, 29, 88, 11, 53, -21, -100, 14, 20, -9, 36, -27, -98, -8, -45, -17, 52, -21, 7, 96, -2, 19, 82, -14, 14, 54, -74, -94, -24, -30, 49, 86, 61, 11, -52, -7, -20, -4, -62, -31, 2, -10, 53, 74, -45, 15, -6, -40, 64, 21, -2, -37, 41, 1, -3, 60, -12, -25, 2, -38, 30, -48, -65, 44, 25, 14, 75, 21, 24, -69, -34, 8, -45, -21, 97, -18, -11, -39, -60, -71, -37, -19, -19, 32, 0, 40, 83, 77, 92, 77, 27, -52, -75, -26, -36, -32, 51, 52, -40, 38, 60, 1, 48, 52, -27, -69, -22, -34, -25, 47, -49, 22, 17, -54, 7, -14, -29, 13, 35, 7, 43, -83, -7, 3, -47, -12, 69, 35, 7, 70, 21, -61, -56, -51, -13, -42, -36, 27, -11, 31, 35, 62, 4, -12, 59, -10, 4, 57, 7, -34, -27, -13, -57, -55, 66, -48, -28, 68, 24, 45, 107, 2, -69, -46, -19, -21, 21, 32, 47, -75, -26, 5, -38, -44, 7, 13, -17, -24, 92, 37, 43, 87, 42, -30, -26, -9, 4, 4, 54, 11, 18, -9, -32, -80, -52, -9, 2, -14, 0, 9, -10, -59, 27, 24, 15, 55, 38, -5, 18, -9, 65, 3, -32, 11, -42, -18, 7, 44, -20, -21, 56, 22, -56, 32, 48, -93, -36, -9, -64, 5, 59, -6, 23, -7, -110, 1, -27, -5, 23, 42, 76, 24, 6, -62, -28, -21, 35, 54, -7, -44, -72, -18, -3, 0, 7, -71, -28, -46, -1, 32, 31, 21, 8, 46, 20, 64, 71, -3, 14, -22, -45, 14, -20, 6, -47, -19, -31, -51, 52, 68, 40, 38, 43, -31, -22, -15, -93, -42, -8, 14, 13, 47, 39, 2, 38, 37, 5, 7, -13, -22, -94, -53, -79, -20, -6, 0, 56, 32, 2, 68, 46, -40, -21, 5, -71, 10, 62, -45, -10, -59, -9, 13, -7, 86, 9, -70, 9, 17, 11, -2, 43, -40, -13, -21, 25, -39, 66, 9, 1, 26, -12, 15, -70, -37, -31, -41, 4, 34, 98, -41, 4, 14, -40, -23, 21, -17, 17, 17, 66, -10, -37, 34, -41, 29, 22, -20, 22, 0, -63, 4, 11, -15, -13, 25, -46, -95, 11, -4, 3, 76, 36, 3, -24, -38, -11, -18, 76, 90, 45, 64, -32, -55, 4, -1, -34, 10, -9, -62, 48, -5, 5, 49, 8, 47, 55, 0, -81, -77, -87, -53, 17, -13, 29, -14, 0, 18, 27, 40, 76, -39, -26, -9, 1, 56, 11, -23, -19, -25, 25, 114, 73, 14, -48, -78, -63, -64, 31, -6, -12, -44, -28, -12, 29, 46, 59, -64, -47, -39, -19, 24, 8, 36, 38, -2, -3, 58, -1, -41, -9, -49, -20, 34, 46, 92, 36, -43, -68, -55, -47, 19, -32, -17, 29, -4, -5, 90, 13, -31, 25, -32, 13, -35, -28, -11, -20, 0, 29, 83, 23, 110, 29, 21, -28, -77, 0, 4, 63, 83, 29, -52, -56, -22, -127, -22, 14, -10, 58, 76, 42, 23, 0, -28, -98, -19, -11, 14, 0, -13, -15, 18, 45, 20, 17, -15, -107, -43, -28, -8, 45, 22, 30, 35, -58, 5, 55, 2, 3, 42, -36, 38, -20, -10, 28, -64, 18, 9, -59, 23, -46, -12, 9, 74, 56, 80, 76, -36, -60, -5, 9, 21, 79, -14, -32, 35, -65, -47, -35, -48, -53, -8, 57, -11, -42, 12, 15, 18, 30, 20, -41, -20, 10, -5, -12, 34, -37, 3, 57, 65, 1, -39, -6, -11, 15, 59, 62, 49, -30, -4, -1, -72, -56, -7, -8, -19, -13, -6, 10, -14, -7, 62, -18, -15, 51, -53, 32, 18, -23, 43, -64, 13, 20, -31, -28, -13, -20, 18, 60, 90, 31, -4, -49, -69, -24, -31, 8, 29, -29, -9, -59, 23, 11, -62, -1, -18, 21, 51, 26, 39, -26, -39, -11, 42, -1, 4, 38, 5, 65, -30, 2, 28, -77, -38, 0, -74, -43, 0, 57, 23, 37, 28, -52, 17, -32, 41, 40, 40, 88, 30, 11, -9, -45, -37, -30, -38, -52, 13, 10, -45, 32, -6, -15, 11, 17, 2, -71, 37, -5, -49, 76, 19, 12, 83, 52, -5, 18, -29, -93, -42, -41, -35, 0, 58, 19, 80, -34, -15, 5, -59, -28, 57, -8, -7, 3, 0, 12, 47, 5, 17, -69, -9, -10, 18, 62, 59, -36, -34, -17, -59, 54, 24, 38, 62, 12, 3, -6, 7, -29, -62, -26, -99, -26, 10, 12, 8, 89, 21, 35, -2, -47, -69, -71, 17, 54, 81, 43, 23, 45, 12, 10, 14, -43, -104, 38, 22, 48, 99, 25, -8, -18, -54, -35, -46, -45, -42, -27, -62, 10, 25, 53, 80, 48, 29, 56, -13, -6, -9, -80, -63, 0, -35, -1, 44, 72, -9, 0, -48, -75, -49, 4, 77, 96, 22, 60, 46, -65, 14, 51, -22, 17, 23, -37, 8, 22, -32, 0, -10, -89, 42, 9, -3, 29, -39, -18, 9, 21, -4, 9, 2, 52, 19, 23, -38, -109, -79, 8, 54, 6, 62, 0, -85, 55, 20, 41, 7, -39, -13, -96, -19, 55, 62, 56, 21, -17, -22, -120, -19, -19, -28, 24, 3, 56, -26, 10, -8, -53, -10, 13, -19, 24, 35, -47, 32, 44, -23, 51, 54, 2, 25, 4, -42, -46, -55, -29, 45, 64, 54, 55, 12, -66, -59, -65, 19, 45, 32, 96, 32, -15, -6, -9, -52, 28, 29, 3, 8, -30, -62, -25, -10, -15, 19, -30, -12, 32, 74, 49, 65, 17, 0, -18, -37, 13, 8, -82, -19, -42, -85, -13, 24, 11, 9, 31, -63, 0, 6, 83, 13, 14, 22, -26, -12, -30, -22, -12, -23, 41, 98, 6, 23, -47, -88, -1, 23, 73, 90, 68, -7, -52, -39, -30, -22, 47, 1, -27, 28, 9, -45, -3, -76, -77, -42, -2, 34, 51, 71, 5, -6, 21, -23, -29, 51, -22, -24, -47, -26, -70, 1, 52, 69, -3, 25, -20, -93, 5, 9, 31, 28, -1, 37, -49, 19, -34, 69, 29, -19, 6, 32, -2, -12, -6, -20, -89, -62, 71, 18, -18, -4, -27, -51, 7, -7, 46, -7, 59, 38, 4, 37, -5, -53, -3, -22, 10, -7, -7, 18, 13, -42, 34, -45, 7, 15, -14, 37, 42, -44, 32, 69, -59, -10, 22, -14, 26, 41, -9, -19, -108, -30, 40, 51, 90, 71, -5, -59, -39, 44, -22, 41, 17, -83, -59, -4, -24, -25, 107, 26, 51, 42, -53, -88, -19, 0, 58, 89, -7, -55, -62, -40, 25, -36, 11, -35, -63, 44, 6, -22, 26, -53, -6, 18, 58, -17, -45, -26, -15, 34, 38, 73, 26, -77, 11, 8, 1, 10, 13, -61, 41, 4, 23, 74, -12, 10, 8, -29, -30, 0, -18, -81, 29, -12, -56, -1, -11, -23, 17, 104, 70, 105, 28, -55, -52, -32, -25, -13, -42, -13, -69, 6, 75, 34, 81, 57, -42, -10, 22, -91, -35, 12, -65, -47, 61, -26, -10, 74, 13, -12, 74, -19, -46, 39, -29, -35, -42, -48, 11, 65, 56, 65, -8, 12, -49, -45, 27, -23, -10, 90, -32, 23, -7, -66, 80, 31, 29, 12, -54, -59, -25, 37, 43, 26, -4, -85, -52, 19, 13, 41, 41, 11, -24, -51, 27, -17, -1, 20, 49, -3, -29, 48, -2, -18, 72, 13, -35, -37, -21, -70, -20, 13, -39, 77, 36, 5, 11, -22, -99, -25, -2, 1, 9, 83, 42, 3, 3, -24, -42, -34, 25, -10, -57, -5, 6, 40, -12, 62, 12, -81, 19, -38, -30, 10, 9, -45, 27, 27, 22, -4, -15, -25, -23, 25, 14, 56, -23, -24, -37, -27, -52, -5, -23, -18, -2, 28, 47, 9, 35, 0, -35, 69, 13, 24, 0, -41, 25, 27, -13, -38, -42, -37, 48, 56, 63, 0, -66, -72, -10, -6, 32, 54, -46, -10, -40, -57, 10, -23, -10, 6, -35, 10, -26, 9, 45, 65, 58, 54, 41, -46, -73, -43, -71, -40, 35, 48, 40, 57, -44, -59, -20, -25, 6, 28, -25, 46, 11, -4, 62, 0, -31, 31, 31, 3, 4, -37, -21, 1, -63, 23, -19, -6, -54, -31, -31, 0, 57, 65, 58, -7, 21, 26, -25, 46, 64, -35, 14, -22, -73, -90, -54, -55, -58, -1, 48, 88, 46, 32, -56, -102, -80, -41, 4, 6, 9, 47, 30, 31, -11, 55, -18, -47, 77, -39, -35, 49, 42, 48, 59, 8, -72, -49, -37, -56, 35, -35, 20, 46, 15, 51, 21, -3, -87, -20, -14, -7, 10, -27, -41, -70, -25, 0, 52, 77, 15, 1, 1, 3, -24, -38, 25, -2, -8, -8, -12, -37, -64, -35, 7, 5, 40, 29, -12, 54, 18, -10, 32, -12, -1, 3, 76, 43, -4, -86, -83, -116, -40, 3, 6, 36, -7, 15, 64, 80, 60, 21, -22, -45, -41, -5, -46, 31, 20, 4, 5, 51, -12, -73, -49, -53, -59, 3, 32, 74, 3, -77, 3, -58, -35, 71, 45, 0, 13, -2, 0, -2, 56, 22, 26, 71, 6, 58, 36, -13, -19, -44, -36, -14, -18, 7, 36, -2, 22, 49, -35, -29, -10, -48, -3, -9, -62, 21, -11, 5, 70, -5, 17, 71, 24, 54, -35, -69, -46, -66, -19, -6, 32, -14, -38, 44, 28, 15, 60, 44, 40, -19, -13, -48, -26, -41, 73, -8, -3, 3, -69, -37, 0, 29, -23, -43, -4, -65, 12, 73, 49, 57, 17, -51, 7, -7, 53, 52, 30, -6, -48, -55, -95, -6, 48, 27, 44, 42, -57, -114, -21, -29, 25, 72, 53, 66, -11, 39, -11, 42, 9, -53, -62, -74, -83, -35, -5, 41, 18, 15, 96, 20, 85, -5, -42, -36, -59, -46, 43, 8, 4, 38, -78, 1, -31, -15, 78, 30, 47, 74, -2, 4, -20, -6, -85, -5, 28, 19, -18, 34, 28, -76, 38, 52, -83, 19, 27, -17, 92, -14, -28, -9, -69, -17, 35, -85, -24, -12, 20, 40, 41, 17, -42, -35, 13, 58, -20, -2, -25, -96, -44, -19, 35, 62, 58, -26, -19, -19, 6, 38, 71, 0, -111, -48, -3, 35, 24, 59, -9, -43, -14, 26, -6, 45, -8, 20, -2, -21, -17, -91, -15, 1, 56, 68, 38, -17, -17, -72, -8, 46, 13, 94, 29, 35, -26, -127, -39, -10, 36, 41, 57, 5, -19, -60, -63, 7, 2, -10, 7, 38, 5, 47, 73, 21, -10, -34, 22, 31, 18, 7, -75, -93, -32, 17, 62, 10, 3, 20, -18, 15, 78, -38, -35, 6, -83, -10, -4, -81, 40, 13, 10, 98, -31, 51, 44, -58, -41, -19, -96, -17, 10, 27, -2, -22, 12, 5, 45, 73, 39, 76, 35, 6, -27, -69, -14, -66, -18, 91, 3, 59, 2, -56, -54, -87, -3, 32, 40, 23, 30, -97, -40, 19, -8, 28, 127, -12, -51, -37, -40, 9, 60, 21, 34, 24, -40, -2, -56, 4, -13, 25, 34, -32, 7, 36, 10, 64, 51, 26, -3, -20, -4, 25, -21, 48, 5, -34, -21, -29, -14, 15, -7, 31, 31, 32, -12, -25, -87, -61, -36, -38, 0, 47, 34, 21, 112, 23, 30, -6, -74, -45, -11, 0, -24, 4, 18, -5, 45, 17, -26, -5, -45, 32, 37, -65, -43, -55, -86, -7, 53, 27, 77, 89, 3, 23, -21, -10, -44, -60, 6, -14, 12, 35, -21, 23, -28, -34, 28, 17, -82, -5, 6, -11, -11, 19, 6, -4, 4, 31, 27, 5, -43, -22, -70, -8, 21, 8, 32, 7, -24, 9, 5, 17, -43, 13, -29, -27, 44, 5, -3, -3, 72, 41, 11, 8, -48, -79, -38, 0, 66, 41, 75, 9, 1, 0, -80, -10, -13, -65, 17, 0, 35, -2, 28, -21, -25, -48, 6, -17, -51, 35, -34, -19, -17, -43, 26, 29, -8, 40, 3, -28, 63, 19, -9, 11, -57, -64, 19, 9, -5, 80, 47, -43, 26, 3, -37, 70, 21, 48, 39, -17, -48, -53, -87, -81, 22, 4, -12, 21, -5, -27, 38, 20, -20, -2, -36, 40, 42, 32, 59, 14, 17, 27, -23, -36, -23, -45, 19, 70, -2, -12, 2, -76, -7, 8, 3, 36, 11, -36, -53, -9, 5, 17, 45, -56, -27, -44, -39, 20, 0, 18, 19, 43, 15, 7, -7, 11, -51, 24, 1, -5, 32, 79, -12, -4, 31, -9, -19, 85, 25, -46, -38, -43, -94, -44, 73, 42, 19, 7, -22, -20, -59, -18, 48, -38, -48, 60, -73, -57, 13, -3, 29, 70, 59, 94, 25, 5, 17, -23, -66, -1, 11, -4, 64, -10, -28, -35, -115, -24, 5, -26, 34, 36, 27, 5, 27, -8, -10, -42, 77, 11, 24, 24, -38, 11, -43, -57, 0, -18, -5, -12, -2, -27, -44, -4, 27, -14, 24, 5, 11, 92, -23, -22, -17, -79, -30, 42, 70, 64, 57, 14, -37, -27, -122, -53, -24, 14, 39, 26, 66, 5, -8, 59, -65, -48, -14, 1, 26, 93, 42, 3, 47, -73, -70, 0, -90, -61, 56, 1, -5, 70, 70, -31, 14, 17, 23, 36, 4, -3, 0, -82, -51, 32, -39, -36, 54, 37, -27, -2, 37, -57, -70, 15, -38, -29, 91, 97, 2, 0, 1, -21, -59, 55, 65, -61, -40, -1, -30, 60, 81, 61, 10, -24, -51, -20, 7, -31, 37, -46, 47, -15, -51, 42, -7, -3, 69, -31, -6, 25, 20, 40, 60, 36, -31, -62, -60, -3, 4, 31, 46, -41, -54, -25, 14, -20, 54, 76, -11, 14, 13, 14, -9, -1, 0, -65, -121, -18, 7, 70, 59, 8, 0, -49, -73, 1, -1, 3, -48, 23, -3, -23, 45, 12, -7, 35, -7, -1, 42, -9, 13, 11, -53, 7, -31, 4, 51, -31, 20, -14, -100, 26, 11, -21, 71, 59, -37, -28, 48, -9, -7, 13, -9, -41, -8, 24, -58, -20, -44, -29, 26, 35, 48, -9, -45, 25, -40, -26, 47, 31, -35, 10, 39, 12, 39, 31, 34, -30, -69, -43, -53, -27, 29, 60, 0, 31, -10, -3, -71, -13, 13, 11, 29, 70, 12, -22, -23, -21, -49, -2, -23, 60, 15, -37, -10, -59, -19, 0, -39, 62, 39, 31, 83, -3, -21, 27, -55, -12, -1, -47, 11, 15, 104, -42, -25, -6, -86, 24, 47, 13, 29, 8, -102, 13, -4, -43, -5, -12, -26, 29, 28, -30, -4, -56, -2, 79, 59, 13, 0, -19, 17, 0, 46, 37, -68, -63, 17, -53, -29, 69, 4, -13, 31, 34, -53, 18, -4, 35, -21, 86, 47, -59, -34, -56, -121, -42, -1, 13, 86, 52, 17, -38, -38, -60, -18, 19, 25, 22, 22, 104, 20, 4, -46, -60, -88, -64, -17, -47, -23, 2, 30, 80, 83, 24, -3, -62, -52, -76, -10, 24, 7, 90, 86, 54, 61, -47, -56, -28, -58, -44, 13, 5, 82, 49, 58, -5, -93, -32, 22, 40, 38, 31, 22, -72, -17, 36, -110, -43, -6, -23, 6, 48, -1, 3, -1, -5, 48, -72, -12, -27, -69, 24, 3, -5, 18, 4, 8, 38, 18, 61, 6, -56, -32, -23, 27, 80, 85, 10, -41, 0, -27, -30, -7, -19, -32, 37, 15, 22, -40, -12, -22, -13, -13, 13, -26, 7, 15, -5, 57, 55, 13, 32, -19, -46, 37, -53, 1, -9, -34, 1, 22, -42, 15, -22, -39, 0, -7, -47, -34, 75, 74, 46, 98, 20, -58, -5, -22, 39, 21, 5, -3, -43, -24, -80, 30, 15, -63, 43, 28, 18, 85, 47, -1, -45, -28, -34, -35, 4, 14, 2, 34, 11, -55, -4, -52, -72, 24, -61, -26, 12, 10, 9, 25, 31, 49, 28, 7, 20, 5, -82, 18, -19, -96, 42, -21, -15, 83, 40, 31, 25, -41, -18, 29, 23, 54, 12, -89, -58, -52, -27, 68, 34, 46, 10, 0, -49, 28, 49, 40, 24, -5, -21, -56, -51, -7, -40, -36, 40, 39, 60, 5, 8, 45, -51, -1, 44, -2, 23, 62, -36, -54, -10, -51, -27, 24, 21, -41, 39, -8, 29, 12, 19, 26, 23, -40, 6, -32, -111, 13, -13, -17, 66, 29, -66, 23, 15, 5, 75, 81, -21, -35, -64, -75, -27, -4, -4, 65, 69, 6, 40, 28, 15, -38, 32, 69, -29, -37, -63, -57, -38, 20, 13, 0, -52, -63, -24, 46, 73, 44, 40, 13, -31, 14, 1, 8, 65, -40, -23, -9, -26, -58, 78, 13, 28, 38, -7, -52, -37, -46, 6, 11, 22, 38, 4, 18, 5, 17, 12, -70, -34, 6, 2, 48, 55, 13, -55, -53, -3, -21, 68, 62, 41, 51, 23, -42, -29, -73, -116, -23, -35, -1, 65, 17, -4, 40, 48, 28, -2, -48, -29, -36, 10, 90, -10, 2, -1, -43, 64, -39, -22, -37, -49, -18, -26, 25, -22, -11, 56, 63, 56, -13, -52, -48, -61, -27, 53, 71, -28, 1, 80, -4, -8, 43, 10, -86, -44, 23, 12, 26, 90, 29, 34, -49, -52, 26, -35, -3, 34, -59, 19, -35, 22, 19, -20, 27, 58, 13, 51, 0, -82, -3, -55, -3, 79, -18, 24, 10, -55, -32, -7, -38, -8, 42, -40, 12, 68, 27, 31, 7, -43, -15, -12, 18, 14, -21, -20, -22, -25, 57, -11, -52, 66, 21, 0, 68, -13, -73, 15, -1, -35, 53, -6, -55, 80, -20, 23, 34, -54, 1, 8, -24, 39, 20, -26, 1, -55, 34, 4, 54, 23, -17, 28, -43, 2, 5, -113, -54, -75, -31, 71, 74, 62, 89, -35, -52, -10, -41, -28, 93, -8, -13, -56, -77, -78, -25, 56, 66, 42, 78, -54, -21, -6, -27, -24, 79, 34, -19, 53, 0, -56, -49, -49, -40, -5, -22, 0, 39, 12, 19, 56, 0, 23, -1, 12, 88, -42, -48, -22, -65, -35, 51, 1, 38, -46, -26, -9, -46, -24, 37, 23, 44, -12, -9, 0, -64, -14, 72, 2, 22, 103, -62, -8, 20, -49, -27, 27, -19, 25, -12, -13, -4, -70, 43, 38, 66, 20, 8, 76, -18, 22, -24, -46, 6, -59, 14, 31, -55, -2, 53, 0, 61, 13, -10, 12, -14, 35, 19, 32, -1, -45, 8, 28, 15, 64, 1, -51, -71, -38, 0, -66, 0, -48, -79, -1, 60, 76, 45, 46, -31, -31, -21, 30, 14, 41, -13, -37, -60, -19, -40, 14, 4, 19, -12, 28, 0, -17, 71, 1, 17, -18, -38, -100, 29, 58, 21, 41, 49, 21, 7, 52, -38, -75, -26, -45, -41, 24, -17, 11, 19, 51, -23, 44, -25, 20, -4, 41, -41, -27, 1, -76, -25, -35, 30, 13, -29, 53, -19, -30, 43, 24, -9, 25, 34, 11, 18, 10, -39, -69, -22, 47, 23, 25, 21, -30, 3, 23, 19, -14, -21, -1, 26, -8, 10, -2, -57, -27, 24, -24, 18, 20, 10, -21, 17, -32, -4, 26, -51, 65, 19, 52, 9, -3, -1, -46, -63, -9, -56, -55, 20, 66, 41, 68, 39, -4, -7, -12, -46, -91, -38, -79, -30, 36, 46, -13, 15, -1, 38, -4, -13, 25, -3, 9, 48, 2, -9, -99, -4, 8, -3, 44, -10, -49, -15, -25, 4, 39, 6, -8, 41, 61, -1, -1, -31, -51, -11, 36, 80, 8, 19, 42, -34, -21, -26, -51, -10, 37, -26, 39, 31, -36, -8, 2, -27, -85, -24, -21, 15, 37, 52, 62, -65, 55, 31, -22, 31, -51, -125, -35, 0, 6, 62, 111, 43, 65, 54, -36, -75, -92, -2, 43, 37, 76, 32, -77, -115, -15, -49, -7, 75, -5, 31, 68, -41, -11, 27, -24, -37, 48, 20, -24, 36, -3, 40, -12, -1, -39, -34, -55, 12, 61, -2, 0, -43, -65, -11, -1, 49, 26, -5, 26, 0, -26, 4, 6, 0, -37, 65, 28, -17, 21, 18, -68, -38, 10, -78, 6, -32, 46, 72, 37, 29, -61, -29, -36, -28, -40, -9, -32, 45, 119, 82, 44, -44, -80, -90, -53, 51, 75, 68, 64, -29, -56, -70, -23, -13, 47, 23, 22, -20, 28, 0, 27, 60, -34, -85, -52, -46, -19, -8, 60, -27, 21, 34, 29, 24, -12, 53, -35, -2, 35, -34, 5, -24, -19, -6, 37, 5, 62, -8, -54, -27, -75, -17, 8, 78, 14, 46, 0, -75, 8, 0, -3, 30, 27, 8, -14, 49, -8, -6, -15, 37, 13, -54, -42, -63, -113, 0, 31, 45, 122, -39, -44, -2, -97, -40, 97, 35, -11, 79, 28, 11, 38, -48, -29, -57, -64, 34, -35, 21, 51, -30, 42, 21, -10, 40, 1, 7, -65, 53, 9, 10, 23, -49, -110, -17, -20, -13, 85, 5, 35, 106, 5, 26, -18, -48, -11, -100, -23, 12, 12, 9, 46, 10, 25, -11, 38, 41, -57, -75, -40, 19, 57, 48, 69, -29, -117, 12, 12, 30, 22, -46, -21, -26, 4, 13, 32, -49, -31, 25, 14, 55, -4, -23, -1, -88, -61, 18, 5, 56, 6, 55, 32, -29, -1, 0, 43, -7, 27, 42, -26, 11, 21, -14, 11, -13, -83, 0, 7, -8, 31, 66, -6, -32, -47, -73, -6, 15, 31, 76, -9, -55, 60, -55, -27, 58, -73, -29, 21, 10, 56, 96, 34, 30, 7, -41, -8, -77, -78, -45, -37, -34, 14, -8, -25, 47, 23, -7, 59, -32, -14, 4, 1, 0, -69, 6, -66, -41, 3, 25, 83, 27, 0, -32, 0, 12, 12, 56, 35, -56, -19, 36, -31, 56, 44, 27, -5, -41, 14, -39, 1, 55, -40, 15, 23, 53, 18, -14, -56, -72, -40, 0, 1, 90, 6, 70, 36, -26, -42, -40, 4, 26, 68, 56, -23, -5, -28, -42, 31, -26, 39, -69, -14, 31, -35, 39, 42, -54, 48, 28, 15, 7, -32, -56, -55, -6, -38, 9, 23, 15, 34, -25, -47, -56, 5, 21, 44, 59, -6, 14, -4, -32, 37, -34, -28, 35, 22, -36, -26, 56, 12, 2, 102, 30, -86, 8, 14, -71, -7, -40, -93, -57, -14, 8, 0, 68, 43, 0, 72, -48, -14, -68, -29, -18, -17, 7, 7, 26, 14, -19, 43, -27, 26, -6, -36, 17, -18, 6, 22, 76, -31, -12, -61, -45, -28, 34, 68, 60, 28, -3, -77, -1, -18, -48, 70, 0, -6, 30, -78, -52, -21, 15, 56, 11, 34, -8, 2, 55, 24, 60, 48, -21, -14, -58, -58, -60, -85, 55, 18, 13, 65, 59, -27, -18, 14, -61, 26, -32, -21, 3, -66, 10, -12, 43, 5, 22, -24, 19, 21, 63, 18, 13, -17, -65, 40, 4, 1, -11, -12, -14, -23, -30, -20, -47, 31, 80, 77, 60, -5, -53, -34, -49, 38, -27, -6, 9, -53, 7, 34, -10, 41, 34, 9, 18, -6, -25, 56, -28, -22, -3, -31, -5, -9, -10, -3, 2, -24, 79, 54, -75, -22, 17, -3, 37, 25, -48, -76, -29, 41, 19, 6, -1, -60, -70, 51, 19, 49, 27, 1, 28, -76, 2, 37, -59, 24, 73, -14, 71, 55, -6, 28, -51, -40, -14, -90, 31, -19, 12, 24, -2, -11, -5, 56, 26, -1, -24, -32, -22, 55, -6, 15, -18, -115, 25, 21, -2, 51, -63, 51, 32, 8, 74, -2, 22, -5, -31, -47, -93, -65, -28, 27, 1, 14, -2, 18, 10, 58, 79, -55, -60, -4, -42, 4, 38, 1, -23, -68, 8, 20, -37, 37, -15, -10, -24, 29, 15, 47, 45, 44, -55, 34, 31, -4, 35, 0, -10, -25, -1, 5, 10, 8, 4, 51, -48, -25, 56, -39, 10, 4, -83, -68, -7, 52, 68, 21, -21, 6, -69, -78, 14, -65, -31, 2, 13, 44, 10, 30, -19, 43, -11, -63, 57, -21, 21, 127, 46, 58, 1, -34, 0, 2, -4, 30, -8, -112, -58, -20, -18, 10, 87, -12, -31, 19, -52, 46, -2, 5, -45, -37, -14, 5, 20, 5, 40, 48, 1, 83, 17, -39, -72, -41, -73, 37, 72, 40, 57, 19, -41, -27, 10, 2, 7, 12, -27, 1, -61, -1, -4, -12, 24, -25, 34, -18, -36, 3, -63, -30, 75, 55, 19, -8, -79, -79, 4, 62, 13, -8, -41, -54, 23, 80, 21, -22, -13, -47, 43, 15, -7, -18, -20, -4, 45, -9, 12, -54, -30, 48, 15, -19, 8, -15, -18, 43, 92, 39, -12, -42, -7, -53, 22, 80, -58, -48, -18, -32, 20, 21, 60, -38, -23, 55, 38, -18, -6, -26, -76, 45, 18, 21, 28, 47, 5, 26, -24, -36, -15, 6, 10, 5, -10, 0, -4, 54, 42, -31, -39, -28, -20, 35, -2, -46, -36, -53, -32, -3, 92, 3, -11, 4, 11, -43, 17, 57, -65, 12, -53, -68, 13, 46, 65, -4, 5, 11, -55, 0, 97, 2, 18, 20, -9, 17, -93, -30, -13, -58, -42, 27, 26, 11, 54, 62, -35, -2, -43, -60, 38, -42, -24, 28, -11, 3, 45, 80, 3, 28, -64, -9, -31, -42, 26, 60, -8, 7, 83, -21, -43, 9, -19, 0, 20, 45, 14, -47, -31, -41, -48, -66, 21, -14, 4, 69, 46, 25, 13, -58, 8, -26, 9, -7, 10, -4, 34, 34, -17, -40, -27, 11, 13, 29, -2, -76, 20, 27, 61, 76, 7, -3, -13, -25, -18, 46, -15, 64, -5, -26, -45, -10, 6, -4, 31, 30, -26, 23, -8, -59, -49, -43, 6, 62, 13, 40, -45, -36, 1, 20, 39, 88, 19, 61, -2, -27, -46, -48, -68, 36, 35, 7, 80, 28, -42, -41, -58, -76, -83, -26, -14, 20, 86, 14, -2, 0, -45, 10, 35, -37, 31, 29, 20, 40, 31, -27, -24, 0, 3, -9, -7, -45, -30, -18, -5, 78, 48, 22, 46, -8, -63, 29, -10, -41, 31, -6, 15, 56, -42, 6, -20, -63, 2, -36, -53, -2, -3, 35, 32, 47, 12, 22, 61, -11, -12, -69, -30, -11, -40, 5, 1, -20, 47, 18, 95, 32, 23, -20, -61, -11, 10, 18, 87, -6, -99, -32, -49, -40, 57, 6, 34, 49, -14, -43, -40, -79, -65, 19, 55, 48, 78, 60, -5, -45, -7, -45, -9, 68, -20, 27, 54, -30, 27, -19, -83, -61, -62, -76, 26, 71, 81, 86, 22, -23, -28, -63, 44, 64, -12, -22, -38, -92, -4, -1, -12, 21, -30, 31, 60, 26, 66, -51, -65, -27, -31, 22, 125, 38, 47, -20, -111, -56, -55, -22, 80, 47, 64, -18, -60, 23, -24, 17, 105, 2, 3, -59, -1, -41, -60, 74, -8, -1, 0, -27, -29, 17, -15, 17, -30, -35, 12, 64, 68, 51, 19, 12, -18, 3, -26, -54, -65, -49, -26, 90, 8, -8, 51, -55, -54, 55, 7, -5, 65, -34, -10, -40, -9, 20, 45, 55, -22, -22, 6, -76, -36, -18, -18, 10, 49, 105, 4, 3, 11, -83, 25, 20, 0, 36, 55, -51, -89, -44, -51, -24, 18, 105, -2, -21, -19, -32, 0, -3, 9, -7, 0, 32, 23, 38, -21, 35, -8, 20, 3, -29, -53, -25, -5, 1, 39, -20, 3, -62, 37, -22, -61, 21, -45, 5, 43, 25, 42, 8, -28, 1, 8, -3, -10, 14, -9, 26, -22, 34, 1, 4, -37, 31, -1, -32, -19, 22, 0, 1, 29, -44, 24, -30, -5, 78, -4, -39, 24, 9, -59, 47, 28, 22, -4, -48, 12, -6, -4, 89, -17, -74, -27, -79, 18, 59, 29, 34, 43, -21, 59, 23, 34, -10, -64, -37, -19, -28, 112, 22, 39, 11, -11, -1, -38, 0, -68, -45, -12, -38, -56, 17, 3, 1, 73, 126, -4, -3, -5, -70, -65, 29, -57, 9, 55, -19, -14, 47, 10, -1, 98, 53, -28, -34, -53, -66, 0, -25, 4, 24, 6, 71, 39, 13, -24, -108, -47, -25, -7, 59, 58, 32, 23, -7, -45, -14, -30, 68, -24, -23, 0, -57, -20, 31, -55, -24, -44, 35, 86, 35, 61, 69, -72, -17, -32, -51, 31, 5, 26, 83, 27, 37, 12, -38, -61, -105, -40, -37, -53, 46, 41, 32, 78, -14, -15, -74, -49, -30, -47, 6, 34, 28, -4, 62, -39, -7, 0, -25, 9, 34, -6, 24, -54, -31, -6, 8, -12, 53, 40, -28, -6, -61, -59, -29, 20, 15, 49, 68, 60, 15, 30, -2, -90, -21, -6, 19, -5, -24, 29, 38, 1, 15, 10, -23, -25, 28, -25, -11, -14, -79, 8, 7, 14, -6, 40, -15, -31, -9, -23, -5, 7, 60, -15, -44, -14, -71, -43, 15, 25, -3, 28, 3, 31, 70, 28, 28, 17, 53, -70, -20, -1, -90, -44, 7, 14, 34, 8, -20, 34, -66, -30, 28, -10, 44, 56, -18, 45, 47, 2, 68, -29, -62, -12, -38, 56, 43, -20, -65, -12, -2, -5, 43, 18, 39, -1, 41, 38, -78, -69, -52, -18, 26, 72, 7, 3, -11, -49, 20, -79, 19, -42, -57, 44, 36, 60, 30, 57, 24, -42, 21, -23, -36, -40, -24, 6, 28, -15, 34, -48, -52, 12, -18, -19, 21, 11, 60, 2, 49, 77, -58, 34, 26, -36, 18, -27, 12, -24, -14, -14, -7, -10, -19, -65, -36, -74, -45, -7, 45, 90, 45, 52, 12, -88, 3, 25, 60, 78, 64, 46, -34, -27, -58, -51, -6, -30, 14, 42, -43, 61, 20, -44, -45, -31, -53, 22, 55, -9, 76, 10, 38, 12, -43, -35, -46, -46, 22, 68, -6, -5, 27, -35, -88, 14, -28, -23, 98, 56, 76, 65, -39, -74, -8, -22, -37, 13, -65, -35, -9, 27, 15, 3, 13, -45, 27, 54, -34, 31, 44, -11, -24, 53, 40, 6, 70, 42, -5, -23, -34, -3, -4, 6, -27, -40, 15, -11, 0, 29, 32, -37, 3, 17, -11, -43, -24, -47, -2, 19, 98, 31, 19, -45, -55, 7, 11, 25, -57, -52, -70, -24, 60, 104, 39, 71, -17, 1, 45, -12, -13, -66, -27, -2, 48, 41, 2, -20, -69, -53, -37, 26, 13, -21, 53, 66, -17, -20, -8, -47, -43, 3, 13, 40, -31, 65, 1, -29, -18, -38, -32, 102, 58, 14, -23, -47, -62, 31, 4, -3, 53, -68, -22, 38, -3, 30, -23, -21, -63, -87, -14, 5, 42, 54, -7, -5, -9, -13, 14, 77, 71, -20, -31, 3, -78, -48, 40, -18, -54, 41, 32, 17, 46, 88, -41, 14, -19, -52, 25, 26, 60, 4, 6, 1, -66, -31, -11, -34, 2, 41, -52, -23, -60, -21, 21, 8, 65, -18, 17, 46, 3, 64, -72, -59, -10, -53, -13, 86, 17, 0, 13, -28, 40, -28, 4, 72, -60, -28, 37, 6, -30, 61, 36, -31, -42, -31, -66, -41, 42, 28, 59, 3, -39, -35, 0, 1, 18, 41, -35, 11, -10, 70, -7, 6, 6, -60, -12, -20, 5, 24, 58, 29, 4, 8, -23, 52, -23, 10, 19, -52, -28, 1, -8, -13, -29, 52, -28, -68, -18, -39, 5, 75, 48, 71, -29, 0, 44, -9, 72, 17, -42, -37, 29, -62, -3, -13, -87, 3, 34, 30, 60, 14, -17, 4, -105, -19, -42, -47, 34, 53, -30, 8, -29, -48, -2, 0, 18, 14, 61, 38, 49, -40, 19, -14, -59, 53, -13, 60, 26, 32, -21, -35, -56, -40, -1, -35, 20, 42, -18, 39, 66, -34, 26, 51, 31, 24, -37, -97, -53, -49, -1, 80, 105, -11, 26, 31, -62, -8, 42, -95, 7, -11, -90, 20, -28, -1, -14, 39, -6, 38, 68, 35, 35, 57, -13, 1, -4, -1, -52, -18, -29, -80, -44, 40, 56, 38, 35, 38, 0, -68, -19, -45, -56, 29, 65, 23, 5, 26, -52, -28, 29, 15, -18, 72, 30, 32, -42, -31, -46, -23, -15, -10, 52, 22, -5, -11, 19, -37, -17, 54, -20, -54, 26, -31, -72, 79, 4, -9, 109, 29, 26, 52, -8, -1, 0, -24, -30, 10, -41, -9, 69, -47, 31, 10, -99, -32, 22, 63, 61, 85, 7, -90, -103, -72, -48, 48, 53, 5, 19, -15, 3, -23, -5, -5, -20, 36, 88, 51, 48, 15, -68, -57, 27, -35, 34, 90, 18, 39, 38, 35, 4, -45, -55, -11, -69, -20, 38, 4, 2, -13, -30, -18, -29, 4, 43, 20, 62, 6, -15, 15, 14, 17, 21, -30, -56, -49, -45, 23, 8, 39, -44, 14, 62, 2, 25, 13, 17, -59, -12, 20, -3, 10, 76, -34, -66, -57, -20, 48, 85, 127, -8, -81, -23, -39, -71, 14, -15, -21, 32, -8, 76, 17, -6, 8, -18, -71, 39, 15, 25, 17, -29, 3, -43, 42, 41, -82, -39, -56, -9, 43, 42, 88, -37, -51, -72, -31, 28, 41, 38, 36, -32, 27, -4, 38, -18, -78, 0, -8, 22, 85, 31, -26, -59, 40, 18, 1, 28, -21, -102, -77, 41, 0, -21, 85, -39, -79, 73, 13, -10, 34, -55, -23, 15, 44, 65, 19, -13, -65, 13, 7, 49, 40, -17, -63, -2, -19, -56, 80, 38, 2, 102, 1, -34, -60, -79, -31, -21, -28, 27, -37, 42, 79, 63, 81, -27, -52, 6, -52, 0, 86, 10, -64, -43, -43, -74, 31, 57, 4, 71, 25, -2, -6, -22, -26, 17, -8, 61, -36, -113, -10, -7, 18, 29, 96, 32, 1, 14, 11, -53, -90, -27, -63, -66, -11, 37, 29, -6, 19, 32, -24, -3, 65, 20, -4, 22, -32, 43, 5, -13, 1, -47, -79, 3, 62, 0, 18, -13, -83, -61, 17, 38, 17, 60, 52, -72, -39, -20, -24, 49, 66, 43, 41, -37, 32, -14, -1, -40, -8, -27, -39, 54, -2, 59, 2, 36, -7, -69, -8, -106, -19, 11, 22, 90, 87, 22, -11, -96, -65, -73, 0, 41, -31, 24, -29, -31, 92, 98, 65, 34, -39, -58, -51, 19, 13, 71, -36, -4, 27, -10, 47, 12, -20, -21, 10, -58, 26, 62, -62, 37, 49, -48, 38, -17, -6, -53, -78, -5, -10, -6, 36, 19, -41, -63, -19, -35, 18, 49, 15, 39, 13, -4, -26, -45, -29, -39, 41, 88, 18, 14, 6, 3, 27, 1, -4, -6, -73, -13, -26, 1, 12, 56, 20, -12, -20, -31, -41, 23, 76, -25, 6, 3, -5, -12, 1, 3, 36, 31, -11, -29, -47, -32, 20, 88, 108, 38, -43, -48, -37, -69, -25, -1, -49, -5, -10, 70, 52, 25, 13, -34, -8, -26, 8, 31, -26, -71, -9, -31, -21, 75, 91, 10, 26, 5, -42, -79, -12, 23, 11, -6, 23, -9, 5, 34, 74, 53, 8, -25, -38, -21, -45, 40, -18, 4, -22, -23, 64, 28, 66, 39, -57, -13, -51, -35, 40, -66, -10, 1, -9, 24, -21, 5, -41, 20, 57, 42, 70, 0, 36, 31, -19, -51, -44, -26, -46, 0, -2, -24, -57, -2, -27, 1, -14, -8, 39, 9, 0, 32, 43, 43, 11, 10, -12, -51, -15, 30, 7, 9, 1, -20, -10, 47, -58, -47, -25, -78, 5, 88, 79, 53, 22, -30, -70, -52, -34, -9, 43, 30, 17, -26, -56, -35, -31, 22, 53, 40, 79, 17, -2, 20, -24, -58, 21, -36, -97, -14, -13, -31, -7, 75, 7, -48, 40, 2, -42, 41, 23, -70, 30, 4, -22, 19, 15, -72, -1, -15, -27, 26, -2, -12, 14, -45, 14, 11, 34, -21, 13, -8, 5, 119, 59, 88, 14, -79, -53, -29, -13, 19, 28, 10, -46, -20, -3, 7, 25, -19, -25, 25, -28, 0, 28, 0, 1, 4, 23, -39, -85, -68, -55, 10, 47, 12, 46, -2, 12, -12, 17, -29, -17, 3, -35, 46, -51, -41, 27, 39, 43, 48, -14, -22, -2, -3, 43, 44, -66, 30, -4, -34, 26, -47, -2, 64, -12, 53, 25, -83, 18, -40, -46, 15, 17, -11, 38, 87, -56, 15, 57, -28, -8, -36, -46, -14, 19, 6, 48, 66, -7, 54, 53, -26, -57, -38, -49, -70, -27, 47, 13, 12 );

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
